VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpu_core
  CLASS BLOCK ;
  FOREIGN gpu_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END ack
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END clk
  PIN command[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END command[0]
  PIN command[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END command[10]
  PIN command[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 0.000 622.160 4.000 ;
    END
  END command[11]
  PIN command[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 664.160 0.000 664.720 4.000 ;
    END
  END command[12]
  PIN command[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 0.000 707.280 4.000 ;
    END
  END command[13]
  PIN command[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END command[14]
  PIN command[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 791.840 0.000 792.400 4.000 ;
    END
  END command[15]
  PIN command[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 834.400 0.000 834.960 4.000 ;
    END
  END command[16]
  PIN command[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 0.000 877.520 4.000 ;
    END
  END command[17]
  PIN command[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 919.520 0.000 920.080 4.000 ;
    END
  END command[18]
  PIN command[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 0.000 962.640 4.000 ;
    END
  END command[19]
  PIN command[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END command[1]
  PIN command[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 0.000 1005.200 4.000 ;
    END
  END command[20]
  PIN command[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1047.200 0.000 1047.760 4.000 ;
    END
  END command[21]
  PIN command[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1089.760 0.000 1090.320 4.000 ;
    END
  END command[22]
  PIN command[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 0.000 1132.880 4.000 ;
    END
  END command[23]
  PIN command[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1174.880 0.000 1175.440 4.000 ;
    END
  END command[24]
  PIN command[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1217.440 0.000 1218.000 4.000 ;
    END
  END command[25]
  PIN command[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1260.000 0.000 1260.560 4.000 ;
    END
  END command[26]
  PIN command[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1302.560 0.000 1303.120 4.000 ;
    END
  END command[27]
  PIN command[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1345.120 0.000 1345.680 4.000 ;
    END
  END command[28]
  PIN command[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1387.680 0.000 1388.240 4.000 ;
    END
  END command[29]
  PIN command[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END command[2]
  PIN command[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1430.240 0.000 1430.800 4.000 ;
    END
  END command[30]
  PIN command[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1472.800 0.000 1473.360 4.000 ;
    END
  END command[31]
  PIN command[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 4.000 ;
    END
  END command[3]
  PIN command[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END command[4]
  PIN command[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END command[5]
  PIN command[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END command[6]
  PIN command[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END command[7]
  PIN command[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 0.000 494.480 4.000 ;
    END
  END command[8]
  PIN command[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 0.000 537.040 4.000 ;
    END
  END command[9]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 43.680 1500.000 44.240 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 267.680 1500.000 268.240 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 290.080 1500.000 290.640 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 312.480 1500.000 313.040 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 334.880 1500.000 335.440 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 357.280 1500.000 357.840 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 379.680 1500.000 380.240 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 402.080 1500.000 402.640 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 424.480 1500.000 425.040 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 446.880 1500.000 447.440 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 469.280 1500.000 469.840 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 66.080 1500.000 66.640 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 491.680 1500.000 492.240 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 514.080 1500.000 514.640 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 536.480 1500.000 537.040 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 558.880 1500.000 559.440 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 581.280 1500.000 581.840 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 603.680 1500.000 604.240 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 626.080 1500.000 626.640 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 648.480 1500.000 649.040 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 670.880 1500.000 671.440 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 693.280 1500.000 693.840 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 88.480 1500.000 89.040 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 715.680 1500.000 716.240 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 738.080 1500.000 738.640 ;
    END
  END data_in[31]
  PIN data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 760.480 1500.000 761.040 ;
    END
  END data_in[32]
  PIN data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 782.880 1500.000 783.440 ;
    END
  END data_in[33]
  PIN data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 805.280 1500.000 805.840 ;
    END
  END data_in[34]
  PIN data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 827.680 1500.000 828.240 ;
    END
  END data_in[35]
  PIN data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 850.080 1500.000 850.640 ;
    END
  END data_in[36]
  PIN data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 872.480 1500.000 873.040 ;
    END
  END data_in[37]
  PIN data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 894.880 1500.000 895.440 ;
    END
  END data_in[38]
  PIN data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 917.280 1500.000 917.840 ;
    END
  END data_in[39]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 110.880 1500.000 111.440 ;
    END
  END data_in[3]
  PIN data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 939.680 1500.000 940.240 ;
    END
  END data_in[40]
  PIN data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 962.080 1500.000 962.640 ;
    END
  END data_in[41]
  PIN data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 984.480 1500.000 985.040 ;
    END
  END data_in[42]
  PIN data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1006.880 1500.000 1007.440 ;
    END
  END data_in[43]
  PIN data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1029.280 1500.000 1029.840 ;
    END
  END data_in[44]
  PIN data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1051.680 1500.000 1052.240 ;
    END
  END data_in[45]
  PIN data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1074.080 1500.000 1074.640 ;
    END
  END data_in[46]
  PIN data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1096.480 1500.000 1097.040 ;
    END
  END data_in[47]
  PIN data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1118.880 1500.000 1119.440 ;
    END
  END data_in[48]
  PIN data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1141.280 1500.000 1141.840 ;
    END
  END data_in[49]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 133.280 1500.000 133.840 ;
    END
  END data_in[4]
  PIN data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1163.680 1500.000 1164.240 ;
    END
  END data_in[50]
  PIN data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1186.080 1500.000 1186.640 ;
    END
  END data_in[51]
  PIN data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1208.480 1500.000 1209.040 ;
    END
  END data_in[52]
  PIN data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1230.880 1500.000 1231.440 ;
    END
  END data_in[53]
  PIN data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1253.280 1500.000 1253.840 ;
    END
  END data_in[54]
  PIN data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1275.680 1500.000 1276.240 ;
    END
  END data_in[55]
  PIN data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1298.080 1500.000 1298.640 ;
    END
  END data_in[56]
  PIN data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1320.480 1500.000 1321.040 ;
    END
  END data_in[57]
  PIN data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1342.880 1500.000 1343.440 ;
    END
  END data_in[58]
  PIN data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1365.280 1500.000 1365.840 ;
    END
  END data_in[59]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 155.680 1500.000 156.240 ;
    END
  END data_in[5]
  PIN data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1387.680 1500.000 1388.240 ;
    END
  END data_in[60]
  PIN data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1410.080 1500.000 1410.640 ;
    END
  END data_in[61]
  PIN data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1432.480 1500.000 1433.040 ;
    END
  END data_in[62]
  PIN data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1454.880 1500.000 1455.440 ;
    END
  END data_in[63]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 178.080 1500.000 178.640 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 200.480 1500.000 201.040 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 222.880 1500.000 223.440 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 245.280 1500.000 245.840 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1454.880 4.000 1455.440 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1230.880 4.000 1231.440 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1208.480 4.000 1209.040 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1186.080 4.000 1186.640 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1163.680 4.000 1164.240 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1141.280 4.000 1141.840 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1118.880 4.000 1119.440 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1096.480 4.000 1097.040 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1074.080 4.000 1074.640 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1051.680 4.000 1052.240 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1029.280 4.000 1029.840 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1432.480 4.000 1433.040 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1006.880 4.000 1007.440 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 984.480 4.000 985.040 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 962.080 4.000 962.640 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 939.680 4.000 940.240 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 917.280 4.000 917.840 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 894.880 4.000 895.440 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 872.480 4.000 873.040 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 850.080 4.000 850.640 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 827.680 4.000 828.240 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 805.280 4.000 805.840 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1410.080 4.000 1410.640 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 782.880 4.000 783.440 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 760.480 4.000 761.040 ;
    END
  END data_out[31]
  PIN data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 738.080 4.000 738.640 ;
    END
  END data_out[32]
  PIN data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 715.680 4.000 716.240 ;
    END
  END data_out[33]
  PIN data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 693.280 4.000 693.840 ;
    END
  END data_out[34]
  PIN data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 670.880 4.000 671.440 ;
    END
  END data_out[35]
  PIN data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 648.480 4.000 649.040 ;
    END
  END data_out[36]
  PIN data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.080 4.000 626.640 ;
    END
  END data_out[37]
  PIN data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 603.680 4.000 604.240 ;
    END
  END data_out[38]
  PIN data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 4.000 581.840 ;
    END
  END data_out[39]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1387.680 4.000 1388.240 ;
    END
  END data_out[3]
  PIN data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 4.000 559.440 ;
    END
  END data_out[40]
  PIN data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 536.480 4.000 537.040 ;
    END
  END data_out[41]
  PIN data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END data_out[42]
  PIN data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.680 4.000 492.240 ;
    END
  END data_out[43]
  PIN data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.280 4.000 469.840 ;
    END
  END data_out[44]
  PIN data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 446.880 4.000 447.440 ;
    END
  END data_out[45]
  PIN data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 424.480 4.000 425.040 ;
    END
  END data_out[46]
  PIN data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.080 4.000 402.640 ;
    END
  END data_out[47]
  PIN data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.680 4.000 380.240 ;
    END
  END data_out[48]
  PIN data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 357.280 4.000 357.840 ;
    END
  END data_out[49]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1365.280 4.000 1365.840 ;
    END
  END data_out[4]
  PIN data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.880 4.000 335.440 ;
    END
  END data_out[50]
  PIN data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END data_out[51]
  PIN data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.080 4.000 290.640 ;
    END
  END data_out[52]
  PIN data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.680 4.000 268.240 ;
    END
  END data_out[53]
  PIN data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 4.000 245.840 ;
    END
  END data_out[54]
  PIN data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.880 4.000 223.440 ;
    END
  END data_out[55]
  PIN data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.480 4.000 201.040 ;
    END
  END data_out[56]
  PIN data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END data_out[57]
  PIN data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 4.000 156.240 ;
    END
  END data_out[58]
  PIN data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 4.000 133.840 ;
    END
  END data_out[59]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1342.880 4.000 1343.440 ;
    END
  END data_out[5]
  PIN data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END data_out[60]
  PIN data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 4.000 89.040 ;
    END
  END data_out[61]
  PIN data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END data_out[62]
  PIN data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END data_out[63]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1320.480 4.000 1321.040 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1298.080 4.000 1298.640 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1275.680 4.000 1276.240 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1253.280 4.000 1253.840 ;
    END
  END data_out[9]
  PIN stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 4.000 ;
    END
  END stb
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1482.060 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1482.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1482.060 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1492.960 1482.060 ;
      LAYER Metal2 ;
        RECT 7.420 4.300 1493.940 1481.950 ;
        RECT 7.420 3.500 25.460 4.300 ;
        RECT 26.620 3.500 68.020 4.300 ;
        RECT 69.180 3.500 110.580 4.300 ;
        RECT 111.740 3.500 153.140 4.300 ;
        RECT 154.300 3.500 195.700 4.300 ;
        RECT 196.860 3.500 238.260 4.300 ;
        RECT 239.420 3.500 280.820 4.300 ;
        RECT 281.980 3.500 323.380 4.300 ;
        RECT 324.540 3.500 365.940 4.300 ;
        RECT 367.100 3.500 408.500 4.300 ;
        RECT 409.660 3.500 451.060 4.300 ;
        RECT 452.220 3.500 493.620 4.300 ;
        RECT 494.780 3.500 536.180 4.300 ;
        RECT 537.340 3.500 578.740 4.300 ;
        RECT 579.900 3.500 621.300 4.300 ;
        RECT 622.460 3.500 663.860 4.300 ;
        RECT 665.020 3.500 706.420 4.300 ;
        RECT 707.580 3.500 748.980 4.300 ;
        RECT 750.140 3.500 791.540 4.300 ;
        RECT 792.700 3.500 834.100 4.300 ;
        RECT 835.260 3.500 876.660 4.300 ;
        RECT 877.820 3.500 919.220 4.300 ;
        RECT 920.380 3.500 961.780 4.300 ;
        RECT 962.940 3.500 1004.340 4.300 ;
        RECT 1005.500 3.500 1046.900 4.300 ;
        RECT 1048.060 3.500 1089.460 4.300 ;
        RECT 1090.620 3.500 1132.020 4.300 ;
        RECT 1133.180 3.500 1174.580 4.300 ;
        RECT 1175.740 3.500 1217.140 4.300 ;
        RECT 1218.300 3.500 1259.700 4.300 ;
        RECT 1260.860 3.500 1302.260 4.300 ;
        RECT 1303.420 3.500 1344.820 4.300 ;
        RECT 1345.980 3.500 1387.380 4.300 ;
        RECT 1388.540 3.500 1429.940 4.300 ;
        RECT 1431.100 3.500 1472.500 4.300 ;
        RECT 1473.660 3.500 1493.940 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1455.740 1496.000 1481.900 ;
        RECT 4.300 1454.580 1495.700 1455.740 ;
        RECT 4.000 1433.340 1496.000 1454.580 ;
        RECT 4.300 1432.180 1495.700 1433.340 ;
        RECT 4.000 1410.940 1496.000 1432.180 ;
        RECT 4.300 1409.780 1495.700 1410.940 ;
        RECT 4.000 1388.540 1496.000 1409.780 ;
        RECT 4.300 1387.380 1495.700 1388.540 ;
        RECT 4.000 1366.140 1496.000 1387.380 ;
        RECT 4.300 1364.980 1495.700 1366.140 ;
        RECT 4.000 1343.740 1496.000 1364.980 ;
        RECT 4.300 1342.580 1495.700 1343.740 ;
        RECT 4.000 1321.340 1496.000 1342.580 ;
        RECT 4.300 1320.180 1495.700 1321.340 ;
        RECT 4.000 1298.940 1496.000 1320.180 ;
        RECT 4.300 1297.780 1495.700 1298.940 ;
        RECT 4.000 1276.540 1496.000 1297.780 ;
        RECT 4.300 1275.380 1495.700 1276.540 ;
        RECT 4.000 1254.140 1496.000 1275.380 ;
        RECT 4.300 1252.980 1495.700 1254.140 ;
        RECT 4.000 1231.740 1496.000 1252.980 ;
        RECT 4.300 1230.580 1495.700 1231.740 ;
        RECT 4.000 1209.340 1496.000 1230.580 ;
        RECT 4.300 1208.180 1495.700 1209.340 ;
        RECT 4.000 1186.940 1496.000 1208.180 ;
        RECT 4.300 1185.780 1495.700 1186.940 ;
        RECT 4.000 1164.540 1496.000 1185.780 ;
        RECT 4.300 1163.380 1495.700 1164.540 ;
        RECT 4.000 1142.140 1496.000 1163.380 ;
        RECT 4.300 1140.980 1495.700 1142.140 ;
        RECT 4.000 1119.740 1496.000 1140.980 ;
        RECT 4.300 1118.580 1495.700 1119.740 ;
        RECT 4.000 1097.340 1496.000 1118.580 ;
        RECT 4.300 1096.180 1495.700 1097.340 ;
        RECT 4.000 1074.940 1496.000 1096.180 ;
        RECT 4.300 1073.780 1495.700 1074.940 ;
        RECT 4.000 1052.540 1496.000 1073.780 ;
        RECT 4.300 1051.380 1495.700 1052.540 ;
        RECT 4.000 1030.140 1496.000 1051.380 ;
        RECT 4.300 1028.980 1495.700 1030.140 ;
        RECT 4.000 1007.740 1496.000 1028.980 ;
        RECT 4.300 1006.580 1495.700 1007.740 ;
        RECT 4.000 985.340 1496.000 1006.580 ;
        RECT 4.300 984.180 1495.700 985.340 ;
        RECT 4.000 962.940 1496.000 984.180 ;
        RECT 4.300 961.780 1495.700 962.940 ;
        RECT 4.000 940.540 1496.000 961.780 ;
        RECT 4.300 939.380 1495.700 940.540 ;
        RECT 4.000 918.140 1496.000 939.380 ;
        RECT 4.300 916.980 1495.700 918.140 ;
        RECT 4.000 895.740 1496.000 916.980 ;
        RECT 4.300 894.580 1495.700 895.740 ;
        RECT 4.000 873.340 1496.000 894.580 ;
        RECT 4.300 872.180 1495.700 873.340 ;
        RECT 4.000 850.940 1496.000 872.180 ;
        RECT 4.300 849.780 1495.700 850.940 ;
        RECT 4.000 828.540 1496.000 849.780 ;
        RECT 4.300 827.380 1495.700 828.540 ;
        RECT 4.000 806.140 1496.000 827.380 ;
        RECT 4.300 804.980 1495.700 806.140 ;
        RECT 4.000 783.740 1496.000 804.980 ;
        RECT 4.300 782.580 1495.700 783.740 ;
        RECT 4.000 761.340 1496.000 782.580 ;
        RECT 4.300 760.180 1495.700 761.340 ;
        RECT 4.000 738.940 1496.000 760.180 ;
        RECT 4.300 737.780 1495.700 738.940 ;
        RECT 4.000 716.540 1496.000 737.780 ;
        RECT 4.300 715.380 1495.700 716.540 ;
        RECT 4.000 694.140 1496.000 715.380 ;
        RECT 4.300 692.980 1495.700 694.140 ;
        RECT 4.000 671.740 1496.000 692.980 ;
        RECT 4.300 670.580 1495.700 671.740 ;
        RECT 4.000 649.340 1496.000 670.580 ;
        RECT 4.300 648.180 1495.700 649.340 ;
        RECT 4.000 626.940 1496.000 648.180 ;
        RECT 4.300 625.780 1495.700 626.940 ;
        RECT 4.000 604.540 1496.000 625.780 ;
        RECT 4.300 603.380 1495.700 604.540 ;
        RECT 4.000 582.140 1496.000 603.380 ;
        RECT 4.300 580.980 1495.700 582.140 ;
        RECT 4.000 559.740 1496.000 580.980 ;
        RECT 4.300 558.580 1495.700 559.740 ;
        RECT 4.000 537.340 1496.000 558.580 ;
        RECT 4.300 536.180 1495.700 537.340 ;
        RECT 4.000 514.940 1496.000 536.180 ;
        RECT 4.300 513.780 1495.700 514.940 ;
        RECT 4.000 492.540 1496.000 513.780 ;
        RECT 4.300 491.380 1495.700 492.540 ;
        RECT 4.000 470.140 1496.000 491.380 ;
        RECT 4.300 468.980 1495.700 470.140 ;
        RECT 4.000 447.740 1496.000 468.980 ;
        RECT 4.300 446.580 1495.700 447.740 ;
        RECT 4.000 425.340 1496.000 446.580 ;
        RECT 4.300 424.180 1495.700 425.340 ;
        RECT 4.000 402.940 1496.000 424.180 ;
        RECT 4.300 401.780 1495.700 402.940 ;
        RECT 4.000 380.540 1496.000 401.780 ;
        RECT 4.300 379.380 1495.700 380.540 ;
        RECT 4.000 358.140 1496.000 379.380 ;
        RECT 4.300 356.980 1495.700 358.140 ;
        RECT 4.000 335.740 1496.000 356.980 ;
        RECT 4.300 334.580 1495.700 335.740 ;
        RECT 4.000 313.340 1496.000 334.580 ;
        RECT 4.300 312.180 1495.700 313.340 ;
        RECT 4.000 290.940 1496.000 312.180 ;
        RECT 4.300 289.780 1495.700 290.940 ;
        RECT 4.000 268.540 1496.000 289.780 ;
        RECT 4.300 267.380 1495.700 268.540 ;
        RECT 4.000 246.140 1496.000 267.380 ;
        RECT 4.300 244.980 1495.700 246.140 ;
        RECT 4.000 223.740 1496.000 244.980 ;
        RECT 4.300 222.580 1495.700 223.740 ;
        RECT 4.000 201.340 1496.000 222.580 ;
        RECT 4.300 200.180 1495.700 201.340 ;
        RECT 4.000 178.940 1496.000 200.180 ;
        RECT 4.300 177.780 1495.700 178.940 ;
        RECT 4.000 156.540 1496.000 177.780 ;
        RECT 4.300 155.380 1495.700 156.540 ;
        RECT 4.000 134.140 1496.000 155.380 ;
        RECT 4.300 132.980 1495.700 134.140 ;
        RECT 4.000 111.740 1496.000 132.980 ;
        RECT 4.300 110.580 1495.700 111.740 ;
        RECT 4.000 89.340 1496.000 110.580 ;
        RECT 4.300 88.180 1495.700 89.340 ;
        RECT 4.000 66.940 1496.000 88.180 ;
        RECT 4.300 65.780 1495.700 66.940 ;
        RECT 4.000 44.540 1496.000 65.780 ;
        RECT 4.300 43.380 1495.700 44.540 ;
        RECT 4.000 15.540 1496.000 43.380 ;
      LAYER Metal4 ;
        RECT 44.380 233.050 98.740 1252.070 ;
        RECT 100.940 233.050 175.540 1252.070 ;
        RECT 177.740 233.050 252.340 1252.070 ;
        RECT 254.540 233.050 329.140 1252.070 ;
        RECT 331.340 233.050 405.940 1252.070 ;
        RECT 408.140 233.050 482.740 1252.070 ;
        RECT 484.940 233.050 559.540 1252.070 ;
        RECT 561.740 233.050 636.340 1252.070 ;
        RECT 638.540 233.050 713.140 1252.070 ;
        RECT 715.340 233.050 789.940 1252.070 ;
        RECT 792.140 233.050 866.740 1252.070 ;
        RECT 868.940 233.050 943.540 1252.070 ;
        RECT 945.740 233.050 1020.340 1252.070 ;
        RECT 1022.540 233.050 1097.140 1252.070 ;
        RECT 1099.340 233.050 1173.940 1252.070 ;
        RECT 1176.140 233.050 1250.740 1252.070 ;
        RECT 1252.940 233.050 1327.540 1252.070 ;
        RECT 1329.740 233.050 1404.340 1252.070 ;
        RECT 1406.540 233.050 1475.460 1252.070 ;
  END
END gpu_core
END LIBRARY

