VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tinyrv
  CLASS BLOCK ;
  FOREIGN tinyrv ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 600.000 ;
  PIN alu_out_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 596.000 246.960 600.000 ;
    END
  END alu_out_out[0]
  PIN alu_out_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 596.000 179.760 600.000 ;
    END
  END alu_out_out[10]
  PIN alu_out_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 596.000 173.040 600.000 ;
    END
  END alu_out_out[11]
  PIN alu_out_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 596.000 166.320 600.000 ;
    END
  END alu_out_out[12]
  PIN alu_out_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 596.000 159.600 600.000 ;
    END
  END alu_out_out[13]
  PIN alu_out_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 596.000 152.880 600.000 ;
    END
  END alu_out_out[14]
  PIN alu_out_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 596.000 146.160 600.000 ;
    END
  END alu_out_out[15]
  PIN alu_out_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 596.000 139.440 600.000 ;
    END
  END alu_out_out[16]
  PIN alu_out_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 596.000 132.720 600.000 ;
    END
  END alu_out_out[17]
  PIN alu_out_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 596.000 126.000 600.000 ;
    END
  END alu_out_out[18]
  PIN alu_out_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 596.000 119.280 600.000 ;
    END
  END alu_out_out[19]
  PIN alu_out_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 596.000 240.240 600.000 ;
    END
  END alu_out_out[1]
  PIN alu_out_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 596.000 112.560 600.000 ;
    END
  END alu_out_out[20]
  PIN alu_out_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 596.000 105.840 600.000 ;
    END
  END alu_out_out[21]
  PIN alu_out_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 596.000 99.120 600.000 ;
    END
  END alu_out_out[22]
  PIN alu_out_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 596.000 92.400 600.000 ;
    END
  END alu_out_out[23]
  PIN alu_out_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 596.000 85.680 600.000 ;
    END
  END alu_out_out[24]
  PIN alu_out_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 596.000 78.960 600.000 ;
    END
  END alu_out_out[25]
  PIN alu_out_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 596.000 72.240 600.000 ;
    END
  END alu_out_out[26]
  PIN alu_out_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 596.000 65.520 600.000 ;
    END
  END alu_out_out[27]
  PIN alu_out_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 596.000 58.800 600.000 ;
    END
  END alu_out_out[28]
  PIN alu_out_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 596.000 52.080 600.000 ;
    END
  END alu_out_out[29]
  PIN alu_out_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 596.000 233.520 600.000 ;
    END
  END alu_out_out[2]
  PIN alu_out_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 596.000 45.360 600.000 ;
    END
  END alu_out_out[30]
  PIN alu_out_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 596.000 38.640 600.000 ;
    END
  END alu_out_out[31]
  PIN alu_out_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 596.000 226.800 600.000 ;
    END
  END alu_out_out[3]
  PIN alu_out_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 596.000 220.080 600.000 ;
    END
  END alu_out_out[4]
  PIN alu_out_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 596.000 213.360 600.000 ;
    END
  END alu_out_out[5]
  PIN alu_out_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 596.000 206.640 600.000 ;
    END
  END alu_out_out[6]
  PIN alu_out_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 596.000 199.920 600.000 ;
    END
  END alu_out_out[7]
  PIN alu_out_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 596.000 193.200 600.000 ;
    END
  END alu_out_out[8]
  PIN alu_out_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 596.000 186.480 600.000 ;
    END
  END alu_out_out[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 4.000 ;
    END
  END clk
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 4.000 ;
    END
  END inst[0]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END inst[10]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END inst[11]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 4.000 ;
    END
  END inst[12]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END inst[13]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 4.000 ;
    END
  END inst[14]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END inst[15]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END inst[16]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END inst[17]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END inst[18]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END inst[19]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END inst[1]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END inst[20]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END inst[21]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 0.000 138.320 4.000 ;
    END
  END inst[22]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 4.000 ;
    END
  END inst[23]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END inst[24]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END inst[25]
  PIN inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END inst[26]
  PIN inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END inst[27]
  PIN inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END inst[28]
  PIN inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 4.000 ;
    END
  END inst[29]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 4.000 ;
    END
  END inst[2]
  PIN inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END inst[30]
  PIN inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END inst[31]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END inst[3]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END inst[4]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END inst[5]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END inst[6]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END inst[7]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 4.000 ;
    END
  END inst[8]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 4.000 ;
    END
  END inst[9]
  PIN mem_load_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 596.000 462.000 600.000 ;
    END
  END mem_load_out[0]
  PIN mem_load_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 596.000 394.800 600.000 ;
    END
  END mem_load_out[10]
  PIN mem_load_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 596.000 388.080 600.000 ;
    END
  END mem_load_out[11]
  PIN mem_load_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 596.000 381.360 600.000 ;
    END
  END mem_load_out[12]
  PIN mem_load_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 596.000 374.640 600.000 ;
    END
  END mem_load_out[13]
  PIN mem_load_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 596.000 367.920 600.000 ;
    END
  END mem_load_out[14]
  PIN mem_load_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 596.000 361.200 600.000 ;
    END
  END mem_load_out[15]
  PIN mem_load_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 596.000 354.480 600.000 ;
    END
  END mem_load_out[16]
  PIN mem_load_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 596.000 347.760 600.000 ;
    END
  END mem_load_out[17]
  PIN mem_load_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 596.000 341.040 600.000 ;
    END
  END mem_load_out[18]
  PIN mem_load_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 596.000 334.320 600.000 ;
    END
  END mem_load_out[19]
  PIN mem_load_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 596.000 455.280 600.000 ;
    END
  END mem_load_out[1]
  PIN mem_load_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 596.000 327.600 600.000 ;
    END
  END mem_load_out[20]
  PIN mem_load_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 596.000 320.880 600.000 ;
    END
  END mem_load_out[21]
  PIN mem_load_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 596.000 314.160 600.000 ;
    END
  END mem_load_out[22]
  PIN mem_load_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 596.000 307.440 600.000 ;
    END
  END mem_load_out[23]
  PIN mem_load_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 596.000 300.720 600.000 ;
    END
  END mem_load_out[24]
  PIN mem_load_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 596.000 294.000 600.000 ;
    END
  END mem_load_out[25]
  PIN mem_load_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 596.000 287.280 600.000 ;
    END
  END mem_load_out[26]
  PIN mem_load_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 596.000 280.560 600.000 ;
    END
  END mem_load_out[27]
  PIN mem_load_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 596.000 273.840 600.000 ;
    END
  END mem_load_out[28]
  PIN mem_load_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 596.000 267.120 600.000 ;
    END
  END mem_load_out[29]
  PIN mem_load_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 596.000 448.560 600.000 ;
    END
  END mem_load_out[2]
  PIN mem_load_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 596.000 260.400 600.000 ;
    END
  END mem_load_out[30]
  PIN mem_load_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 596.000 253.680 600.000 ;
    END
  END mem_load_out[31]
  PIN mem_load_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 596.000 441.840 600.000 ;
    END
  END mem_load_out[3]
  PIN mem_load_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 596.000 435.120 600.000 ;
    END
  END mem_load_out[4]
  PIN mem_load_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 596.000 428.400 600.000 ;
    END
  END mem_load_out[5]
  PIN mem_load_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 596.000 421.680 600.000 ;
    END
  END mem_load_out[6]
  PIN mem_load_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 596.000 414.960 600.000 ;
    END
  END mem_load_out[7]
  PIN mem_load_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 596.000 408.240 600.000 ;
    END
  END mem_load_out[8]
  PIN mem_load_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 596.000 401.520 600.000 ;
    END
  END mem_load_out[9]
  PIN pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END pc[0]
  PIN pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END pc[10]
  PIN pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 0.000 232.400 4.000 ;
    END
  END pc[11]
  PIN pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 4.000 ;
    END
  END pc[12]
  PIN pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 4.000 ;
    END
  END pc[13]
  PIN pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END pc[14]
  PIN pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END pc[15]
  PIN pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 0.000 254.800 4.000 ;
    END
  END pc[16]
  PIN pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END pc[17]
  PIN pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END pc[18]
  PIN pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END pc[19]
  PIN pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END pc[1]
  PIN pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 0.000 272.720 4.000 ;
    END
  END pc[20]
  PIN pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 4.000 ;
    END
  END pc[21]
  PIN pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 4.000 ;
    END
  END pc[22]
  PIN pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END pc[23]
  PIN pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END pc[24]
  PIN pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 0.000 295.120 4.000 ;
    END
  END pc[25]
  PIN pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 4.000 ;
    END
  END pc[26]
  PIN pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 0.000 304.080 4.000 ;
    END
  END pc[27]
  PIN pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END pc[28]
  PIN pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END pc[29]
  PIN pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END pc[2]
  PIN pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END pc[30]
  PIN pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 4.000 ;
    END
  END pc[31]
  PIN pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END pc[3]
  PIN pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 4.000 ;
    END
  END pc[4]
  PIN pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END pc[5]
  PIN pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 4.000 ;
    END
  END pc[6]
  PIN pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END pc[7]
  PIN pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END pc[8]
  PIN pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END pc[9]
  PIN pc_next[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 0.000 326.480 4.000 ;
    END
  END pc_next[0]
  PIN pc_next[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 0.000 371.280 4.000 ;
    END
  END pc_next[10]
  PIN pc_next[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END pc_next[11]
  PIN pc_next[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 0.000 380.240 4.000 ;
    END
  END pc_next[12]
  PIN pc_next[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 0.000 384.720 4.000 ;
    END
  END pc_next[13]
  PIN pc_next[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 0.000 389.200 4.000 ;
    END
  END pc_next[14]
  PIN pc_next[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 0.000 393.680 4.000 ;
    END
  END pc_next[15]
  PIN pc_next[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END pc_next[16]
  PIN pc_next[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END pc_next[17]
  PIN pc_next[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END pc_next[18]
  PIN pc_next[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END pc_next[19]
  PIN pc_next[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END pc_next[1]
  PIN pc_next[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 0.000 416.080 4.000 ;
    END
  END pc_next[20]
  PIN pc_next[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 0.000 420.560 4.000 ;
    END
  END pc_next[21]
  PIN pc_next[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END pc_next[22]
  PIN pc_next[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END pc_next[23]
  PIN pc_next[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 0.000 434.000 4.000 ;
    END
  END pc_next[24]
  PIN pc_next[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END pc_next[25]
  PIN pc_next[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 0.000 442.960 4.000 ;
    END
  END pc_next[26]
  PIN pc_next[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END pc_next[27]
  PIN pc_next[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END pc_next[28]
  PIN pc_next[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 0.000 456.400 4.000 ;
    END
  END pc_next[29]
  PIN pc_next[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 0.000 335.440 4.000 ;
    END
  END pc_next[2]
  PIN pc_next[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 0.000 460.880 4.000 ;
    END
  END pc_next[30]
  PIN pc_next[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END pc_next[31]
  PIN pc_next[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 0.000 339.920 4.000 ;
    END
  END pc_next[3]
  PIN pc_next[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END pc_next[4]
  PIN pc_next[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END pc_next[5]
  PIN pc_next[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END pc_next[6]
  PIN pc_next[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END pc_next[7]
  PIN pc_next[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 0.000 362.320 4.000 ;
    END
  END pc_next[8]
  PIN pc_next[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END pc_next[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 495.510 585.610 ;
      LAYER Metal2 ;
        RECT 5.180 595.700 37.780 596.820 ;
        RECT 38.940 595.700 44.500 596.820 ;
        RECT 45.660 595.700 51.220 596.820 ;
        RECT 52.380 595.700 57.940 596.820 ;
        RECT 59.100 595.700 64.660 596.820 ;
        RECT 65.820 595.700 71.380 596.820 ;
        RECT 72.540 595.700 78.100 596.820 ;
        RECT 79.260 595.700 84.820 596.820 ;
        RECT 85.980 595.700 91.540 596.820 ;
        RECT 92.700 595.700 98.260 596.820 ;
        RECT 99.420 595.700 104.980 596.820 ;
        RECT 106.140 595.700 111.700 596.820 ;
        RECT 112.860 595.700 118.420 596.820 ;
        RECT 119.580 595.700 125.140 596.820 ;
        RECT 126.300 595.700 131.860 596.820 ;
        RECT 133.020 595.700 138.580 596.820 ;
        RECT 139.740 595.700 145.300 596.820 ;
        RECT 146.460 595.700 152.020 596.820 ;
        RECT 153.180 595.700 158.740 596.820 ;
        RECT 159.900 595.700 165.460 596.820 ;
        RECT 166.620 595.700 172.180 596.820 ;
        RECT 173.340 595.700 178.900 596.820 ;
        RECT 180.060 595.700 185.620 596.820 ;
        RECT 186.780 595.700 192.340 596.820 ;
        RECT 193.500 595.700 199.060 596.820 ;
        RECT 200.220 595.700 205.780 596.820 ;
        RECT 206.940 595.700 212.500 596.820 ;
        RECT 213.660 595.700 219.220 596.820 ;
        RECT 220.380 595.700 225.940 596.820 ;
        RECT 227.100 595.700 232.660 596.820 ;
        RECT 233.820 595.700 239.380 596.820 ;
        RECT 240.540 595.700 246.100 596.820 ;
        RECT 247.260 595.700 252.820 596.820 ;
        RECT 253.980 595.700 259.540 596.820 ;
        RECT 260.700 595.700 266.260 596.820 ;
        RECT 267.420 595.700 272.980 596.820 ;
        RECT 274.140 595.700 279.700 596.820 ;
        RECT 280.860 595.700 286.420 596.820 ;
        RECT 287.580 595.700 293.140 596.820 ;
        RECT 294.300 595.700 299.860 596.820 ;
        RECT 301.020 595.700 306.580 596.820 ;
        RECT 307.740 595.700 313.300 596.820 ;
        RECT 314.460 595.700 320.020 596.820 ;
        RECT 321.180 595.700 326.740 596.820 ;
        RECT 327.900 595.700 333.460 596.820 ;
        RECT 334.620 595.700 340.180 596.820 ;
        RECT 341.340 595.700 346.900 596.820 ;
        RECT 348.060 595.700 353.620 596.820 ;
        RECT 354.780 595.700 360.340 596.820 ;
        RECT 361.500 595.700 367.060 596.820 ;
        RECT 368.220 595.700 373.780 596.820 ;
        RECT 374.940 595.700 380.500 596.820 ;
        RECT 381.660 595.700 387.220 596.820 ;
        RECT 388.380 595.700 393.940 596.820 ;
        RECT 395.100 595.700 400.660 596.820 ;
        RECT 401.820 595.700 407.380 596.820 ;
        RECT 408.540 595.700 414.100 596.820 ;
        RECT 415.260 595.700 420.820 596.820 ;
        RECT 421.980 595.700 427.540 596.820 ;
        RECT 428.700 595.700 434.260 596.820 ;
        RECT 435.420 595.700 440.980 596.820 ;
        RECT 442.140 595.700 447.700 596.820 ;
        RECT 448.860 595.700 454.420 596.820 ;
        RECT 455.580 595.700 461.140 596.820 ;
        RECT 462.300 595.700 497.700 596.820 ;
        RECT 5.180 4.300 497.700 595.700 ;
        RECT 5.180 2.890 34.420 4.300 ;
        RECT 35.580 2.890 38.900 4.300 ;
        RECT 40.060 2.890 43.380 4.300 ;
        RECT 44.540 2.890 47.860 4.300 ;
        RECT 49.020 2.890 52.340 4.300 ;
        RECT 53.500 2.890 56.820 4.300 ;
        RECT 57.980 2.890 61.300 4.300 ;
        RECT 62.460 2.890 65.780 4.300 ;
        RECT 66.940 2.890 70.260 4.300 ;
        RECT 71.420 2.890 74.740 4.300 ;
        RECT 75.900 2.890 79.220 4.300 ;
        RECT 80.380 2.890 83.700 4.300 ;
        RECT 84.860 2.890 88.180 4.300 ;
        RECT 89.340 2.890 92.660 4.300 ;
        RECT 93.820 2.890 97.140 4.300 ;
        RECT 98.300 2.890 101.620 4.300 ;
        RECT 102.780 2.890 106.100 4.300 ;
        RECT 107.260 2.890 110.580 4.300 ;
        RECT 111.740 2.890 115.060 4.300 ;
        RECT 116.220 2.890 119.540 4.300 ;
        RECT 120.700 2.890 124.020 4.300 ;
        RECT 125.180 2.890 128.500 4.300 ;
        RECT 129.660 2.890 132.980 4.300 ;
        RECT 134.140 2.890 137.460 4.300 ;
        RECT 138.620 2.890 141.940 4.300 ;
        RECT 143.100 2.890 146.420 4.300 ;
        RECT 147.580 2.890 150.900 4.300 ;
        RECT 152.060 2.890 155.380 4.300 ;
        RECT 156.540 2.890 159.860 4.300 ;
        RECT 161.020 2.890 164.340 4.300 ;
        RECT 165.500 2.890 168.820 4.300 ;
        RECT 169.980 2.890 173.300 4.300 ;
        RECT 174.460 2.890 177.780 4.300 ;
        RECT 178.940 2.890 182.260 4.300 ;
        RECT 183.420 2.890 186.740 4.300 ;
        RECT 187.900 2.890 191.220 4.300 ;
        RECT 192.380 2.890 195.700 4.300 ;
        RECT 196.860 2.890 200.180 4.300 ;
        RECT 201.340 2.890 204.660 4.300 ;
        RECT 205.820 2.890 209.140 4.300 ;
        RECT 210.300 2.890 213.620 4.300 ;
        RECT 214.780 2.890 218.100 4.300 ;
        RECT 219.260 2.890 222.580 4.300 ;
        RECT 223.740 2.890 227.060 4.300 ;
        RECT 228.220 2.890 231.540 4.300 ;
        RECT 232.700 2.890 236.020 4.300 ;
        RECT 237.180 2.890 240.500 4.300 ;
        RECT 241.660 2.890 244.980 4.300 ;
        RECT 246.140 2.890 249.460 4.300 ;
        RECT 250.620 2.890 253.940 4.300 ;
        RECT 255.100 2.890 258.420 4.300 ;
        RECT 259.580 2.890 262.900 4.300 ;
        RECT 264.060 2.890 267.380 4.300 ;
        RECT 268.540 2.890 271.860 4.300 ;
        RECT 273.020 2.890 276.340 4.300 ;
        RECT 277.500 2.890 280.820 4.300 ;
        RECT 281.980 2.890 285.300 4.300 ;
        RECT 286.460 2.890 289.780 4.300 ;
        RECT 290.940 2.890 294.260 4.300 ;
        RECT 295.420 2.890 298.740 4.300 ;
        RECT 299.900 2.890 303.220 4.300 ;
        RECT 304.380 2.890 307.700 4.300 ;
        RECT 308.860 2.890 312.180 4.300 ;
        RECT 313.340 2.890 316.660 4.300 ;
        RECT 317.820 2.890 321.140 4.300 ;
        RECT 322.300 2.890 325.620 4.300 ;
        RECT 326.780 2.890 330.100 4.300 ;
        RECT 331.260 2.890 334.580 4.300 ;
        RECT 335.740 2.890 339.060 4.300 ;
        RECT 340.220 2.890 343.540 4.300 ;
        RECT 344.700 2.890 348.020 4.300 ;
        RECT 349.180 2.890 352.500 4.300 ;
        RECT 353.660 2.890 356.980 4.300 ;
        RECT 358.140 2.890 361.460 4.300 ;
        RECT 362.620 2.890 365.940 4.300 ;
        RECT 367.100 2.890 370.420 4.300 ;
        RECT 371.580 2.890 374.900 4.300 ;
        RECT 376.060 2.890 379.380 4.300 ;
        RECT 380.540 2.890 383.860 4.300 ;
        RECT 385.020 2.890 388.340 4.300 ;
        RECT 389.500 2.890 392.820 4.300 ;
        RECT 393.980 2.890 397.300 4.300 ;
        RECT 398.460 2.890 401.780 4.300 ;
        RECT 402.940 2.890 406.260 4.300 ;
        RECT 407.420 2.890 410.740 4.300 ;
        RECT 411.900 2.890 415.220 4.300 ;
        RECT 416.380 2.890 419.700 4.300 ;
        RECT 420.860 2.890 424.180 4.300 ;
        RECT 425.340 2.890 428.660 4.300 ;
        RECT 429.820 2.890 433.140 4.300 ;
        RECT 434.300 2.890 437.620 4.300 ;
        RECT 438.780 2.890 442.100 4.300 ;
        RECT 443.260 2.890 446.580 4.300 ;
        RECT 447.740 2.890 451.060 4.300 ;
        RECT 452.220 2.890 455.540 4.300 ;
        RECT 456.700 2.890 460.020 4.300 ;
        RECT 461.180 2.890 464.500 4.300 ;
        RECT 465.660 2.890 497.700 4.300 ;
      LAYER Metal3 ;
        RECT 5.130 2.380 497.750 590.100 ;
      LAYER Metal4 ;
        RECT 20.300 584.680 490.420 590.150 ;
        RECT 20.300 15.080 21.940 584.680 ;
        RECT 24.140 15.080 98.740 584.680 ;
        RECT 100.940 15.080 175.540 584.680 ;
        RECT 177.740 15.080 252.340 584.680 ;
        RECT 254.540 15.080 329.140 584.680 ;
        RECT 331.340 15.080 405.940 584.680 ;
        RECT 408.140 15.080 482.740 584.680 ;
        RECT 484.940 15.080 490.420 584.680 ;
        RECT 20.300 2.330 490.420 15.080 ;
  END
END tinyrv
END LIBRARY

