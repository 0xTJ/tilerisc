magic
tech gf180mcuD
magscale 1 5
timestamp 1701106896
<< obsm1 >>
rect 672 1538 249312 398302
<< obsm2 >>
rect 854 1549 249186 398291
<< metal3 >>
rect 0 252000 400 252056
rect 0 245616 400 245672
rect 249600 245616 250000 245672
rect 249600 244944 250000 245000
rect 249600 244608 250000 244664
rect 249600 244272 250000 244328
rect 0 243936 400 243992
rect 249600 243936 250000 243992
rect 249600 243600 250000 243656
rect 0 243264 400 243320
rect 0 242928 400 242984
rect 0 241584 400 241640
rect 0 240576 400 240632
rect 249600 240240 250000 240296
rect 0 239904 400 239960
rect 249600 239904 250000 239960
rect 249600 239568 250000 239624
rect 0 239232 400 239288
rect 0 238224 400 238280
rect 0 237888 400 237944
rect 249600 237552 250000 237608
rect 0 235200 400 235256
rect 0 234864 400 234920
rect 0 231504 400 231560
rect 249600 230832 250000 230888
rect 249600 230496 250000 230552
rect 0 229824 400 229880
rect 0 229488 400 229544
rect 0 229152 400 229208
rect 0 228816 400 228872
rect 0 226128 400 226184
rect 249600 225792 250000 225848
rect 249600 225120 250000 225176
rect 249600 224448 250000 224504
rect 249600 224112 250000 224168
rect 0 220416 400 220472
rect 0 220080 400 220136
rect 249600 220080 250000 220136
rect 0 218400 400 218456
rect 0 218064 400 218120
rect 249600 217728 250000 217784
rect 249600 216720 250000 216776
rect 0 216384 400 216440
rect 0 215712 400 215768
rect 249600 215712 250000 215768
rect 0 214032 400 214088
rect 0 211680 400 211736
rect 249600 211680 250000 211736
rect 0 211344 400 211400
rect 0 211008 400 211064
rect 0 210672 400 210728
rect 0 210336 400 210392
rect 249600 210336 250000 210392
rect 0 210000 400 210056
rect 0 209664 400 209720
rect 0 209328 400 209384
rect 249600 207312 250000 207368
rect 0 206976 400 207032
rect 249600 205632 250000 205688
rect 249600 205296 250000 205352
rect 249600 204288 250000 204344
rect 249600 203616 250000 203672
rect 249600 202944 250000 203000
rect 0 202272 400 202328
rect 249600 202272 250000 202328
rect 0 201936 400 201992
rect 249600 201936 250000 201992
rect 0 201600 400 201656
rect 249600 201600 250000 201656
rect 0 201264 400 201320
rect 0 197904 400 197960
rect 0 197568 400 197624
rect 0 196224 400 196280
rect 249600 196224 250000 196280
rect 0 195888 400 195944
rect 249600 195888 250000 195944
rect 249600 195552 250000 195608
rect 0 195216 400 195272
rect 249600 194544 250000 194600
rect 249600 193200 250000 193256
rect 249600 192864 250000 192920
rect 0 192528 400 192584
rect 249600 192192 250000 192248
rect 249600 191520 250000 191576
rect 0 191184 400 191240
rect 249600 191184 250000 191240
rect 0 189504 400 189560
rect 249600 188160 250000 188216
rect 249600 185136 250000 185192
rect 249600 184800 250000 184856
rect 0 184464 400 184520
rect 0 184128 400 184184
rect 249600 183792 250000 183848
rect 0 183456 400 183512
rect 0 181776 400 181832
rect 249600 181776 250000 181832
rect 0 181440 400 181496
rect 0 181104 400 181160
rect 0 180768 400 180824
rect 0 180432 400 180488
rect 0 180096 400 180152
rect 0 179760 400 179816
rect 0 179424 400 179480
rect 249600 179424 250000 179480
rect 0 179088 400 179144
rect 0 178752 400 178808
rect 0 178416 400 178472
rect 0 178080 400 178136
rect 249600 177744 250000 177800
rect 0 177408 400 177464
rect 0 177072 400 177128
rect 249600 177072 250000 177128
rect 0 176400 400 176456
rect 249600 176064 250000 176120
rect 249600 175728 250000 175784
rect 249600 175392 250000 175448
rect 0 171696 400 171752
rect 249600 170352 250000 170408
rect 0 170016 400 170072
rect 249600 170016 250000 170072
rect 249600 169680 250000 169736
rect 249600 169344 250000 169400
rect 0 169008 400 169064
rect 249600 169008 250000 169064
rect 0 168672 400 168728
rect 0 168336 400 168392
rect 249600 163296 250000 163352
rect 0 162960 400 163016
rect 249600 162960 250000 163016
rect 249600 162624 250000 162680
rect 249600 161952 250000 162008
rect 0 159936 400 159992
rect 0 158592 400 158648
rect 0 157920 400 157976
rect 249600 157584 250000 157640
rect 249600 155232 250000 155288
rect 249600 153888 250000 153944
rect 249600 153552 250000 153608
<< obsm3 >>
rect 400 252086 249600 398286
rect 430 251970 249600 252086
rect 400 245702 249600 251970
rect 430 245586 249570 245702
rect 400 245030 249600 245586
rect 400 244914 249570 245030
rect 400 244694 249600 244914
rect 400 244578 249570 244694
rect 400 244358 249600 244578
rect 400 244242 249570 244358
rect 400 244022 249600 244242
rect 430 243906 249570 244022
rect 400 243686 249600 243906
rect 400 243570 249570 243686
rect 400 243350 249600 243570
rect 430 243234 249600 243350
rect 400 243014 249600 243234
rect 430 242898 249600 243014
rect 400 241670 249600 242898
rect 430 241554 249600 241670
rect 400 240662 249600 241554
rect 430 240546 249600 240662
rect 400 240326 249600 240546
rect 400 240210 249570 240326
rect 400 239990 249600 240210
rect 430 239874 249570 239990
rect 400 239654 249600 239874
rect 400 239538 249570 239654
rect 400 239318 249600 239538
rect 430 239202 249600 239318
rect 400 238310 249600 239202
rect 430 238194 249600 238310
rect 400 237974 249600 238194
rect 430 237858 249600 237974
rect 400 237638 249600 237858
rect 400 237522 249570 237638
rect 400 235286 249600 237522
rect 430 235170 249600 235286
rect 400 234950 249600 235170
rect 430 234834 249600 234950
rect 400 231590 249600 234834
rect 430 231474 249600 231590
rect 400 230918 249600 231474
rect 400 230802 249570 230918
rect 400 230582 249600 230802
rect 400 230466 249570 230582
rect 400 229910 249600 230466
rect 430 229794 249600 229910
rect 400 229574 249600 229794
rect 430 229458 249600 229574
rect 400 229238 249600 229458
rect 430 229122 249600 229238
rect 400 228902 249600 229122
rect 430 228786 249600 228902
rect 400 226214 249600 228786
rect 430 226098 249600 226214
rect 400 225878 249600 226098
rect 400 225762 249570 225878
rect 400 225206 249600 225762
rect 400 225090 249570 225206
rect 400 224534 249600 225090
rect 400 224418 249570 224534
rect 400 224198 249600 224418
rect 400 224082 249570 224198
rect 400 220502 249600 224082
rect 430 220386 249600 220502
rect 400 220166 249600 220386
rect 430 220050 249570 220166
rect 400 218486 249600 220050
rect 430 218370 249600 218486
rect 400 218150 249600 218370
rect 430 218034 249600 218150
rect 400 217814 249600 218034
rect 400 217698 249570 217814
rect 400 216806 249600 217698
rect 400 216690 249570 216806
rect 400 216470 249600 216690
rect 430 216354 249600 216470
rect 400 215798 249600 216354
rect 430 215682 249570 215798
rect 400 214118 249600 215682
rect 430 214002 249600 214118
rect 400 211766 249600 214002
rect 430 211650 249570 211766
rect 400 211430 249600 211650
rect 430 211314 249600 211430
rect 400 211094 249600 211314
rect 430 210978 249600 211094
rect 400 210758 249600 210978
rect 430 210642 249600 210758
rect 400 210422 249600 210642
rect 430 210306 249570 210422
rect 400 210086 249600 210306
rect 430 209970 249600 210086
rect 400 209750 249600 209970
rect 430 209634 249600 209750
rect 400 209414 249600 209634
rect 430 209298 249600 209414
rect 400 207398 249600 209298
rect 400 207282 249570 207398
rect 400 207062 249600 207282
rect 430 206946 249600 207062
rect 400 205718 249600 206946
rect 400 205602 249570 205718
rect 400 205382 249600 205602
rect 400 205266 249570 205382
rect 400 204374 249600 205266
rect 400 204258 249570 204374
rect 400 203702 249600 204258
rect 400 203586 249570 203702
rect 400 203030 249600 203586
rect 400 202914 249570 203030
rect 400 202358 249600 202914
rect 430 202242 249570 202358
rect 400 202022 249600 202242
rect 430 201906 249570 202022
rect 400 201686 249600 201906
rect 430 201570 249570 201686
rect 400 201350 249600 201570
rect 430 201234 249600 201350
rect 400 197990 249600 201234
rect 430 197874 249600 197990
rect 400 197654 249600 197874
rect 430 197538 249600 197654
rect 400 196310 249600 197538
rect 430 196194 249570 196310
rect 400 195974 249600 196194
rect 430 195858 249570 195974
rect 400 195638 249600 195858
rect 400 195522 249570 195638
rect 400 195302 249600 195522
rect 430 195186 249600 195302
rect 400 194630 249600 195186
rect 400 194514 249570 194630
rect 400 193286 249600 194514
rect 400 193170 249570 193286
rect 400 192950 249600 193170
rect 400 192834 249570 192950
rect 400 192614 249600 192834
rect 430 192498 249600 192614
rect 400 192278 249600 192498
rect 400 192162 249570 192278
rect 400 191606 249600 192162
rect 400 191490 249570 191606
rect 400 191270 249600 191490
rect 430 191154 249570 191270
rect 400 189590 249600 191154
rect 430 189474 249600 189590
rect 400 188246 249600 189474
rect 400 188130 249570 188246
rect 400 185222 249600 188130
rect 400 185106 249570 185222
rect 400 184886 249600 185106
rect 400 184770 249570 184886
rect 400 184550 249600 184770
rect 430 184434 249600 184550
rect 400 184214 249600 184434
rect 430 184098 249600 184214
rect 400 183878 249600 184098
rect 400 183762 249570 183878
rect 400 183542 249600 183762
rect 430 183426 249600 183542
rect 400 181862 249600 183426
rect 430 181746 249570 181862
rect 400 181526 249600 181746
rect 430 181410 249600 181526
rect 400 181190 249600 181410
rect 430 181074 249600 181190
rect 400 180854 249600 181074
rect 430 180738 249600 180854
rect 400 180518 249600 180738
rect 430 180402 249600 180518
rect 400 180182 249600 180402
rect 430 180066 249600 180182
rect 400 179846 249600 180066
rect 430 179730 249600 179846
rect 400 179510 249600 179730
rect 430 179394 249570 179510
rect 400 179174 249600 179394
rect 430 179058 249600 179174
rect 400 178838 249600 179058
rect 430 178722 249600 178838
rect 400 178502 249600 178722
rect 430 178386 249600 178502
rect 400 178166 249600 178386
rect 430 178050 249600 178166
rect 400 177830 249600 178050
rect 400 177714 249570 177830
rect 400 177494 249600 177714
rect 430 177378 249600 177494
rect 400 177158 249600 177378
rect 430 177042 249570 177158
rect 400 176486 249600 177042
rect 430 176370 249600 176486
rect 400 176150 249600 176370
rect 400 176034 249570 176150
rect 400 175814 249600 176034
rect 400 175698 249570 175814
rect 400 175478 249600 175698
rect 400 175362 249570 175478
rect 400 171782 249600 175362
rect 430 171666 249600 171782
rect 400 170438 249600 171666
rect 400 170322 249570 170438
rect 400 170102 249600 170322
rect 430 169986 249570 170102
rect 400 169766 249600 169986
rect 400 169650 249570 169766
rect 400 169430 249600 169650
rect 400 169314 249570 169430
rect 400 169094 249600 169314
rect 430 168978 249570 169094
rect 400 168758 249600 168978
rect 430 168642 249600 168758
rect 400 168422 249600 168642
rect 430 168306 249600 168422
rect 400 163382 249600 168306
rect 400 163266 249570 163382
rect 400 163046 249600 163266
rect 430 162930 249570 163046
rect 400 162710 249600 162930
rect 400 162594 249570 162710
rect 400 162038 249600 162594
rect 400 161922 249570 162038
rect 400 160022 249600 161922
rect 430 159906 249600 160022
rect 400 158678 249600 159906
rect 430 158562 249600 158678
rect 400 158006 249600 158562
rect 430 157890 249600 158006
rect 400 157670 249600 157890
rect 400 157554 249570 157670
rect 400 155318 249600 157554
rect 400 155202 249570 155318
rect 400 153974 249600 155202
rect 400 153858 249570 153974
rect 400 153638 249600 153858
rect 400 153522 249570 153638
rect 400 1554 249600 153522
<< metal4 >>
rect 2224 1538 2384 398302
rect 9904 1538 10064 398302
rect 17584 1538 17744 398302
rect 25264 1538 25424 398302
rect 32944 1538 33104 398302
rect 40624 1538 40784 398302
rect 48304 1538 48464 398302
rect 55984 1538 56144 398302
rect 63664 1538 63824 398302
rect 71344 1538 71504 398302
rect 79024 1538 79184 398302
rect 86704 1538 86864 398302
rect 94384 1538 94544 398302
rect 102064 1538 102224 398302
rect 109744 1538 109904 398302
rect 117424 1538 117584 398302
rect 125104 1538 125264 398302
rect 132784 1538 132944 398302
rect 140464 1538 140624 398302
rect 148144 1538 148304 398302
rect 155824 1538 155984 398302
rect 163504 1538 163664 398302
rect 171184 1538 171344 398302
rect 178864 1538 179024 398302
rect 186544 1538 186704 398302
rect 194224 1538 194384 398302
rect 201904 1538 202064 398302
rect 209584 1538 209744 398302
rect 217264 1538 217424 398302
rect 224944 1538 225104 398302
rect 232624 1538 232784 398302
rect 240304 1538 240464 398302
rect 247984 1538 248144 398302
<< obsm4 >>
rect 100926 150761 102034 252159
rect 102254 150761 109714 252159
rect 109934 150761 117394 252159
rect 117614 150761 125074 252159
rect 125294 150761 132754 252159
rect 132974 150761 140434 252159
rect 140654 150761 148114 252159
rect 148334 150761 149282 252159
<< labels >>
rlabel metal3 s 0 195216 400 195272 6 ack
port 1 nsew signal output
rlabel metal3 s 0 252000 400 252056 6 clk
port 2 nsew signal input
rlabel metal3 s 0 197568 400 197624 6 cyc
port 3 nsew signal input
rlabel metal3 s 249600 245616 250000 245672 6 dat_in[0]
port 4 nsew signal input
rlabel metal3 s 249600 157584 250000 157640 6 dat_in[10]
port 5 nsew signal input
rlabel metal3 s 249600 155232 250000 155288 6 dat_in[11]
port 6 nsew signal input
rlabel metal3 s 249600 163296 250000 163352 6 dat_in[12]
port 7 nsew signal input
rlabel metal3 s 249600 161952 250000 162008 6 dat_in[13]
port 8 nsew signal input
rlabel metal3 s 249600 162960 250000 163016 6 dat_in[14]
port 9 nsew signal input
rlabel metal3 s 249600 162624 250000 162680 6 dat_in[15]
port 10 nsew signal input
rlabel metal3 s 0 235200 400 235256 6 dat_in[16]
port 11 nsew signal input
rlabel metal3 s 249600 230496 250000 230552 6 dat_in[17]
port 12 nsew signal input
rlabel metal3 s 249600 230832 250000 230888 6 dat_in[18]
port 13 nsew signal input
rlabel metal3 s 0 228816 400 228872 6 dat_in[19]
port 14 nsew signal input
rlabel metal3 s 249600 244272 250000 244328 6 dat_in[1]
port 15 nsew signal input
rlabel metal3 s 249600 211680 250000 211736 6 dat_in[20]
port 16 nsew signal input
rlabel metal3 s 249600 210336 250000 210392 6 dat_in[21]
port 17 nsew signal input
rlabel metal3 s 249600 207312 250000 207368 6 dat_in[22]
port 18 nsew signal input
rlabel metal3 s 249600 205632 250000 205688 6 dat_in[23]
port 19 nsew signal input
rlabel metal3 s 249600 181776 250000 181832 6 dat_in[24]
port 20 nsew signal input
rlabel metal3 s 249600 175728 250000 175784 6 dat_in[25]
port 21 nsew signal input
rlabel metal3 s 249600 176064 250000 176120 6 dat_in[26]
port 22 nsew signal input
rlabel metal3 s 249600 175392 250000 175448 6 dat_in[27]
port 23 nsew signal input
rlabel metal3 s 249600 183792 250000 183848 6 dat_in[28]
port 24 nsew signal input
rlabel metal3 s 249600 179424 250000 179480 6 dat_in[29]
port 25 nsew signal input
rlabel metal3 s 249600 243936 250000 243992 6 dat_in[2]
port 26 nsew signal input
rlabel metal3 s 249600 177744 250000 177800 6 dat_in[30]
port 27 nsew signal input
rlabel metal3 s 249600 191184 250000 191240 6 dat_in[31]
port 28 nsew signal input
rlabel metal3 s 0 243936 400 243992 6 dat_in[32]
port 29 nsew signal input
rlabel metal3 s 0 243264 400 243320 6 dat_in[33]
port 30 nsew signal input
rlabel metal3 s 0 242928 400 242984 6 dat_in[34]
port 31 nsew signal input
rlabel metal3 s 0 245616 400 245672 6 dat_in[35]
port 32 nsew signal input
rlabel metal3 s 0 220416 400 220472 6 dat_in[36]
port 33 nsew signal input
rlabel metal3 s 0 220080 400 220136 6 dat_in[37]
port 34 nsew signal input
rlabel metal3 s 0 218064 400 218120 6 dat_in[38]
port 35 nsew signal input
rlabel metal3 s 0 218400 400 218456 6 dat_in[39]
port 36 nsew signal input
rlabel metal3 s 249600 243600 250000 243656 6 dat_in[3]
port 37 nsew signal input
rlabel metal3 s 0 162960 400 163016 6 dat_in[40]
port 38 nsew signal input
rlabel metal3 s 0 159936 400 159992 6 dat_in[41]
port 39 nsew signal input
rlabel metal3 s 0 157920 400 157976 6 dat_in[42]
port 40 nsew signal input
rlabel metal3 s 0 158592 400 158648 6 dat_in[43]
port 41 nsew signal input
rlabel metal3 s 0 171696 400 171752 6 dat_in[44]
port 42 nsew signal input
rlabel metal3 s 0 168672 400 168728 6 dat_in[45]
port 43 nsew signal input
rlabel metal3 s 0 170016 400 170072 6 dat_in[46]
port 44 nsew signal input
rlabel metal3 s 0 168336 400 168392 6 dat_in[47]
port 45 nsew signal input
rlabel metal3 s 0 231504 400 231560 6 dat_in[48]
port 46 nsew signal input
rlabel metal3 s 0 237888 400 237944 6 dat_in[49]
port 47 nsew signal input
rlabel metal3 s 249600 220080 250000 220136 6 dat_in[4]
port 48 nsew signal input
rlabel metal3 s 0 239232 400 239288 6 dat_in[50]
port 49 nsew signal input
rlabel metal3 s 0 234864 400 234920 6 dat_in[51]
port 50 nsew signal input
rlabel metal3 s 0 210672 400 210728 6 dat_in[52]
port 51 nsew signal input
rlabel metal3 s 0 209328 400 209384 6 dat_in[53]
port 52 nsew signal input
rlabel metal3 s 0 211680 400 211736 6 dat_in[54]
port 53 nsew signal input
rlabel metal3 s 0 210336 400 210392 6 dat_in[55]
port 54 nsew signal input
rlabel metal3 s 0 178080 400 178136 6 dat_in[56]
port 55 nsew signal input
rlabel metal3 s 0 177072 400 177128 6 dat_in[57]
port 56 nsew signal input
rlabel metal3 s 0 176400 400 176456 6 dat_in[58]
port 57 nsew signal input
rlabel metal3 s 0 178416 400 178472 6 dat_in[59]
port 58 nsew signal input
rlabel metal3 s 249600 217728 250000 217784 6 dat_in[5]
port 59 nsew signal input
rlabel metal3 s 0 178752 400 178808 6 dat_in[60]
port 60 nsew signal input
rlabel metal3 s 0 179088 400 179144 6 dat_in[61]
port 61 nsew signal input
rlabel metal3 s 0 180768 400 180824 6 dat_in[62]
port 62 nsew signal input
rlabel metal3 s 0 180432 400 180488 6 dat_in[63]
port 63 nsew signal input
rlabel metal3 s 249600 216720 250000 216776 6 dat_in[6]
port 64 nsew signal input
rlabel metal3 s 249600 215712 250000 215768 6 dat_in[7]
port 65 nsew signal input
rlabel metal3 s 249600 153552 250000 153608 6 dat_in[8]
port 66 nsew signal input
rlabel metal3 s 249600 153888 250000 153944 6 dat_in[9]
port 67 nsew signal input
rlabel metal3 s 249600 225120 250000 225176 6 dat_out[0]
port 68 nsew signal output
rlabel metal3 s 249600 169008 250000 169064 6 dat_out[10]
port 69 nsew signal output
rlabel metal3 s 249600 169680 250000 169736 6 dat_out[11]
port 70 nsew signal output
rlabel metal3 s 249600 169344 250000 169400 6 dat_out[12]
port 71 nsew signal output
rlabel metal3 s 249600 170352 250000 170408 6 dat_out[13]
port 72 nsew signal output
rlabel metal3 s 249600 170016 250000 170072 6 dat_out[14]
port 73 nsew signal output
rlabel metal3 s 249600 177072 250000 177128 6 dat_out[15]
port 74 nsew signal output
rlabel metal3 s 0 226128 400 226184 6 dat_out[16]
port 75 nsew signal output
rlabel metal3 s 0 229488 400 229544 6 dat_out[17]
port 76 nsew signal output
rlabel metal3 s 0 229824 400 229880 6 dat_out[18]
port 77 nsew signal output
rlabel metal3 s 0 229152 400 229208 6 dat_out[19]
port 78 nsew signal output
rlabel metal3 s 249600 237552 250000 237608 6 dat_out[1]
port 79 nsew signal output
rlabel metal3 s 0 214032 400 214088 6 dat_out[20]
port 80 nsew signal output
rlabel metal3 s 0 211008 400 211064 6 dat_out[21]
port 81 nsew signal output
rlabel metal3 s 0 209664 400 209720 6 dat_out[22]
port 82 nsew signal output
rlabel metal3 s 0 206976 400 207032 6 dat_out[23]
port 83 nsew signal output
rlabel metal3 s 249600 185136 250000 185192 6 dat_out[24]
port 84 nsew signal output
rlabel metal3 s 0 181776 400 181832 6 dat_out[25]
port 85 nsew signal output
rlabel metal3 s 249600 184800 250000 184856 6 dat_out[26]
port 86 nsew signal output
rlabel metal3 s 0 181104 400 181160 6 dat_out[27]
port 87 nsew signal output
rlabel metal3 s 249600 188160 250000 188216 6 dat_out[28]
port 88 nsew signal output
rlabel metal3 s 0 189504 400 189560 6 dat_out[29]
port 89 nsew signal output
rlabel metal3 s 249600 240240 250000 240296 6 dat_out[2]
port 90 nsew signal output
rlabel metal3 s 0 191184 400 191240 6 dat_out[30]
port 91 nsew signal output
rlabel metal3 s 0 192528 400 192584 6 dat_out[31]
port 92 nsew signal output
rlabel metal3 s 249600 225792 250000 225848 6 dat_out[32]
port 93 nsew signal output
rlabel metal3 s 249600 239568 250000 239624 6 dat_out[33]
port 94 nsew signal output
rlabel metal3 s 249600 244944 250000 245000 6 dat_out[34]
port 95 nsew signal output
rlabel metal3 s 249600 244608 250000 244664 6 dat_out[35]
port 96 nsew signal output
rlabel metal3 s 249600 224448 250000 224504 6 dat_out[36]
port 97 nsew signal output
rlabel metal3 s 249600 203616 250000 203672 6 dat_out[37]
port 98 nsew signal output
rlabel metal3 s 249600 202944 250000 203000 6 dat_out[38]
port 99 nsew signal output
rlabel metal3 s 249600 201936 250000 201992 6 dat_out[39]
port 100 nsew signal output
rlabel metal3 s 249600 239904 250000 239960 6 dat_out[3]
port 101 nsew signal output
rlabel metal3 s 249600 195552 250000 195608 6 dat_out[40]
port 102 nsew signal output
rlabel metal3 s 249600 192864 250000 192920 6 dat_out[41]
port 103 nsew signal output
rlabel metal3 s 249600 191520 250000 191576 6 dat_out[42]
port 104 nsew signal output
rlabel metal3 s 249600 192192 250000 192248 6 dat_out[43]
port 105 nsew signal output
rlabel metal3 s 249600 193200 250000 193256 6 dat_out[44]
port 106 nsew signal output
rlabel metal3 s 249600 194544 250000 194600 6 dat_out[45]
port 107 nsew signal output
rlabel metal3 s 249600 195888 250000 195944 6 dat_out[46]
port 108 nsew signal output
rlabel metal3 s 249600 196224 250000 196280 6 dat_out[47]
port 109 nsew signal output
rlabel metal3 s 0 240576 400 240632 6 dat_out[48]
port 110 nsew signal output
rlabel metal3 s 0 238224 400 238280 6 dat_out[49]
port 111 nsew signal output
rlabel metal3 s 249600 224112 250000 224168 6 dat_out[4]
port 112 nsew signal output
rlabel metal3 s 0 241584 400 241640 6 dat_out[50]
port 113 nsew signal output
rlabel metal3 s 0 239904 400 239960 6 dat_out[51]
port 114 nsew signal output
rlabel metal3 s 0 215712 400 215768 6 dat_out[52]
port 115 nsew signal output
rlabel metal3 s 0 210000 400 210056 6 dat_out[53]
port 116 nsew signal output
rlabel metal3 s 0 216384 400 216440 6 dat_out[54]
port 117 nsew signal output
rlabel metal3 s 0 211344 400 211400 6 dat_out[55]
port 118 nsew signal output
rlabel metal3 s 0 181440 400 181496 6 dat_out[56]
port 119 nsew signal output
rlabel metal3 s 0 179760 400 179816 6 dat_out[57]
port 120 nsew signal output
rlabel metal3 s 0 180096 400 180152 6 dat_out[58]
port 121 nsew signal output
rlabel metal3 s 0 179424 400 179480 6 dat_out[59]
port 122 nsew signal output
rlabel metal3 s 249600 205296 250000 205352 6 dat_out[5]
port 123 nsew signal output
rlabel metal3 s 0 177408 400 177464 6 dat_out[60]
port 124 nsew signal output
rlabel metal3 s 0 184128 400 184184 6 dat_out[61]
port 125 nsew signal output
rlabel metal3 s 0 183456 400 183512 6 dat_out[62]
port 126 nsew signal output
rlabel metal3 s 0 184464 400 184520 6 dat_out[63]
port 127 nsew signal output
rlabel metal3 s 249600 204288 250000 204344 6 dat_out[6]
port 128 nsew signal output
rlabel metal3 s 249600 202272 250000 202328 6 dat_out[7]
port 129 nsew signal output
rlabel metal3 s 249600 201600 250000 201656 6 dat_out[8]
port 130 nsew signal output
rlabel metal3 s 0 169008 400 169064 6 dat_out[9]
port 131 nsew signal output
rlabel metal3 s 0 196224 400 196280 6 mat_idx[0]
port 132 nsew signal input
rlabel metal3 s 0 195888 400 195944 6 mat_idx[1]
port 133 nsew signal input
rlabel metal4 s 2224 1538 2384 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 398302 6 vdd
port 134 nsew power bidirectional
rlabel metal3 s 0 202272 400 202328 6 vector_idx[0]
port 135 nsew signal input
rlabel metal3 s 0 201600 400 201656 6 vector_idx[1]
port 136 nsew signal input
rlabel metal3 s 0 201936 400 201992 6 vector_type[0]
port 137 nsew signal input
rlabel metal3 s 0 201264 400 201320 6 vector_type[1]
port 138 nsew signal input
rlabel metal4 s 9904 1538 10064 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 398302 6 vss
port 139 nsew ground bidirectional
rlabel metal3 s 0 197904 400 197960 6 we
port 140 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 250000 400000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 47553456
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/gpu_core/runs/23_11_27_12_19/results/signoff/gpu_core.magic.gds
string GDS_START 414952
<< end >>

