magic
tech gf180mcuD
magscale 1 10
timestamp 1700139166
<< metal2 >>
rect 3744 55272 3856 55976
rect 3724 55176 3856 55272
rect 4444 55272 4556 55976
rect 5344 55272 5456 55976
rect 4444 55176 4564 55272
rect 5344 55176 5460 55272
rect 13444 55176 13556 55976
rect 14144 55272 14256 55976
rect 14140 55176 14256 55272
rect 14544 55176 14656 55976
rect 14994 55176 15106 55976
rect 15444 55176 15556 55976
rect 16044 55176 16156 55976
rect 24244 55272 24356 55976
rect 24220 55176 24356 55272
rect 25044 55272 25156 55976
rect 25044 55176 25172 55272
rect 25744 55176 25856 55976
rect 30944 55272 31056 55976
rect 30940 55176 31056 55272
rect 31944 55176 32056 55976
rect 32744 55272 32856 55976
rect 32732 55176 32856 55272
rect 33344 55272 33456 55976
rect 33344 55176 33460 55272
rect 36844 55176 36956 55976
rect 46568 55176 46680 55976
rect 52944 55272 53056 55976
rect 52944 55176 53060 55272
rect 54644 55176 54756 55976
rect 56344 55176 56456 55976
rect 59244 55176 59356 55976
rect 63344 55272 63456 55976
rect 63344 55176 63476 55272
rect 63744 55176 63856 55976
rect 64944 55176 65056 55976
rect 73044 55176 73156 55976
rect 73744 55272 73856 55976
rect 73724 55176 73856 55272
rect 74144 55176 74256 55976
rect 74544 55272 74656 55976
rect 74544 55176 74676 55272
rect 74944 55176 75056 55976
rect 75644 55272 75756 55976
rect 75628 55176 75756 55272
rect 83844 55272 83956 55976
rect 83844 55176 83972 55272
rect 84644 55176 84756 55976
rect 85344 55176 85456 55976
rect 3724 54964 3780 55176
rect 3724 54908 3836 54964
rect 3780 54712 3836 54908
rect 4508 54712 4564 55176
rect 5404 54712 5460 55176
rect 13468 54712 13524 55176
rect 14140 54712 14196 55176
rect 14588 54712 14644 55176
rect 15036 54712 15092 55176
rect 15484 54712 15540 55176
rect 16044 54712 16100 55176
rect 24220 54712 24276 55176
rect 25116 54712 25172 55176
rect 25788 54712 25844 55176
rect 30940 54712 30996 55176
rect 31948 54964 32004 55176
rect 31948 54908 32060 54964
rect 32004 54712 32060 54908
rect 32732 54712 32788 55176
rect 33404 54712 33460 55176
rect 36876 54712 36932 55176
rect 46620 54712 46676 55176
rect 53004 54712 53060 55176
rect 54684 54712 54740 55176
rect 56364 54712 56420 55176
rect 59276 54712 59332 55176
rect 63420 54712 63476 55176
rect 63756 54712 63812 55176
rect 64988 54712 65044 55176
rect 73052 54712 73108 55176
rect 73724 54712 73780 55176
rect 74172 54712 74228 55176
rect 74620 54712 74676 55176
rect 74956 54712 75012 55176
rect 75628 54712 75684 55176
rect 83916 54712 83972 55176
rect 84700 54712 84756 55176
rect 85372 54712 85428 55176
<< metal3 >>
rect 1844 52225 2014 52274
rect 1844 52169 1901 52225
rect 1957 52169 2014 52225
rect 1844 52101 2014 52169
rect 1844 52045 1901 52101
rect 1957 52045 2014 52101
rect 1844 51977 2014 52045
rect 1844 51921 1901 51977
rect 1957 51921 2014 51977
rect 1844 51853 2014 51921
rect 1844 51797 1901 51853
rect 1957 51797 2014 51853
rect 1844 51729 2014 51797
rect 1844 51673 1901 51729
rect 1957 51673 2014 51729
rect 1844 51605 2014 51673
rect 1844 51549 1901 51605
rect 1957 51549 2014 51605
rect 1844 51481 2014 51549
rect 1844 51425 1901 51481
rect 1957 51425 2014 51481
rect 1844 51357 2014 51425
rect 1844 51301 1901 51357
rect 1957 51301 2014 51357
rect 1844 51233 2014 51301
rect 1844 51177 1901 51233
rect 1957 51177 2014 51233
rect 1844 51109 2014 51177
rect 1844 51053 1901 51109
rect 1957 51053 2014 51109
rect 1844 51004 2014 51053
rect 86526 52225 86630 52274
rect 86526 52169 86550 52225
rect 86606 52169 86630 52225
rect 86526 52101 86630 52169
rect 86526 52045 86550 52101
rect 86606 52045 86630 52101
rect 86526 51977 86630 52045
rect 86526 51921 86550 51977
rect 86606 51921 86630 51977
rect 86526 51853 86630 51921
rect 86526 51797 86550 51853
rect 86606 51797 86630 51853
rect 86526 51729 86630 51797
rect 86526 51673 86550 51729
rect 86606 51673 86630 51729
rect 86526 51605 86630 51673
rect 86526 51549 86550 51605
rect 86606 51549 86630 51605
rect 86526 51481 86630 51549
rect 86526 51425 86550 51481
rect 86606 51425 86630 51481
rect 86526 51357 86630 51425
rect 86526 51301 86550 51357
rect 86606 51301 86630 51357
rect 86526 51233 86630 51301
rect 86526 51177 86550 51233
rect 86606 51177 86630 51233
rect 86526 51109 86630 51177
rect 86526 51053 86550 51109
rect 86606 51053 86630 51109
rect 86526 51004 86630 51053
rect 86650 52225 87126 52274
rect 86650 52169 86674 52225
rect 86730 52169 86798 52225
rect 86854 52169 86922 52225
rect 86978 52169 87046 52225
rect 87102 52169 87126 52225
rect 86650 52101 87126 52169
rect 86650 52045 86674 52101
rect 86730 52045 86798 52101
rect 86854 52045 86922 52101
rect 86978 52045 87046 52101
rect 87102 52045 87126 52101
rect 86650 51977 87126 52045
rect 86650 51921 86674 51977
rect 86730 51921 86798 51977
rect 86854 51921 86922 51977
rect 86978 51921 87046 51977
rect 87102 51921 87126 51977
rect 86650 51853 87126 51921
rect 86650 51797 86674 51853
rect 86730 51797 86798 51853
rect 86854 51797 86922 51853
rect 86978 51797 87046 51853
rect 87102 51797 87126 51853
rect 86650 51729 87126 51797
rect 86650 51673 86674 51729
rect 86730 51673 86798 51729
rect 86854 51673 86922 51729
rect 86978 51673 87046 51729
rect 87102 51673 87126 51729
rect 86650 51605 87126 51673
rect 86650 51549 86674 51605
rect 86730 51549 86798 51605
rect 86854 51549 86922 51605
rect 86978 51549 87046 51605
rect 87102 51549 87126 51605
rect 86650 51481 87126 51549
rect 86650 51425 86674 51481
rect 86730 51425 86798 51481
rect 86854 51425 86922 51481
rect 86978 51425 87046 51481
rect 87102 51425 87126 51481
rect 86650 51357 87126 51425
rect 86650 51301 86674 51357
rect 86730 51301 86798 51357
rect 86854 51301 86922 51357
rect 86978 51301 87046 51357
rect 87102 51301 87126 51357
rect 86650 51233 87126 51301
rect 86650 51177 86674 51233
rect 86730 51177 86798 51233
rect 86854 51177 86922 51233
rect 86978 51177 87046 51233
rect 87102 51177 87126 51233
rect 86650 51109 87126 51177
rect 86650 51053 86674 51109
rect 86730 51053 86798 51109
rect 86854 51053 86922 51109
rect 86978 51053 87046 51109
rect 87102 51053 87126 51109
rect 86650 51004 87126 51053
rect 86526 48991 86630 49010
rect 86526 48935 86550 48991
rect 86606 48935 86630 48991
rect 86526 48867 86630 48935
rect 86526 48811 86550 48867
rect 86606 48811 86630 48867
rect 86526 48743 86630 48811
rect 86526 48687 86550 48743
rect 86606 48687 86630 48743
rect 86526 48619 86630 48687
rect 86526 48563 86550 48619
rect 86606 48563 86630 48619
rect 86526 48544 86630 48563
rect 86650 48991 87126 49010
rect 86650 48935 86674 48991
rect 86730 48935 86798 48991
rect 86854 48935 86922 48991
rect 86978 48935 87046 48991
rect 87102 48935 87126 48991
rect 86650 48867 87126 48935
rect 86650 48811 86674 48867
rect 86730 48811 86798 48867
rect 86854 48811 86922 48867
rect 86978 48811 87046 48867
rect 87102 48811 87126 48867
rect 86650 48743 87126 48811
rect 86650 48687 86674 48743
rect 86730 48687 86798 48743
rect 86854 48687 86922 48743
rect 86978 48687 87046 48743
rect 87102 48687 87126 48743
rect 86650 48619 87126 48687
rect 86650 48563 86674 48619
rect 86730 48563 86798 48619
rect 86854 48563 86922 48619
rect 86978 48563 87046 48619
rect 87102 48563 87126 48619
rect 86650 48544 87126 48563
rect 86526 48495 86630 48514
rect 86526 48439 86550 48495
rect 86606 48439 86630 48495
rect 86526 48371 86630 48439
rect 86526 48315 86550 48371
rect 86606 48315 86630 48371
rect 86526 48247 86630 48315
rect 86526 48191 86550 48247
rect 86606 48191 86630 48247
rect 86526 48123 86630 48191
rect 86526 48067 86550 48123
rect 86606 48067 86630 48123
rect 86526 48048 86630 48067
rect 86650 48495 87126 48514
rect 86650 48439 86674 48495
rect 86730 48439 86798 48495
rect 86854 48439 86922 48495
rect 86978 48439 87046 48495
rect 87102 48439 87126 48495
rect 86650 48371 87126 48439
rect 86650 48315 86674 48371
rect 86730 48315 86798 48371
rect 86854 48315 86922 48371
rect 86978 48315 87046 48371
rect 87102 48315 87126 48371
rect 86650 48247 87126 48315
rect 86650 48191 86674 48247
rect 86730 48191 86798 48247
rect 86854 48191 86922 48247
rect 86978 48191 87046 48247
rect 87102 48191 87126 48247
rect 86650 48123 87126 48191
rect 86650 48067 86674 48123
rect 86730 48067 86798 48123
rect 86854 48067 86922 48123
rect 86978 48067 87046 48123
rect 87102 48067 87126 48123
rect 86650 48048 87126 48067
rect 86526 47999 86630 48018
rect 86526 47943 86550 47999
rect 86606 47943 86630 47999
rect 86526 47875 86630 47943
rect 86526 47819 86550 47875
rect 86606 47819 86630 47875
rect 86526 47751 86630 47819
rect 1906 47701 2382 47732
rect 1906 47645 1930 47701
rect 1986 47645 2054 47701
rect 2110 47645 2178 47701
rect 2234 47645 2302 47701
rect 2358 47645 2382 47701
rect 1906 47577 2382 47645
rect 1906 47521 1930 47577
rect 1986 47521 2054 47577
rect 2110 47521 2178 47577
rect 2234 47521 2302 47577
rect 2358 47521 2382 47577
rect 86526 47695 86550 47751
rect 86606 47695 86630 47751
rect 86526 47627 86630 47695
rect 86526 47571 86550 47627
rect 86606 47571 86630 47627
rect 86526 47552 86630 47571
rect 86650 47999 87126 48018
rect 86650 47943 86674 47999
rect 86730 47943 86798 47999
rect 86854 47943 86922 47999
rect 86978 47943 87046 47999
rect 87102 47943 87126 47999
rect 86650 47875 87126 47943
rect 86650 47819 86674 47875
rect 86730 47819 86798 47875
rect 86854 47819 86922 47875
rect 86978 47819 87046 47875
rect 87102 47819 87126 47875
rect 86650 47751 87126 47819
rect 86650 47695 86674 47751
rect 86730 47695 86798 47751
rect 86854 47695 86922 47751
rect 86978 47695 87046 47751
rect 87102 47695 87126 47751
rect 86650 47627 87126 47695
rect 86650 47571 86674 47627
rect 86730 47571 86798 47627
rect 86854 47571 86922 47627
rect 86978 47571 87046 47627
rect 87102 47571 87126 47627
rect 86650 47552 87126 47571
rect 1906 47453 2382 47521
rect 1906 47397 1930 47453
rect 1986 47397 2054 47453
rect 2110 47397 2178 47453
rect 2234 47397 2302 47453
rect 2358 47397 2382 47453
rect 1906 47329 2382 47397
rect 1906 47273 1930 47329
rect 1986 47273 2054 47329
rect 2110 47273 2178 47329
rect 2234 47273 2302 47329
rect 2358 47273 2382 47329
rect 1906 47242 2382 47273
rect 86526 47503 86630 47522
rect 86526 47447 86550 47503
rect 86606 47447 86630 47503
rect 86526 47379 86630 47447
rect 86526 47323 86550 47379
rect 86606 47323 86630 47379
rect 86526 47255 86630 47323
rect 86526 47199 86550 47255
rect 86606 47199 86630 47255
rect 86526 47180 86630 47199
rect 86650 47503 87126 47522
rect 86650 47447 86674 47503
rect 86730 47447 86798 47503
rect 86854 47447 86922 47503
rect 86978 47447 87046 47503
rect 87102 47447 87126 47503
rect 86650 47379 87126 47447
rect 86650 47323 86674 47379
rect 86730 47323 86798 47379
rect 86854 47323 86922 47379
rect 86978 47323 87046 47379
rect 87102 47323 87126 47379
rect 86650 47255 87126 47323
rect 86650 47199 86674 47255
rect 86730 47199 86798 47255
rect 86854 47199 86922 47255
rect 86978 47199 87046 47255
rect 87102 47199 87126 47255
rect 86650 47180 87126 47199
rect 1044 42689 1148 42740
rect 1044 42633 1068 42689
rect 1124 42633 1148 42689
rect 1044 42565 1148 42633
rect 1044 42509 1068 42565
rect 1124 42509 1148 42565
rect 1044 42441 1148 42509
rect 1044 42385 1068 42441
rect 1124 42385 1148 42441
rect 1044 42317 1148 42385
rect 1044 42261 1068 42317
rect 1124 42261 1148 42317
rect 1044 42193 1148 42261
rect 1044 42137 1068 42193
rect 1124 42137 1148 42193
rect 1044 42069 1148 42137
rect 1044 42013 1068 42069
rect 1124 42013 1148 42069
rect 1044 41945 1148 42013
rect 1044 41889 1068 41945
rect 1124 41889 1148 41945
rect 1044 41821 1148 41889
rect 1044 41765 1068 41821
rect 1124 41765 1148 41821
rect 1044 41697 1148 41765
rect 1044 41641 1068 41697
rect 1124 41641 1148 41697
rect 1044 41573 1148 41641
rect 1044 41517 1068 41573
rect 1124 41517 1148 41573
rect 1044 41449 1148 41517
rect 1044 41393 1068 41449
rect 1124 41393 1148 41449
rect 1044 41325 1148 41393
rect 1044 41269 1068 41325
rect 1124 41269 1148 41325
rect 1044 41201 1148 41269
rect 1044 41145 1068 41201
rect 1124 41145 1148 41201
rect 1044 41077 1148 41145
rect 1044 41021 1068 41077
rect 1124 41021 1148 41077
rect 1044 40953 1148 41021
rect 1044 40897 1068 40953
rect 1124 40897 1148 40953
rect 1044 40829 1148 40897
rect 1044 40773 1068 40829
rect 1124 40773 1148 40829
rect 1044 40705 1148 40773
rect 1044 40649 1068 40705
rect 1124 40649 1148 40705
rect 1044 40598 1148 40649
rect 1168 42689 1644 42740
rect 1168 42633 1192 42689
rect 1248 42633 1316 42689
rect 1372 42633 1440 42689
rect 1496 42633 1564 42689
rect 1620 42633 1644 42689
rect 1168 42565 1644 42633
rect 1168 42509 1192 42565
rect 1248 42509 1316 42565
rect 1372 42509 1440 42565
rect 1496 42509 1564 42565
rect 1620 42509 1644 42565
rect 1168 42441 1644 42509
rect 1168 42385 1192 42441
rect 1248 42385 1316 42441
rect 1372 42385 1440 42441
rect 1496 42385 1564 42441
rect 1620 42385 1644 42441
rect 1168 42317 1644 42385
rect 1168 42261 1192 42317
rect 1248 42261 1316 42317
rect 1372 42261 1440 42317
rect 1496 42261 1564 42317
rect 1620 42261 1644 42317
rect 1168 42193 1644 42261
rect 1168 42137 1192 42193
rect 1248 42137 1316 42193
rect 1372 42137 1440 42193
rect 1496 42137 1564 42193
rect 1620 42137 1644 42193
rect 1168 42069 1644 42137
rect 1168 42013 1192 42069
rect 1248 42013 1316 42069
rect 1372 42013 1440 42069
rect 1496 42013 1564 42069
rect 1620 42013 1644 42069
rect 1168 41945 1644 42013
rect 1168 41889 1192 41945
rect 1248 41889 1316 41945
rect 1372 41889 1440 41945
rect 1496 41889 1564 41945
rect 1620 41889 1644 41945
rect 1168 41821 1644 41889
rect 1168 41765 1192 41821
rect 1248 41765 1316 41821
rect 1372 41765 1440 41821
rect 1496 41765 1564 41821
rect 1620 41765 1644 41821
rect 1168 41697 1644 41765
rect 1168 41641 1192 41697
rect 1248 41641 1316 41697
rect 1372 41641 1440 41697
rect 1496 41641 1564 41697
rect 1620 41641 1644 41697
rect 1168 41573 1644 41641
rect 1168 41517 1192 41573
rect 1248 41517 1316 41573
rect 1372 41517 1440 41573
rect 1496 41517 1564 41573
rect 1620 41517 1644 41573
rect 1168 41449 1644 41517
rect 1168 41393 1192 41449
rect 1248 41393 1316 41449
rect 1372 41393 1440 41449
rect 1496 41393 1564 41449
rect 1620 41393 1644 41449
rect 1168 41325 1644 41393
rect 1168 41269 1192 41325
rect 1248 41269 1316 41325
rect 1372 41269 1440 41325
rect 1496 41269 1564 41325
rect 1620 41269 1644 41325
rect 1168 41201 1644 41269
rect 1168 41145 1192 41201
rect 1248 41145 1316 41201
rect 1372 41145 1440 41201
rect 1496 41145 1564 41201
rect 1620 41145 1644 41201
rect 1168 41077 1644 41145
rect 1168 41021 1192 41077
rect 1248 41021 1316 41077
rect 1372 41021 1440 41077
rect 1496 41021 1564 41077
rect 1620 41021 1644 41077
rect 1168 40953 1644 41021
rect 1168 40897 1192 40953
rect 1248 40897 1316 40953
rect 1372 40897 1440 40953
rect 1496 40897 1564 40953
rect 1620 40897 1644 40953
rect 1168 40829 1644 40897
rect 1168 40773 1192 40829
rect 1248 40773 1316 40829
rect 1372 40773 1440 40829
rect 1496 40773 1564 40829
rect 1620 40773 1644 40829
rect 1168 40705 1644 40773
rect 1168 40649 1192 40705
rect 1248 40649 1316 40705
rect 1372 40649 1440 40705
rect 1496 40649 1564 40705
rect 1620 40649 1644 40705
rect 1168 40598 1644 40649
rect 85726 42689 85830 42740
rect 85726 42633 85750 42689
rect 85806 42633 85830 42689
rect 85726 42565 85830 42633
rect 85726 42509 85750 42565
rect 85806 42509 85830 42565
rect 85726 42441 85830 42509
rect 85726 42385 85750 42441
rect 85806 42385 85830 42441
rect 85726 42317 85830 42385
rect 85726 42261 85750 42317
rect 85806 42261 85830 42317
rect 85726 42193 85830 42261
rect 85726 42137 85750 42193
rect 85806 42137 85830 42193
rect 85726 42069 85830 42137
rect 85726 42013 85750 42069
rect 85806 42013 85830 42069
rect 85726 41945 85830 42013
rect 85726 41889 85750 41945
rect 85806 41889 85830 41945
rect 85726 41821 85830 41889
rect 85726 41765 85750 41821
rect 85806 41765 85830 41821
rect 85726 41697 85830 41765
rect 85726 41641 85750 41697
rect 85806 41641 85830 41697
rect 85726 41573 85830 41641
rect 85726 41517 85750 41573
rect 85806 41517 85830 41573
rect 85726 41449 85830 41517
rect 85726 41393 85750 41449
rect 85806 41393 85830 41449
rect 85726 41325 85830 41393
rect 85726 41269 85750 41325
rect 85806 41269 85830 41325
rect 85726 41201 85830 41269
rect 85726 41145 85750 41201
rect 85806 41145 85830 41201
rect 85726 41077 85830 41145
rect 85726 41021 85750 41077
rect 85806 41021 85830 41077
rect 85726 40953 85830 41021
rect 85726 40897 85750 40953
rect 85806 40897 85830 40953
rect 85726 40829 85830 40897
rect 85726 40773 85750 40829
rect 85806 40773 85830 40829
rect 85726 40705 85830 40773
rect 85726 40649 85750 40705
rect 85806 40649 85830 40705
rect 85726 40598 85830 40649
rect 85850 42689 86326 42740
rect 85850 42633 85874 42689
rect 85930 42633 85998 42689
rect 86054 42633 86122 42689
rect 86178 42633 86246 42689
rect 86302 42633 86326 42689
rect 85850 42565 86326 42633
rect 85850 42509 85874 42565
rect 85930 42509 85998 42565
rect 86054 42509 86122 42565
rect 86178 42509 86246 42565
rect 86302 42509 86326 42565
rect 85850 42441 86326 42509
rect 85850 42385 85874 42441
rect 85930 42385 85998 42441
rect 86054 42385 86122 42441
rect 86178 42385 86246 42441
rect 86302 42385 86326 42441
rect 85850 42317 86326 42385
rect 85850 42261 85874 42317
rect 85930 42261 85998 42317
rect 86054 42261 86122 42317
rect 86178 42261 86246 42317
rect 86302 42261 86326 42317
rect 85850 42193 86326 42261
rect 85850 42137 85874 42193
rect 85930 42137 85998 42193
rect 86054 42137 86122 42193
rect 86178 42137 86246 42193
rect 86302 42137 86326 42193
rect 85850 42069 86326 42137
rect 85850 42013 85874 42069
rect 85930 42013 85998 42069
rect 86054 42013 86122 42069
rect 86178 42013 86246 42069
rect 86302 42013 86326 42069
rect 85850 41945 86326 42013
rect 85850 41889 85874 41945
rect 85930 41889 85998 41945
rect 86054 41889 86122 41945
rect 86178 41889 86246 41945
rect 86302 41889 86326 41945
rect 85850 41821 86326 41889
rect 85850 41765 85874 41821
rect 85930 41765 85998 41821
rect 86054 41765 86122 41821
rect 86178 41765 86246 41821
rect 86302 41765 86326 41821
rect 85850 41697 86326 41765
rect 85850 41641 85874 41697
rect 85930 41641 85998 41697
rect 86054 41641 86122 41697
rect 86178 41641 86246 41697
rect 86302 41641 86326 41697
rect 85850 41573 86326 41641
rect 85850 41517 85874 41573
rect 85930 41517 85998 41573
rect 86054 41517 86122 41573
rect 86178 41517 86246 41573
rect 86302 41517 86326 41573
rect 85850 41449 86326 41517
rect 85850 41393 85874 41449
rect 85930 41393 85998 41449
rect 86054 41393 86122 41449
rect 86178 41393 86246 41449
rect 86302 41393 86326 41449
rect 85850 41325 86326 41393
rect 85850 41269 85874 41325
rect 85930 41269 85998 41325
rect 86054 41269 86122 41325
rect 86178 41269 86246 41325
rect 86302 41269 86326 41325
rect 85850 41201 86326 41269
rect 85850 41145 85874 41201
rect 85930 41145 85998 41201
rect 86054 41145 86122 41201
rect 86178 41145 86246 41201
rect 86302 41145 86326 41201
rect 85850 41077 86326 41145
rect 85850 41021 85874 41077
rect 85930 41021 85998 41077
rect 86054 41021 86122 41077
rect 86178 41021 86246 41077
rect 86302 41021 86326 41077
rect 85850 40953 86326 41021
rect 85850 40897 85874 40953
rect 85930 40897 85998 40953
rect 86054 40897 86122 40953
rect 86178 40897 86246 40953
rect 86302 40897 86326 40953
rect 85850 40829 86326 40897
rect 85850 40773 85874 40829
rect 85930 40773 85998 40829
rect 86054 40773 86122 40829
rect 86178 40773 86246 40829
rect 86302 40773 86326 40829
rect 85850 40705 86326 40773
rect 85850 40649 85874 40705
rect 85930 40649 85998 40705
rect 86054 40649 86122 40705
rect 86178 40649 86246 40705
rect 86302 40649 86326 40705
rect 85850 40598 86326 40649
rect 1844 40387 1948 40448
rect 1844 40331 1868 40387
rect 1924 40331 1948 40387
rect 1844 40263 1948 40331
rect 1844 40207 1868 40263
rect 1924 40207 1948 40263
rect 1844 40139 1948 40207
rect 1844 40083 1868 40139
rect 1924 40083 1948 40139
rect 1844 40015 1948 40083
rect 1844 39959 1868 40015
rect 1924 39959 1948 40015
rect 1844 39891 1948 39959
rect 1844 39835 1868 39891
rect 1924 39835 1948 39891
rect 1844 39767 1948 39835
rect 1844 39711 1868 39767
rect 1924 39711 1948 39767
rect 1844 39643 1948 39711
rect 1844 39587 1868 39643
rect 1924 39587 1948 39643
rect 1844 39519 1948 39587
rect 1844 39463 1868 39519
rect 1924 39463 1948 39519
rect 1844 39395 1948 39463
rect 1844 39339 1868 39395
rect 1924 39339 1948 39395
rect 1844 39271 1948 39339
rect 1844 39215 1868 39271
rect 1924 39215 1948 39271
rect 1844 39147 1948 39215
rect 1844 39091 1868 39147
rect 1924 39091 1948 39147
rect 1844 39023 1948 39091
rect 1844 38967 1868 39023
rect 1924 38967 1948 39023
rect 1844 38899 1948 38967
rect 1844 38843 1868 38899
rect 1924 38843 1948 38899
rect 1844 38775 1948 38843
rect 1844 38719 1868 38775
rect 1924 38719 1948 38775
rect 1844 38651 1948 38719
rect 1844 38595 1868 38651
rect 1924 38595 1948 38651
rect 1844 38527 1948 38595
rect 1844 38471 1868 38527
rect 1924 38471 1948 38527
rect 1844 38403 1948 38471
rect 1844 38347 1868 38403
rect 1924 38347 1948 38403
rect 1844 38279 1948 38347
rect 1844 38223 1868 38279
rect 1924 38223 1948 38279
rect 1844 38155 1948 38223
rect 1844 38099 1868 38155
rect 1924 38099 1948 38155
rect 1844 38031 1948 38099
rect 1844 37975 1868 38031
rect 1924 37975 1948 38031
rect 1844 37907 1948 37975
rect 1844 37851 1868 37907
rect 1924 37851 1948 37907
rect 1844 37783 1948 37851
rect 1844 37727 1868 37783
rect 1924 37727 1948 37783
rect 1844 37659 1948 37727
rect 1844 37603 1868 37659
rect 1924 37603 1948 37659
rect 1844 37535 1948 37603
rect 1844 37479 1868 37535
rect 1924 37479 1948 37535
rect 1844 37411 1948 37479
rect 1844 37355 1868 37411
rect 1924 37355 1948 37411
rect 1844 37287 1948 37355
rect 1844 37231 1868 37287
rect 1924 37231 1948 37287
rect 1844 37163 1948 37231
rect 1844 37107 1868 37163
rect 1924 37107 1948 37163
rect 1844 37046 1948 37107
rect 1968 40387 2444 40448
rect 1968 40331 1992 40387
rect 2048 40331 2116 40387
rect 2172 40331 2240 40387
rect 2296 40331 2364 40387
rect 2420 40331 2444 40387
rect 1968 40263 2444 40331
rect 1968 40207 1992 40263
rect 2048 40207 2116 40263
rect 2172 40207 2240 40263
rect 2296 40207 2364 40263
rect 2420 40207 2444 40263
rect 1968 40139 2444 40207
rect 1968 40083 1992 40139
rect 2048 40083 2116 40139
rect 2172 40083 2240 40139
rect 2296 40083 2364 40139
rect 2420 40083 2444 40139
rect 1968 40015 2444 40083
rect 1968 39959 1992 40015
rect 2048 39959 2116 40015
rect 2172 39959 2240 40015
rect 2296 39959 2364 40015
rect 2420 39959 2444 40015
rect 1968 39891 2444 39959
rect 1968 39835 1992 39891
rect 2048 39835 2116 39891
rect 2172 39835 2240 39891
rect 2296 39835 2364 39891
rect 2420 39835 2444 39891
rect 1968 39767 2444 39835
rect 1968 39711 1992 39767
rect 2048 39711 2116 39767
rect 2172 39711 2240 39767
rect 2296 39711 2364 39767
rect 2420 39711 2444 39767
rect 1968 39643 2444 39711
rect 1968 39587 1992 39643
rect 2048 39587 2116 39643
rect 2172 39587 2240 39643
rect 2296 39587 2364 39643
rect 2420 39587 2444 39643
rect 1968 39519 2444 39587
rect 1968 39463 1992 39519
rect 2048 39463 2116 39519
rect 2172 39463 2240 39519
rect 2296 39463 2364 39519
rect 2420 39463 2444 39519
rect 1968 39395 2444 39463
rect 1968 39339 1992 39395
rect 2048 39339 2116 39395
rect 2172 39339 2240 39395
rect 2296 39339 2364 39395
rect 2420 39339 2444 39395
rect 1968 39271 2444 39339
rect 1968 39215 1992 39271
rect 2048 39215 2116 39271
rect 2172 39215 2240 39271
rect 2296 39215 2364 39271
rect 2420 39215 2444 39271
rect 1968 39147 2444 39215
rect 1968 39091 1992 39147
rect 2048 39091 2116 39147
rect 2172 39091 2240 39147
rect 2296 39091 2364 39147
rect 2420 39091 2444 39147
rect 1968 39023 2444 39091
rect 1968 38967 1992 39023
rect 2048 38967 2116 39023
rect 2172 38967 2240 39023
rect 2296 38967 2364 39023
rect 2420 38967 2444 39023
rect 1968 38899 2444 38967
rect 1968 38843 1992 38899
rect 2048 38843 2116 38899
rect 2172 38843 2240 38899
rect 2296 38843 2364 38899
rect 2420 38843 2444 38899
rect 1968 38775 2444 38843
rect 1968 38719 1992 38775
rect 2048 38719 2116 38775
rect 2172 38719 2240 38775
rect 2296 38719 2364 38775
rect 2420 38719 2444 38775
rect 1968 38651 2444 38719
rect 1968 38595 1992 38651
rect 2048 38595 2116 38651
rect 2172 38595 2240 38651
rect 2296 38595 2364 38651
rect 2420 38595 2444 38651
rect 1968 38527 2444 38595
rect 1968 38471 1992 38527
rect 2048 38471 2116 38527
rect 2172 38471 2240 38527
rect 2296 38471 2364 38527
rect 2420 38471 2444 38527
rect 1968 38403 2444 38471
rect 1968 38347 1992 38403
rect 2048 38347 2116 38403
rect 2172 38347 2240 38403
rect 2296 38347 2364 38403
rect 2420 38347 2444 38403
rect 1968 38279 2444 38347
rect 1968 38223 1992 38279
rect 2048 38223 2116 38279
rect 2172 38223 2240 38279
rect 2296 38223 2364 38279
rect 2420 38223 2444 38279
rect 1968 38155 2444 38223
rect 1968 38099 1992 38155
rect 2048 38099 2116 38155
rect 2172 38099 2240 38155
rect 2296 38099 2364 38155
rect 2420 38099 2444 38155
rect 1968 38031 2444 38099
rect 1968 37975 1992 38031
rect 2048 37975 2116 38031
rect 2172 37975 2240 38031
rect 2296 37975 2364 38031
rect 2420 37975 2444 38031
rect 1968 37907 2444 37975
rect 1968 37851 1992 37907
rect 2048 37851 2116 37907
rect 2172 37851 2240 37907
rect 2296 37851 2364 37907
rect 2420 37851 2444 37907
rect 1968 37783 2444 37851
rect 1968 37727 1992 37783
rect 2048 37727 2116 37783
rect 2172 37727 2240 37783
rect 2296 37727 2364 37783
rect 2420 37727 2444 37783
rect 1968 37659 2444 37727
rect 1968 37603 1992 37659
rect 2048 37603 2116 37659
rect 2172 37603 2240 37659
rect 2296 37603 2364 37659
rect 2420 37603 2444 37659
rect 1968 37535 2444 37603
rect 1968 37479 1992 37535
rect 2048 37479 2116 37535
rect 2172 37479 2240 37535
rect 2296 37479 2364 37535
rect 2420 37479 2444 37535
rect 1968 37411 2444 37479
rect 1968 37355 1992 37411
rect 2048 37355 2116 37411
rect 2172 37355 2240 37411
rect 2296 37355 2364 37411
rect 2420 37355 2444 37411
rect 1968 37287 2444 37355
rect 1968 37231 1992 37287
rect 2048 37231 2116 37287
rect 2172 37231 2240 37287
rect 2296 37231 2364 37287
rect 2420 37231 2444 37287
rect 1968 37163 2444 37231
rect 1968 37107 1992 37163
rect 2048 37107 2116 37163
rect 2172 37107 2240 37163
rect 2296 37107 2364 37163
rect 2420 37107 2444 37163
rect 1968 37046 2444 37107
rect 86526 40387 86630 40448
rect 86526 40331 86550 40387
rect 86606 40331 86630 40387
rect 86526 40263 86630 40331
rect 86526 40207 86550 40263
rect 86606 40207 86630 40263
rect 86526 40139 86630 40207
rect 86526 40083 86550 40139
rect 86606 40083 86630 40139
rect 86526 40015 86630 40083
rect 86526 39959 86550 40015
rect 86606 39959 86630 40015
rect 86526 39891 86630 39959
rect 86526 39835 86550 39891
rect 86606 39835 86630 39891
rect 86526 39767 86630 39835
rect 86526 39711 86550 39767
rect 86606 39711 86630 39767
rect 86526 39643 86630 39711
rect 86526 39587 86550 39643
rect 86606 39587 86630 39643
rect 86526 39519 86630 39587
rect 86526 39463 86550 39519
rect 86606 39463 86630 39519
rect 86526 39395 86630 39463
rect 86526 39339 86550 39395
rect 86606 39339 86630 39395
rect 86526 39271 86630 39339
rect 86526 39215 86550 39271
rect 86606 39215 86630 39271
rect 86526 39147 86630 39215
rect 86526 39091 86550 39147
rect 86606 39091 86630 39147
rect 86526 39023 86630 39091
rect 86526 38967 86550 39023
rect 86606 38967 86630 39023
rect 86526 38899 86630 38967
rect 86526 38843 86550 38899
rect 86606 38843 86630 38899
rect 86526 38775 86630 38843
rect 86526 38719 86550 38775
rect 86606 38719 86630 38775
rect 86526 38651 86630 38719
rect 86526 38595 86550 38651
rect 86606 38595 86630 38651
rect 86526 38527 86630 38595
rect 86526 38471 86550 38527
rect 86606 38471 86630 38527
rect 86526 38403 86630 38471
rect 86526 38347 86550 38403
rect 86606 38347 86630 38403
rect 86526 38279 86630 38347
rect 86526 38223 86550 38279
rect 86606 38223 86630 38279
rect 86526 38155 86630 38223
rect 86526 38099 86550 38155
rect 86606 38099 86630 38155
rect 86526 38031 86630 38099
rect 86526 37975 86550 38031
rect 86606 37975 86630 38031
rect 86526 37907 86630 37975
rect 86526 37851 86550 37907
rect 86606 37851 86630 37907
rect 86526 37783 86630 37851
rect 86526 37727 86550 37783
rect 86606 37727 86630 37783
rect 86526 37659 86630 37727
rect 86526 37603 86550 37659
rect 86606 37603 86630 37659
rect 86526 37535 86630 37603
rect 86526 37479 86550 37535
rect 86606 37479 86630 37535
rect 86526 37411 86630 37479
rect 86526 37355 86550 37411
rect 86606 37355 86630 37411
rect 86526 37287 86630 37355
rect 86526 37231 86550 37287
rect 86606 37231 86630 37287
rect 86526 37163 86630 37231
rect 86526 37107 86550 37163
rect 86606 37107 86630 37163
rect 86526 37046 86630 37107
rect 86650 40387 87126 40448
rect 86650 40331 86674 40387
rect 86730 40331 86798 40387
rect 86854 40331 86922 40387
rect 86978 40331 87046 40387
rect 87102 40331 87126 40387
rect 86650 40263 87126 40331
rect 86650 40207 86674 40263
rect 86730 40207 86798 40263
rect 86854 40207 86922 40263
rect 86978 40207 87046 40263
rect 87102 40207 87126 40263
rect 86650 40139 87126 40207
rect 86650 40083 86674 40139
rect 86730 40083 86798 40139
rect 86854 40083 86922 40139
rect 86978 40083 87046 40139
rect 87102 40083 87126 40139
rect 86650 40015 87126 40083
rect 86650 39959 86674 40015
rect 86730 39959 86798 40015
rect 86854 39959 86922 40015
rect 86978 39959 87046 40015
rect 87102 39959 87126 40015
rect 86650 39891 87126 39959
rect 86650 39835 86674 39891
rect 86730 39835 86798 39891
rect 86854 39835 86922 39891
rect 86978 39835 87046 39891
rect 87102 39835 87126 39891
rect 86650 39767 87126 39835
rect 86650 39711 86674 39767
rect 86730 39711 86798 39767
rect 86854 39711 86922 39767
rect 86978 39711 87046 39767
rect 87102 39711 87126 39767
rect 86650 39643 87126 39711
rect 86650 39587 86674 39643
rect 86730 39587 86798 39643
rect 86854 39587 86922 39643
rect 86978 39587 87046 39643
rect 87102 39587 87126 39643
rect 86650 39519 87126 39587
rect 86650 39463 86674 39519
rect 86730 39463 86798 39519
rect 86854 39463 86922 39519
rect 86978 39463 87046 39519
rect 87102 39463 87126 39519
rect 86650 39395 87126 39463
rect 86650 39339 86674 39395
rect 86730 39339 86798 39395
rect 86854 39339 86922 39395
rect 86978 39339 87046 39395
rect 87102 39339 87126 39395
rect 86650 39271 87126 39339
rect 86650 39215 86674 39271
rect 86730 39215 86798 39271
rect 86854 39215 86922 39271
rect 86978 39215 87046 39271
rect 87102 39215 87126 39271
rect 86650 39147 87126 39215
rect 86650 39091 86674 39147
rect 86730 39091 86798 39147
rect 86854 39091 86922 39147
rect 86978 39091 87046 39147
rect 87102 39091 87126 39147
rect 86650 39023 87126 39091
rect 86650 38967 86674 39023
rect 86730 38967 86798 39023
rect 86854 38967 86922 39023
rect 86978 38967 87046 39023
rect 87102 38967 87126 39023
rect 86650 38899 87126 38967
rect 86650 38843 86674 38899
rect 86730 38843 86798 38899
rect 86854 38843 86922 38899
rect 86978 38843 87046 38899
rect 87102 38843 87126 38899
rect 86650 38775 87126 38843
rect 86650 38719 86674 38775
rect 86730 38719 86798 38775
rect 86854 38719 86922 38775
rect 86978 38719 87046 38775
rect 87102 38719 87126 38775
rect 86650 38651 87126 38719
rect 86650 38595 86674 38651
rect 86730 38595 86798 38651
rect 86854 38595 86922 38651
rect 86978 38595 87046 38651
rect 87102 38595 87126 38651
rect 86650 38527 87126 38595
rect 86650 38471 86674 38527
rect 86730 38471 86798 38527
rect 86854 38471 86922 38527
rect 86978 38471 87046 38527
rect 87102 38471 87126 38527
rect 86650 38403 87126 38471
rect 86650 38347 86674 38403
rect 86730 38347 86798 38403
rect 86854 38347 86922 38403
rect 86978 38347 87046 38403
rect 87102 38347 87126 38403
rect 86650 38279 87126 38347
rect 86650 38223 86674 38279
rect 86730 38223 86798 38279
rect 86854 38223 86922 38279
rect 86978 38223 87046 38279
rect 87102 38223 87126 38279
rect 86650 38155 87126 38223
rect 86650 38099 86674 38155
rect 86730 38099 86798 38155
rect 86854 38099 86922 38155
rect 86978 38099 87046 38155
rect 87102 38099 87126 38155
rect 86650 38031 87126 38099
rect 86650 37975 86674 38031
rect 86730 37975 86798 38031
rect 86854 37975 86922 38031
rect 86978 37975 87046 38031
rect 87102 37975 87126 38031
rect 86650 37907 87126 37975
rect 86650 37851 86674 37907
rect 86730 37851 86798 37907
rect 86854 37851 86922 37907
rect 86978 37851 87046 37907
rect 87102 37851 87126 37907
rect 86650 37783 87126 37851
rect 86650 37727 86674 37783
rect 86730 37727 86798 37783
rect 86854 37727 86922 37783
rect 86978 37727 87046 37783
rect 87102 37727 87126 37783
rect 86650 37659 87126 37727
rect 86650 37603 86674 37659
rect 86730 37603 86798 37659
rect 86854 37603 86922 37659
rect 86978 37603 87046 37659
rect 87102 37603 87126 37659
rect 86650 37535 87126 37603
rect 86650 37479 86674 37535
rect 86730 37479 86798 37535
rect 86854 37479 86922 37535
rect 86978 37479 87046 37535
rect 87102 37479 87126 37535
rect 86650 37411 87126 37479
rect 86650 37355 86674 37411
rect 86730 37355 86798 37411
rect 86854 37355 86922 37411
rect 86978 37355 87046 37411
rect 87102 37355 87126 37411
rect 86650 37287 87126 37355
rect 86650 37231 86674 37287
rect 86730 37231 86798 37287
rect 86854 37231 86922 37287
rect 86978 37231 87046 37287
rect 87102 37231 87126 37287
rect 86650 37163 87126 37231
rect 86650 37107 86674 37163
rect 86730 37107 86798 37163
rect 86854 37107 86922 37163
rect 86978 37107 87046 37163
rect 87102 37107 87126 37163
rect 86650 37046 87126 37107
rect 86526 33456 86630 33494
rect 86526 33400 86550 33456
rect 86606 33400 86630 33456
rect 86526 33332 86630 33400
rect 86526 33276 86550 33332
rect 86606 33276 86630 33332
rect 86526 33208 86630 33276
rect 86526 33152 86550 33208
rect 86606 33152 86630 33208
rect 86526 33084 86630 33152
rect 86526 33028 86550 33084
rect 86606 33028 86630 33084
rect 86526 32960 86630 33028
rect 86526 32904 86550 32960
rect 86606 32904 86630 32960
rect 86526 32836 86630 32904
rect 86526 32780 86550 32836
rect 86606 32780 86630 32836
rect 86526 32712 86630 32780
rect 86526 32656 86550 32712
rect 86606 32656 86630 32712
rect 86526 32588 86630 32656
rect 86526 32532 86550 32588
rect 86606 32532 86630 32588
rect 86526 32494 86630 32532
rect 86650 33456 87126 33494
rect 86650 33400 86674 33456
rect 86730 33400 86798 33456
rect 86854 33400 86922 33456
rect 86978 33400 87046 33456
rect 87102 33400 87126 33456
rect 86650 33332 87126 33400
rect 86650 33276 86674 33332
rect 86730 33276 86798 33332
rect 86854 33276 86922 33332
rect 86978 33276 87046 33332
rect 87102 33276 87126 33332
rect 86650 33208 87126 33276
rect 86650 33152 86674 33208
rect 86730 33152 86798 33208
rect 86854 33152 86922 33208
rect 86978 33152 87046 33208
rect 87102 33152 87126 33208
rect 86650 33084 87126 33152
rect 86650 33028 86674 33084
rect 86730 33028 86798 33084
rect 86854 33028 86922 33084
rect 86978 33028 87046 33084
rect 87102 33028 87126 33084
rect 86650 32960 87126 33028
rect 86650 32904 86674 32960
rect 86730 32904 86798 32960
rect 86854 32904 86922 32960
rect 86978 32904 87046 32960
rect 87102 32904 87126 32960
rect 86650 32836 87126 32904
rect 86650 32780 86674 32836
rect 86730 32780 86798 32836
rect 86854 32780 86922 32836
rect 86978 32780 87046 32836
rect 87102 32780 87126 32836
rect 86650 32712 87126 32780
rect 86650 32656 86674 32712
rect 86730 32656 86798 32712
rect 86854 32656 86922 32712
rect 86978 32656 87046 32712
rect 87102 32656 87126 32712
rect 86650 32588 87126 32656
rect 86650 32532 86674 32588
rect 86730 32532 86798 32588
rect 86854 32532 86922 32588
rect 86978 32532 87046 32588
rect 87102 32532 87126 32588
rect 86650 32494 87126 32532
rect 1044 31800 1148 31838
rect 1044 31744 1068 31800
rect 1124 31744 1148 31800
rect 1044 31676 1148 31744
rect 1044 31620 1068 31676
rect 1124 31620 1148 31676
rect 1044 31552 1148 31620
rect 1044 31496 1068 31552
rect 1124 31496 1148 31552
rect 1044 31428 1148 31496
rect 1044 31372 1068 31428
rect 1124 31372 1148 31428
rect 1044 31304 1148 31372
rect 1044 31248 1068 31304
rect 1124 31248 1148 31304
rect 1044 31180 1148 31248
rect 1044 31124 1068 31180
rect 1124 31124 1148 31180
rect 1044 31056 1148 31124
rect 1044 31000 1068 31056
rect 1124 31000 1148 31056
rect 1044 30932 1148 31000
rect 1044 30876 1068 30932
rect 1124 30876 1148 30932
rect 1044 30838 1148 30876
rect 1168 31800 1644 31838
rect 1168 31744 1192 31800
rect 1248 31744 1316 31800
rect 1372 31744 1440 31800
rect 1496 31744 1564 31800
rect 1620 31744 1644 31800
rect 1168 31676 1644 31744
rect 1168 31620 1192 31676
rect 1248 31620 1316 31676
rect 1372 31620 1440 31676
rect 1496 31620 1564 31676
rect 1620 31620 1644 31676
rect 1168 31552 1644 31620
rect 1168 31496 1192 31552
rect 1248 31496 1316 31552
rect 1372 31496 1440 31552
rect 1496 31496 1564 31552
rect 1620 31496 1644 31552
rect 1168 31428 1644 31496
rect 1168 31372 1192 31428
rect 1248 31372 1316 31428
rect 1372 31372 1440 31428
rect 1496 31372 1564 31428
rect 1620 31372 1644 31428
rect 1168 31304 1644 31372
rect 1168 31248 1192 31304
rect 1248 31248 1316 31304
rect 1372 31248 1440 31304
rect 1496 31248 1564 31304
rect 1620 31248 1644 31304
rect 1168 31180 1644 31248
rect 1168 31124 1192 31180
rect 1248 31124 1316 31180
rect 1372 31124 1440 31180
rect 1496 31124 1564 31180
rect 1620 31124 1644 31180
rect 1168 31056 1644 31124
rect 1168 31000 1192 31056
rect 1248 31000 1316 31056
rect 1372 31000 1440 31056
rect 1496 31000 1564 31056
rect 1620 31000 1644 31056
rect 1168 30932 1644 31000
rect 1168 30876 1192 30932
rect 1248 30876 1316 30932
rect 1372 30876 1440 30932
rect 1496 30876 1564 30932
rect 1620 30876 1644 30932
rect 1168 30838 1644 30876
rect 85726 31800 85830 31838
rect 85726 31744 85750 31800
rect 85806 31744 85830 31800
rect 85726 31676 85830 31744
rect 85726 31620 85750 31676
rect 85806 31620 85830 31676
rect 85726 31552 85830 31620
rect 85726 31496 85750 31552
rect 85806 31496 85830 31552
rect 85726 31428 85830 31496
rect 85726 31372 85750 31428
rect 85806 31372 85830 31428
rect 85726 31304 85830 31372
rect 85726 31248 85750 31304
rect 85806 31248 85830 31304
rect 85726 31180 85830 31248
rect 85726 31124 85750 31180
rect 85806 31124 85830 31180
rect 85726 31056 85830 31124
rect 85726 31000 85750 31056
rect 85806 31000 85830 31056
rect 85726 30932 85830 31000
rect 85726 30876 85750 30932
rect 85806 30876 85830 30932
rect 85726 30838 85830 30876
rect 85850 31800 86326 31838
rect 85850 31744 85874 31800
rect 85930 31744 85998 31800
rect 86054 31744 86122 31800
rect 86178 31744 86246 31800
rect 86302 31744 86326 31800
rect 85850 31676 86326 31744
rect 85850 31620 85874 31676
rect 85930 31620 85998 31676
rect 86054 31620 86122 31676
rect 86178 31620 86246 31676
rect 86302 31620 86326 31676
rect 85850 31552 86326 31620
rect 85850 31496 85874 31552
rect 85930 31496 85998 31552
rect 86054 31496 86122 31552
rect 86178 31496 86246 31552
rect 86302 31496 86326 31552
rect 85850 31428 86326 31496
rect 85850 31372 85874 31428
rect 85930 31372 85998 31428
rect 86054 31372 86122 31428
rect 86178 31372 86246 31428
rect 86302 31372 86326 31428
rect 85850 31304 86326 31372
rect 85850 31248 85874 31304
rect 85930 31248 85998 31304
rect 86054 31248 86122 31304
rect 86178 31248 86246 31304
rect 86302 31248 86326 31304
rect 85850 31180 86326 31248
rect 85850 31124 85874 31180
rect 85930 31124 85998 31180
rect 86054 31124 86122 31180
rect 86178 31124 86246 31180
rect 86302 31124 86326 31180
rect 85850 31056 86326 31124
rect 85850 31000 85874 31056
rect 85930 31000 85998 31056
rect 86054 31000 86122 31056
rect 86178 31000 86246 31056
rect 86302 31000 86326 31056
rect 85850 30932 86326 31000
rect 85850 30876 85874 30932
rect 85930 30876 85998 30932
rect 86054 30876 86122 30932
rect 86178 30876 86246 30932
rect 86302 30876 86326 30932
rect 85850 30838 86326 30876
rect 1906 20059 2382 20116
rect 1906 20003 1930 20059
rect 1986 20003 2054 20059
rect 2110 20003 2178 20059
rect 2234 20003 2302 20059
rect 2358 20003 2382 20059
rect 1906 19935 2382 20003
rect 1906 19879 1930 19935
rect 1986 19879 2054 19935
rect 2110 19879 2178 19935
rect 2234 19879 2302 19935
rect 2358 19879 2382 19935
rect 1906 19811 2382 19879
rect 1906 19755 1930 19811
rect 1986 19755 2054 19811
rect 2110 19755 2178 19811
rect 2234 19755 2302 19811
rect 2358 19755 2382 19811
rect 1906 19687 2382 19755
rect 1906 19631 1930 19687
rect 1986 19631 2054 19687
rect 2110 19631 2178 19687
rect 2234 19631 2302 19687
rect 2358 19631 2382 19687
rect 1906 19574 2382 19631
rect 86588 20059 87064 20116
rect 86588 20003 86612 20059
rect 86668 20003 86736 20059
rect 86792 20003 86860 20059
rect 86916 20003 86984 20059
rect 87040 20003 87064 20059
rect 86588 19935 87064 20003
rect 86588 19879 86612 19935
rect 86668 19879 86736 19935
rect 86792 19879 86860 19935
rect 86916 19879 86984 19935
rect 87040 19879 87064 19935
rect 86588 19811 87064 19879
rect 86588 19755 86612 19811
rect 86668 19755 86736 19811
rect 86792 19755 86860 19811
rect 86916 19755 86984 19811
rect 87040 19755 87064 19811
rect 86588 19687 87064 19755
rect 86588 19631 86612 19687
rect 86668 19631 86736 19687
rect 86792 19631 86860 19687
rect 86916 19631 86984 19687
rect 87040 19631 87064 19687
rect 86588 19574 87064 19631
rect 1106 18864 1582 18876
rect 1106 18808 1130 18864
rect 1186 18808 1254 18864
rect 1310 18808 1378 18864
rect 1434 18808 1502 18864
rect 1558 18808 1582 18864
rect 1106 18740 1582 18808
rect 1106 18684 1130 18740
rect 1186 18684 1254 18740
rect 1310 18684 1378 18740
rect 1434 18684 1502 18740
rect 1558 18684 1582 18740
rect 1106 18616 1582 18684
rect 1106 18560 1130 18616
rect 1186 18560 1254 18616
rect 1310 18560 1378 18616
rect 1434 18560 1502 18616
rect 1558 18560 1582 18616
rect 1106 18492 1582 18560
rect 1106 18436 1130 18492
rect 1186 18436 1254 18492
rect 1310 18436 1378 18492
rect 1434 18436 1502 18492
rect 1558 18436 1582 18492
rect 1106 18424 1582 18436
rect 85788 18864 86264 18876
rect 85788 18808 85812 18864
rect 85868 18808 85936 18864
rect 85992 18808 86060 18864
rect 86116 18808 86184 18864
rect 86240 18808 86264 18864
rect 85788 18740 86264 18808
rect 85788 18684 85812 18740
rect 85868 18684 85936 18740
rect 85992 18684 86060 18740
rect 86116 18684 86184 18740
rect 86240 18684 86264 18740
rect 85788 18616 86264 18684
rect 85788 18560 85812 18616
rect 85868 18560 85936 18616
rect 85992 18560 86060 18616
rect 86116 18560 86184 18616
rect 86240 18560 86264 18616
rect 85788 18492 86264 18560
rect 85788 18436 85812 18492
rect 85868 18436 85936 18492
rect 85992 18436 86060 18492
rect 86116 18436 86184 18492
rect 86240 18436 86264 18492
rect 85788 18424 86264 18436
rect 86588 17964 87064 17976
rect 86588 17908 86612 17964
rect 86668 17908 86736 17964
rect 86792 17908 86860 17964
rect 86916 17908 86984 17964
rect 87040 17908 87064 17964
rect 1906 17840 2382 17900
rect 1906 17784 1930 17840
rect 1986 17784 2054 17840
rect 2110 17784 2178 17840
rect 2234 17784 2302 17840
rect 2358 17784 2382 17840
rect 1906 17716 2382 17784
rect 1906 17660 1930 17716
rect 1986 17660 2054 17716
rect 2110 17660 2178 17716
rect 2234 17660 2302 17716
rect 2358 17660 2382 17716
rect 1906 17600 2382 17660
rect 86588 17840 87064 17908
rect 86588 17784 86612 17840
rect 86668 17784 86736 17840
rect 86792 17784 86860 17840
rect 86916 17784 86984 17840
rect 87040 17784 87064 17840
rect 86588 17716 87064 17784
rect 86588 17660 86612 17716
rect 86668 17660 86736 17716
rect 86792 17660 86860 17716
rect 86916 17660 86984 17716
rect 87040 17660 87064 17716
rect 86588 17592 87064 17660
rect 86588 17536 86612 17592
rect 86668 17536 86736 17592
rect 86792 17536 86860 17592
rect 86916 17536 86984 17592
rect 87040 17536 87064 17592
rect 86588 17524 87064 17536
rect 1106 17064 1582 17076
rect 1106 17008 1130 17064
rect 1186 17008 1254 17064
rect 1310 17008 1378 17064
rect 1434 17008 1502 17064
rect 1558 17008 1582 17064
rect 1106 16940 1582 17008
rect 1106 16884 1130 16940
rect 1186 16884 1254 16940
rect 1310 16884 1378 16940
rect 1434 16884 1502 16940
rect 1558 16884 1582 16940
rect 1106 16816 1582 16884
rect 1106 16760 1130 16816
rect 1186 16760 1254 16816
rect 1310 16760 1378 16816
rect 1434 16760 1502 16816
rect 1558 16760 1582 16816
rect 1106 16692 1582 16760
rect 1106 16636 1130 16692
rect 1186 16636 1254 16692
rect 1310 16636 1378 16692
rect 1434 16636 1502 16692
rect 1558 16636 1582 16692
rect 1106 16624 1582 16636
rect 85788 17064 86264 17076
rect 85788 17008 85812 17064
rect 85868 17008 85936 17064
rect 85992 17008 86060 17064
rect 86116 17008 86184 17064
rect 86240 17008 86264 17064
rect 85788 16940 86264 17008
rect 85788 16884 85812 16940
rect 85868 16884 85936 16940
rect 85992 16884 86060 16940
rect 86116 16884 86184 16940
rect 86240 16884 86264 16940
rect 85788 16816 86264 16884
rect 85788 16760 85812 16816
rect 85868 16760 85936 16816
rect 85992 16760 86060 16816
rect 86116 16760 86184 16816
rect 86240 16760 86264 16816
rect 85788 16692 86264 16760
rect 85788 16636 85812 16692
rect 85868 16636 85936 16692
rect 85992 16636 86060 16692
rect 86116 16636 86184 16692
rect 86240 16636 86264 16692
rect 85788 16624 86264 16636
rect 86588 16164 87064 16176
rect 86588 16108 86612 16164
rect 86668 16108 86736 16164
rect 86792 16108 86860 16164
rect 86916 16108 86984 16164
rect 87040 16108 87064 16164
rect 1906 16040 2382 16100
rect 1906 15984 1930 16040
rect 1986 15984 2054 16040
rect 2110 15984 2178 16040
rect 2234 15984 2302 16040
rect 2358 15984 2382 16040
rect 1906 15916 2382 15984
rect 1906 15860 1930 15916
rect 1986 15860 2054 15916
rect 2110 15860 2178 15916
rect 2234 15860 2302 15916
rect 2358 15860 2382 15916
rect 1906 15800 2382 15860
rect 86588 16040 87064 16108
rect 86588 15984 86612 16040
rect 86668 15984 86736 16040
rect 86792 15984 86860 16040
rect 86916 15984 86984 16040
rect 87040 15984 87064 16040
rect 86588 15916 87064 15984
rect 86588 15860 86612 15916
rect 86668 15860 86736 15916
rect 86792 15860 86860 15916
rect 86916 15860 86984 15916
rect 87040 15860 87064 15916
rect 86588 15792 87064 15860
rect 86588 15736 86612 15792
rect 86668 15736 86736 15792
rect 86792 15736 86860 15792
rect 86916 15736 86984 15792
rect 87040 15736 87064 15792
rect 86588 15724 87064 15736
rect 1106 15264 1582 15276
rect 1106 15208 1130 15264
rect 1186 15208 1254 15264
rect 1310 15208 1378 15264
rect 1434 15208 1502 15264
rect 1558 15208 1582 15264
rect 1106 15140 1582 15208
rect 1106 15084 1130 15140
rect 1186 15084 1254 15140
rect 1310 15084 1378 15140
rect 1434 15084 1502 15140
rect 1558 15084 1582 15140
rect 1106 15016 1582 15084
rect 1106 14960 1130 15016
rect 1186 14960 1254 15016
rect 1310 14960 1378 15016
rect 1434 14960 1502 15016
rect 1558 14960 1582 15016
rect 1106 14892 1582 14960
rect 1106 14836 1130 14892
rect 1186 14836 1254 14892
rect 1310 14836 1378 14892
rect 1434 14836 1502 14892
rect 1558 14836 1582 14892
rect 1106 14824 1582 14836
rect 85788 15264 86264 15276
rect 85788 15208 85812 15264
rect 85868 15208 85936 15264
rect 85992 15208 86060 15264
rect 86116 15208 86184 15264
rect 86240 15208 86264 15264
rect 85788 15140 86264 15208
rect 85788 15084 85812 15140
rect 85868 15084 85936 15140
rect 85992 15084 86060 15140
rect 86116 15084 86184 15140
rect 86240 15084 86264 15140
rect 85788 15016 86264 15084
rect 85788 14960 85812 15016
rect 85868 14960 85936 15016
rect 85992 14960 86060 15016
rect 86116 14960 86184 15016
rect 86240 14960 86264 15016
rect 85788 14892 86264 14960
rect 85788 14836 85812 14892
rect 85868 14836 85936 14892
rect 85992 14836 86060 14892
rect 86116 14836 86184 14892
rect 86240 14836 86264 14892
rect 85788 14824 86264 14836
rect 86588 14364 87064 14376
rect 86588 14308 86612 14364
rect 86668 14308 86736 14364
rect 86792 14308 86860 14364
rect 86916 14308 86984 14364
rect 87040 14308 87064 14364
rect 1906 14240 2382 14300
rect 1906 14184 1930 14240
rect 1986 14184 2054 14240
rect 2110 14184 2178 14240
rect 2234 14184 2302 14240
rect 2358 14184 2382 14240
rect 1906 14116 2382 14184
rect 1906 14060 1930 14116
rect 1986 14060 2054 14116
rect 2110 14060 2178 14116
rect 2234 14060 2302 14116
rect 2358 14060 2382 14116
rect 1906 14000 2382 14060
rect 86588 14240 87064 14308
rect 86588 14184 86612 14240
rect 86668 14184 86736 14240
rect 86792 14184 86860 14240
rect 86916 14184 86984 14240
rect 87040 14184 87064 14240
rect 86588 14116 87064 14184
rect 86588 14060 86612 14116
rect 86668 14060 86736 14116
rect 86792 14060 86860 14116
rect 86916 14060 86984 14116
rect 87040 14060 87064 14116
rect 86588 13992 87064 14060
rect 86588 13936 86612 13992
rect 86668 13936 86736 13992
rect 86792 13936 86860 13992
rect 86916 13936 86984 13992
rect 87040 13936 87064 13992
rect 86588 13924 87064 13936
rect 1106 13464 1582 13476
rect 1106 13408 1130 13464
rect 1186 13408 1254 13464
rect 1310 13408 1378 13464
rect 1434 13408 1502 13464
rect 1558 13408 1582 13464
rect 1106 13340 1582 13408
rect 1106 13284 1130 13340
rect 1186 13284 1254 13340
rect 1310 13284 1378 13340
rect 1434 13284 1502 13340
rect 1558 13284 1582 13340
rect 1106 13216 1582 13284
rect 1106 13160 1130 13216
rect 1186 13160 1254 13216
rect 1310 13160 1378 13216
rect 1434 13160 1502 13216
rect 1558 13160 1582 13216
rect 1106 13092 1582 13160
rect 1106 13036 1130 13092
rect 1186 13036 1254 13092
rect 1310 13036 1378 13092
rect 1434 13036 1502 13092
rect 1558 13036 1582 13092
rect 1106 13024 1582 13036
rect 85788 13464 86264 13476
rect 85788 13408 85812 13464
rect 85868 13408 85936 13464
rect 85992 13408 86060 13464
rect 86116 13408 86184 13464
rect 86240 13408 86264 13464
rect 85788 13340 86264 13408
rect 85788 13284 85812 13340
rect 85868 13284 85936 13340
rect 85992 13284 86060 13340
rect 86116 13284 86184 13340
rect 86240 13284 86264 13340
rect 85788 13216 86264 13284
rect 85788 13160 85812 13216
rect 85868 13160 85936 13216
rect 85992 13160 86060 13216
rect 86116 13160 86184 13216
rect 86240 13160 86264 13216
rect 85788 13092 86264 13160
rect 85788 13036 85812 13092
rect 85868 13036 85936 13092
rect 85992 13036 86060 13092
rect 86116 13036 86184 13092
rect 86240 13036 86264 13092
rect 85788 13024 86264 13036
rect 86588 12564 87064 12576
rect 86588 12508 86612 12564
rect 86668 12508 86736 12564
rect 86792 12508 86860 12564
rect 86916 12508 86984 12564
rect 87040 12508 87064 12564
rect 1906 12440 2382 12500
rect 1906 12384 1930 12440
rect 1986 12384 2054 12440
rect 2110 12384 2178 12440
rect 2234 12384 2302 12440
rect 2358 12384 2382 12440
rect 1906 12316 2382 12384
rect 1906 12260 1930 12316
rect 1986 12260 2054 12316
rect 2110 12260 2178 12316
rect 2234 12260 2302 12316
rect 2358 12260 2382 12316
rect 1906 12200 2382 12260
rect 86588 12440 87064 12508
rect 86588 12384 86612 12440
rect 86668 12384 86736 12440
rect 86792 12384 86860 12440
rect 86916 12384 86984 12440
rect 87040 12384 87064 12440
rect 86588 12316 87064 12384
rect 86588 12260 86612 12316
rect 86668 12260 86736 12316
rect 86792 12260 86860 12316
rect 86916 12260 86984 12316
rect 87040 12260 87064 12316
rect 86588 12192 87064 12260
rect 86588 12136 86612 12192
rect 86668 12136 86736 12192
rect 86792 12136 86860 12192
rect 86916 12136 86984 12192
rect 87040 12136 87064 12192
rect 86588 12124 87064 12136
rect 1106 11664 1582 11676
rect 1106 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1582 11664
rect 1106 11540 1582 11608
rect 1106 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1582 11540
rect 1106 11416 1582 11484
rect 1106 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1582 11416
rect 1106 11292 1582 11360
rect 1106 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1582 11292
rect 1106 11224 1582 11236
rect 85788 11664 86264 11676
rect 85788 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86264 11664
rect 85788 11540 86264 11608
rect 85788 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86264 11540
rect 85788 11416 86264 11484
rect 85788 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86264 11416
rect 85788 11292 86264 11360
rect 85788 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86264 11292
rect 85788 11224 86264 11236
rect 86588 10764 87064 10776
rect 86588 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87064 10764
rect 1906 10640 2382 10700
rect 1906 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2382 10640
rect 1906 10516 2382 10584
rect 1906 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2382 10516
rect 1906 10400 2382 10460
rect 86588 10640 87064 10708
rect 86588 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87064 10640
rect 86588 10516 87064 10584
rect 86588 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87064 10516
rect 86588 10392 87064 10460
rect 86588 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87064 10392
rect 86588 10324 87064 10336
rect 1106 9864 1582 9876
rect 1106 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1582 9864
rect 1106 9740 1582 9808
rect 1106 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1582 9740
rect 1106 9616 1582 9684
rect 1106 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1582 9616
rect 1106 9492 1582 9560
rect 1106 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1582 9492
rect 1106 9424 1582 9436
rect 85788 9864 86264 9876
rect 85788 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86264 9864
rect 85788 9740 86264 9808
rect 85788 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86264 9740
rect 85788 9616 86264 9684
rect 85788 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86264 9616
rect 85788 9492 86264 9560
rect 85788 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86264 9492
rect 85788 9424 86264 9436
rect 86588 8964 87064 8976
rect 86588 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87064 8964
rect 1906 8840 2382 8900
rect 1906 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2382 8840
rect 1906 8716 2382 8784
rect 1906 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2382 8716
rect 1906 8600 2382 8660
rect 86588 8840 87064 8908
rect 86588 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87064 8840
rect 86588 8716 87064 8784
rect 86588 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87064 8716
rect 86588 8592 87064 8660
rect 86588 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87064 8592
rect 86588 8524 87064 8536
rect 1106 8064 1582 8076
rect 1106 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1582 8064
rect 1106 7940 1582 8008
rect 1106 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1582 7940
rect 1106 7816 1582 7884
rect 1106 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1582 7816
rect 1106 7692 1582 7760
rect 1106 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1582 7692
rect 1106 7624 1582 7636
rect 85788 8064 86264 8076
rect 85788 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86264 8064
rect 85788 7940 86264 8008
rect 85788 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86264 7940
rect 85788 7816 86264 7884
rect 85788 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86264 7816
rect 85788 7692 86264 7760
rect 85788 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86264 7692
rect 85788 7624 86264 7636
rect 86588 7164 87064 7176
rect 86588 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87064 7164
rect 1906 7040 2382 7100
rect 1906 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2382 7040
rect 1906 6916 2382 6984
rect 1906 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2382 6916
rect 1906 6800 2382 6860
rect 86588 7040 87064 7108
rect 86588 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87064 7040
rect 86588 6916 87064 6984
rect 86588 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87064 6916
rect 86588 6792 87064 6860
rect 86588 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87064 6792
rect 86588 6724 87064 6736
rect 1106 6264 1582 6276
rect 1106 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1582 6264
rect 1106 6140 1582 6208
rect 1106 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1582 6140
rect 1106 6016 1582 6084
rect 1106 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1582 6016
rect 1106 5892 1582 5960
rect 1106 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1582 5892
rect 1106 5824 1582 5836
rect 85788 6264 86264 6276
rect 85788 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86264 6264
rect 85788 6140 86264 6208
rect 85788 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86264 6140
rect 85788 6016 86264 6084
rect 85788 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86264 6016
rect 85788 5892 86264 5960
rect 85788 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86264 5892
rect 85788 5824 86264 5836
rect 86588 5364 87064 5376
rect 86588 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87064 5364
rect 1906 5240 2382 5300
rect 1906 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2382 5240
rect 1906 5116 2382 5184
rect 1906 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2382 5116
rect 1906 5000 2382 5060
rect 86588 5240 87064 5308
rect 86588 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87064 5240
rect 86588 5116 87064 5184
rect 86588 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87064 5116
rect 86588 4992 87064 5060
rect 86588 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87064 4992
rect 86588 4924 87064 4936
rect 1106 4464 1582 4476
rect 1106 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1582 4464
rect 1106 4340 1582 4408
rect 1106 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1582 4340
rect 1106 4216 1582 4284
rect 1106 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1582 4216
rect 1106 4092 1582 4160
rect 1106 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1582 4092
rect 1106 4024 1582 4036
rect 85788 4464 86264 4476
rect 85788 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86264 4464
rect 85788 4340 86264 4408
rect 85788 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86264 4340
rect 85788 4216 86264 4284
rect 85788 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86264 4216
rect 85788 4092 86264 4160
rect 85788 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86264 4092
rect 85788 4024 86264 4036
rect 86588 3632 87064 3700
rect 86588 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87064 3632
rect 86588 3508 87064 3576
rect 1906 3440 2382 3500
rect 1906 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2382 3440
rect 1906 3316 2382 3384
rect 1906 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2382 3316
rect 1906 3200 2382 3260
rect 86588 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87064 3508
rect 86588 3384 87064 3452
rect 86588 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87064 3384
rect 86588 3260 87064 3328
rect 86588 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87064 3260
rect 86588 3136 87064 3204
<< via3 >>
rect 1901 52169 1957 52225
rect 1901 52045 1957 52101
rect 1901 51921 1957 51977
rect 1901 51797 1957 51853
rect 1901 51673 1957 51729
rect 1901 51549 1957 51605
rect 1901 51425 1957 51481
rect 1901 51301 1957 51357
rect 1901 51177 1957 51233
rect 1901 51053 1957 51109
rect 86550 52169 86606 52225
rect 86550 52045 86606 52101
rect 86550 51921 86606 51977
rect 86550 51797 86606 51853
rect 86550 51673 86606 51729
rect 86550 51549 86606 51605
rect 86550 51425 86606 51481
rect 86550 51301 86606 51357
rect 86550 51177 86606 51233
rect 86550 51053 86606 51109
rect 86674 52169 86730 52225
rect 86798 52169 86854 52225
rect 86922 52169 86978 52225
rect 87046 52169 87102 52225
rect 86674 52045 86730 52101
rect 86798 52045 86854 52101
rect 86922 52045 86978 52101
rect 87046 52045 87102 52101
rect 86674 51921 86730 51977
rect 86798 51921 86854 51977
rect 86922 51921 86978 51977
rect 87046 51921 87102 51977
rect 86674 51797 86730 51853
rect 86798 51797 86854 51853
rect 86922 51797 86978 51853
rect 87046 51797 87102 51853
rect 86674 51673 86730 51729
rect 86798 51673 86854 51729
rect 86922 51673 86978 51729
rect 87046 51673 87102 51729
rect 86674 51549 86730 51605
rect 86798 51549 86854 51605
rect 86922 51549 86978 51605
rect 87046 51549 87102 51605
rect 86674 51425 86730 51481
rect 86798 51425 86854 51481
rect 86922 51425 86978 51481
rect 87046 51425 87102 51481
rect 86674 51301 86730 51357
rect 86798 51301 86854 51357
rect 86922 51301 86978 51357
rect 87046 51301 87102 51357
rect 86674 51177 86730 51233
rect 86798 51177 86854 51233
rect 86922 51177 86978 51233
rect 87046 51177 87102 51233
rect 86674 51053 86730 51109
rect 86798 51053 86854 51109
rect 86922 51053 86978 51109
rect 87046 51053 87102 51109
rect 86550 48935 86606 48991
rect 86550 48811 86606 48867
rect 86550 48687 86606 48743
rect 86550 48563 86606 48619
rect 86674 48935 86730 48991
rect 86798 48935 86854 48991
rect 86922 48935 86978 48991
rect 87046 48935 87102 48991
rect 86674 48811 86730 48867
rect 86798 48811 86854 48867
rect 86922 48811 86978 48867
rect 87046 48811 87102 48867
rect 86674 48687 86730 48743
rect 86798 48687 86854 48743
rect 86922 48687 86978 48743
rect 87046 48687 87102 48743
rect 86674 48563 86730 48619
rect 86798 48563 86854 48619
rect 86922 48563 86978 48619
rect 87046 48563 87102 48619
rect 86550 48439 86606 48495
rect 86550 48315 86606 48371
rect 86550 48191 86606 48247
rect 86550 48067 86606 48123
rect 86674 48439 86730 48495
rect 86798 48439 86854 48495
rect 86922 48439 86978 48495
rect 87046 48439 87102 48495
rect 86674 48315 86730 48371
rect 86798 48315 86854 48371
rect 86922 48315 86978 48371
rect 87046 48315 87102 48371
rect 86674 48191 86730 48247
rect 86798 48191 86854 48247
rect 86922 48191 86978 48247
rect 87046 48191 87102 48247
rect 86674 48067 86730 48123
rect 86798 48067 86854 48123
rect 86922 48067 86978 48123
rect 87046 48067 87102 48123
rect 86550 47943 86606 47999
rect 86550 47819 86606 47875
rect 1930 47645 1986 47701
rect 2054 47645 2110 47701
rect 2178 47645 2234 47701
rect 2302 47645 2358 47701
rect 1930 47521 1986 47577
rect 2054 47521 2110 47577
rect 2178 47521 2234 47577
rect 2302 47521 2358 47577
rect 86550 47695 86606 47751
rect 86550 47571 86606 47627
rect 86674 47943 86730 47999
rect 86798 47943 86854 47999
rect 86922 47943 86978 47999
rect 87046 47943 87102 47999
rect 86674 47819 86730 47875
rect 86798 47819 86854 47875
rect 86922 47819 86978 47875
rect 87046 47819 87102 47875
rect 86674 47695 86730 47751
rect 86798 47695 86854 47751
rect 86922 47695 86978 47751
rect 87046 47695 87102 47751
rect 86674 47571 86730 47627
rect 86798 47571 86854 47627
rect 86922 47571 86978 47627
rect 87046 47571 87102 47627
rect 1930 47397 1986 47453
rect 2054 47397 2110 47453
rect 2178 47397 2234 47453
rect 2302 47397 2358 47453
rect 1930 47273 1986 47329
rect 2054 47273 2110 47329
rect 2178 47273 2234 47329
rect 2302 47273 2358 47329
rect 86550 47447 86606 47503
rect 86550 47323 86606 47379
rect 86550 47199 86606 47255
rect 86674 47447 86730 47503
rect 86798 47447 86854 47503
rect 86922 47447 86978 47503
rect 87046 47447 87102 47503
rect 86674 47323 86730 47379
rect 86798 47323 86854 47379
rect 86922 47323 86978 47379
rect 87046 47323 87102 47379
rect 86674 47199 86730 47255
rect 86798 47199 86854 47255
rect 86922 47199 86978 47255
rect 87046 47199 87102 47255
rect 1068 42633 1124 42689
rect 1068 42509 1124 42565
rect 1068 42385 1124 42441
rect 1068 42261 1124 42317
rect 1068 42137 1124 42193
rect 1068 42013 1124 42069
rect 1068 41889 1124 41945
rect 1068 41765 1124 41821
rect 1068 41641 1124 41697
rect 1068 41517 1124 41573
rect 1068 41393 1124 41449
rect 1068 41269 1124 41325
rect 1068 41145 1124 41201
rect 1068 41021 1124 41077
rect 1068 40897 1124 40953
rect 1068 40773 1124 40829
rect 1068 40649 1124 40705
rect 1192 42633 1248 42689
rect 1316 42633 1372 42689
rect 1440 42633 1496 42689
rect 1564 42633 1620 42689
rect 1192 42509 1248 42565
rect 1316 42509 1372 42565
rect 1440 42509 1496 42565
rect 1564 42509 1620 42565
rect 1192 42385 1248 42441
rect 1316 42385 1372 42441
rect 1440 42385 1496 42441
rect 1564 42385 1620 42441
rect 1192 42261 1248 42317
rect 1316 42261 1372 42317
rect 1440 42261 1496 42317
rect 1564 42261 1620 42317
rect 1192 42137 1248 42193
rect 1316 42137 1372 42193
rect 1440 42137 1496 42193
rect 1564 42137 1620 42193
rect 1192 42013 1248 42069
rect 1316 42013 1372 42069
rect 1440 42013 1496 42069
rect 1564 42013 1620 42069
rect 1192 41889 1248 41945
rect 1316 41889 1372 41945
rect 1440 41889 1496 41945
rect 1564 41889 1620 41945
rect 1192 41765 1248 41821
rect 1316 41765 1372 41821
rect 1440 41765 1496 41821
rect 1564 41765 1620 41821
rect 1192 41641 1248 41697
rect 1316 41641 1372 41697
rect 1440 41641 1496 41697
rect 1564 41641 1620 41697
rect 1192 41517 1248 41573
rect 1316 41517 1372 41573
rect 1440 41517 1496 41573
rect 1564 41517 1620 41573
rect 1192 41393 1248 41449
rect 1316 41393 1372 41449
rect 1440 41393 1496 41449
rect 1564 41393 1620 41449
rect 1192 41269 1248 41325
rect 1316 41269 1372 41325
rect 1440 41269 1496 41325
rect 1564 41269 1620 41325
rect 1192 41145 1248 41201
rect 1316 41145 1372 41201
rect 1440 41145 1496 41201
rect 1564 41145 1620 41201
rect 1192 41021 1248 41077
rect 1316 41021 1372 41077
rect 1440 41021 1496 41077
rect 1564 41021 1620 41077
rect 1192 40897 1248 40953
rect 1316 40897 1372 40953
rect 1440 40897 1496 40953
rect 1564 40897 1620 40953
rect 1192 40773 1248 40829
rect 1316 40773 1372 40829
rect 1440 40773 1496 40829
rect 1564 40773 1620 40829
rect 1192 40649 1248 40705
rect 1316 40649 1372 40705
rect 1440 40649 1496 40705
rect 1564 40649 1620 40705
rect 85750 42633 85806 42689
rect 85750 42509 85806 42565
rect 85750 42385 85806 42441
rect 85750 42261 85806 42317
rect 85750 42137 85806 42193
rect 85750 42013 85806 42069
rect 85750 41889 85806 41945
rect 85750 41765 85806 41821
rect 85750 41641 85806 41697
rect 85750 41517 85806 41573
rect 85750 41393 85806 41449
rect 85750 41269 85806 41325
rect 85750 41145 85806 41201
rect 85750 41021 85806 41077
rect 85750 40897 85806 40953
rect 85750 40773 85806 40829
rect 85750 40649 85806 40705
rect 85874 42633 85930 42689
rect 85998 42633 86054 42689
rect 86122 42633 86178 42689
rect 86246 42633 86302 42689
rect 85874 42509 85930 42565
rect 85998 42509 86054 42565
rect 86122 42509 86178 42565
rect 86246 42509 86302 42565
rect 85874 42385 85930 42441
rect 85998 42385 86054 42441
rect 86122 42385 86178 42441
rect 86246 42385 86302 42441
rect 85874 42261 85930 42317
rect 85998 42261 86054 42317
rect 86122 42261 86178 42317
rect 86246 42261 86302 42317
rect 85874 42137 85930 42193
rect 85998 42137 86054 42193
rect 86122 42137 86178 42193
rect 86246 42137 86302 42193
rect 85874 42013 85930 42069
rect 85998 42013 86054 42069
rect 86122 42013 86178 42069
rect 86246 42013 86302 42069
rect 85874 41889 85930 41945
rect 85998 41889 86054 41945
rect 86122 41889 86178 41945
rect 86246 41889 86302 41945
rect 85874 41765 85930 41821
rect 85998 41765 86054 41821
rect 86122 41765 86178 41821
rect 86246 41765 86302 41821
rect 85874 41641 85930 41697
rect 85998 41641 86054 41697
rect 86122 41641 86178 41697
rect 86246 41641 86302 41697
rect 85874 41517 85930 41573
rect 85998 41517 86054 41573
rect 86122 41517 86178 41573
rect 86246 41517 86302 41573
rect 85874 41393 85930 41449
rect 85998 41393 86054 41449
rect 86122 41393 86178 41449
rect 86246 41393 86302 41449
rect 85874 41269 85930 41325
rect 85998 41269 86054 41325
rect 86122 41269 86178 41325
rect 86246 41269 86302 41325
rect 85874 41145 85930 41201
rect 85998 41145 86054 41201
rect 86122 41145 86178 41201
rect 86246 41145 86302 41201
rect 85874 41021 85930 41077
rect 85998 41021 86054 41077
rect 86122 41021 86178 41077
rect 86246 41021 86302 41077
rect 85874 40897 85930 40953
rect 85998 40897 86054 40953
rect 86122 40897 86178 40953
rect 86246 40897 86302 40953
rect 85874 40773 85930 40829
rect 85998 40773 86054 40829
rect 86122 40773 86178 40829
rect 86246 40773 86302 40829
rect 85874 40649 85930 40705
rect 85998 40649 86054 40705
rect 86122 40649 86178 40705
rect 86246 40649 86302 40705
rect 1868 40331 1924 40387
rect 1868 40207 1924 40263
rect 1868 40083 1924 40139
rect 1868 39959 1924 40015
rect 1868 39835 1924 39891
rect 1868 39711 1924 39767
rect 1868 39587 1924 39643
rect 1868 39463 1924 39519
rect 1868 39339 1924 39395
rect 1868 39215 1924 39271
rect 1868 39091 1924 39147
rect 1868 38967 1924 39023
rect 1868 38843 1924 38899
rect 1868 38719 1924 38775
rect 1868 38595 1924 38651
rect 1868 38471 1924 38527
rect 1868 38347 1924 38403
rect 1868 38223 1924 38279
rect 1868 38099 1924 38155
rect 1868 37975 1924 38031
rect 1868 37851 1924 37907
rect 1868 37727 1924 37783
rect 1868 37603 1924 37659
rect 1868 37479 1924 37535
rect 1868 37355 1924 37411
rect 1868 37231 1924 37287
rect 1868 37107 1924 37163
rect 1992 40331 2048 40387
rect 2116 40331 2172 40387
rect 2240 40331 2296 40387
rect 2364 40331 2420 40387
rect 1992 40207 2048 40263
rect 2116 40207 2172 40263
rect 2240 40207 2296 40263
rect 2364 40207 2420 40263
rect 1992 40083 2048 40139
rect 2116 40083 2172 40139
rect 2240 40083 2296 40139
rect 2364 40083 2420 40139
rect 1992 39959 2048 40015
rect 2116 39959 2172 40015
rect 2240 39959 2296 40015
rect 2364 39959 2420 40015
rect 1992 39835 2048 39891
rect 2116 39835 2172 39891
rect 2240 39835 2296 39891
rect 2364 39835 2420 39891
rect 1992 39711 2048 39767
rect 2116 39711 2172 39767
rect 2240 39711 2296 39767
rect 2364 39711 2420 39767
rect 1992 39587 2048 39643
rect 2116 39587 2172 39643
rect 2240 39587 2296 39643
rect 2364 39587 2420 39643
rect 1992 39463 2048 39519
rect 2116 39463 2172 39519
rect 2240 39463 2296 39519
rect 2364 39463 2420 39519
rect 1992 39339 2048 39395
rect 2116 39339 2172 39395
rect 2240 39339 2296 39395
rect 2364 39339 2420 39395
rect 1992 39215 2048 39271
rect 2116 39215 2172 39271
rect 2240 39215 2296 39271
rect 2364 39215 2420 39271
rect 1992 39091 2048 39147
rect 2116 39091 2172 39147
rect 2240 39091 2296 39147
rect 2364 39091 2420 39147
rect 1992 38967 2048 39023
rect 2116 38967 2172 39023
rect 2240 38967 2296 39023
rect 2364 38967 2420 39023
rect 1992 38843 2048 38899
rect 2116 38843 2172 38899
rect 2240 38843 2296 38899
rect 2364 38843 2420 38899
rect 1992 38719 2048 38775
rect 2116 38719 2172 38775
rect 2240 38719 2296 38775
rect 2364 38719 2420 38775
rect 1992 38595 2048 38651
rect 2116 38595 2172 38651
rect 2240 38595 2296 38651
rect 2364 38595 2420 38651
rect 1992 38471 2048 38527
rect 2116 38471 2172 38527
rect 2240 38471 2296 38527
rect 2364 38471 2420 38527
rect 1992 38347 2048 38403
rect 2116 38347 2172 38403
rect 2240 38347 2296 38403
rect 2364 38347 2420 38403
rect 1992 38223 2048 38279
rect 2116 38223 2172 38279
rect 2240 38223 2296 38279
rect 2364 38223 2420 38279
rect 1992 38099 2048 38155
rect 2116 38099 2172 38155
rect 2240 38099 2296 38155
rect 2364 38099 2420 38155
rect 1992 37975 2048 38031
rect 2116 37975 2172 38031
rect 2240 37975 2296 38031
rect 2364 37975 2420 38031
rect 1992 37851 2048 37907
rect 2116 37851 2172 37907
rect 2240 37851 2296 37907
rect 2364 37851 2420 37907
rect 1992 37727 2048 37783
rect 2116 37727 2172 37783
rect 2240 37727 2296 37783
rect 2364 37727 2420 37783
rect 1992 37603 2048 37659
rect 2116 37603 2172 37659
rect 2240 37603 2296 37659
rect 2364 37603 2420 37659
rect 1992 37479 2048 37535
rect 2116 37479 2172 37535
rect 2240 37479 2296 37535
rect 2364 37479 2420 37535
rect 1992 37355 2048 37411
rect 2116 37355 2172 37411
rect 2240 37355 2296 37411
rect 2364 37355 2420 37411
rect 1992 37231 2048 37287
rect 2116 37231 2172 37287
rect 2240 37231 2296 37287
rect 2364 37231 2420 37287
rect 1992 37107 2048 37163
rect 2116 37107 2172 37163
rect 2240 37107 2296 37163
rect 2364 37107 2420 37163
rect 86550 40331 86606 40387
rect 86550 40207 86606 40263
rect 86550 40083 86606 40139
rect 86550 39959 86606 40015
rect 86550 39835 86606 39891
rect 86550 39711 86606 39767
rect 86550 39587 86606 39643
rect 86550 39463 86606 39519
rect 86550 39339 86606 39395
rect 86550 39215 86606 39271
rect 86550 39091 86606 39147
rect 86550 38967 86606 39023
rect 86550 38843 86606 38899
rect 86550 38719 86606 38775
rect 86550 38595 86606 38651
rect 86550 38471 86606 38527
rect 86550 38347 86606 38403
rect 86550 38223 86606 38279
rect 86550 38099 86606 38155
rect 86550 37975 86606 38031
rect 86550 37851 86606 37907
rect 86550 37727 86606 37783
rect 86550 37603 86606 37659
rect 86550 37479 86606 37535
rect 86550 37355 86606 37411
rect 86550 37231 86606 37287
rect 86550 37107 86606 37163
rect 86674 40331 86730 40387
rect 86798 40331 86854 40387
rect 86922 40331 86978 40387
rect 87046 40331 87102 40387
rect 86674 40207 86730 40263
rect 86798 40207 86854 40263
rect 86922 40207 86978 40263
rect 87046 40207 87102 40263
rect 86674 40083 86730 40139
rect 86798 40083 86854 40139
rect 86922 40083 86978 40139
rect 87046 40083 87102 40139
rect 86674 39959 86730 40015
rect 86798 39959 86854 40015
rect 86922 39959 86978 40015
rect 87046 39959 87102 40015
rect 86674 39835 86730 39891
rect 86798 39835 86854 39891
rect 86922 39835 86978 39891
rect 87046 39835 87102 39891
rect 86674 39711 86730 39767
rect 86798 39711 86854 39767
rect 86922 39711 86978 39767
rect 87046 39711 87102 39767
rect 86674 39587 86730 39643
rect 86798 39587 86854 39643
rect 86922 39587 86978 39643
rect 87046 39587 87102 39643
rect 86674 39463 86730 39519
rect 86798 39463 86854 39519
rect 86922 39463 86978 39519
rect 87046 39463 87102 39519
rect 86674 39339 86730 39395
rect 86798 39339 86854 39395
rect 86922 39339 86978 39395
rect 87046 39339 87102 39395
rect 86674 39215 86730 39271
rect 86798 39215 86854 39271
rect 86922 39215 86978 39271
rect 87046 39215 87102 39271
rect 86674 39091 86730 39147
rect 86798 39091 86854 39147
rect 86922 39091 86978 39147
rect 87046 39091 87102 39147
rect 86674 38967 86730 39023
rect 86798 38967 86854 39023
rect 86922 38967 86978 39023
rect 87046 38967 87102 39023
rect 86674 38843 86730 38899
rect 86798 38843 86854 38899
rect 86922 38843 86978 38899
rect 87046 38843 87102 38899
rect 86674 38719 86730 38775
rect 86798 38719 86854 38775
rect 86922 38719 86978 38775
rect 87046 38719 87102 38775
rect 86674 38595 86730 38651
rect 86798 38595 86854 38651
rect 86922 38595 86978 38651
rect 87046 38595 87102 38651
rect 86674 38471 86730 38527
rect 86798 38471 86854 38527
rect 86922 38471 86978 38527
rect 87046 38471 87102 38527
rect 86674 38347 86730 38403
rect 86798 38347 86854 38403
rect 86922 38347 86978 38403
rect 87046 38347 87102 38403
rect 86674 38223 86730 38279
rect 86798 38223 86854 38279
rect 86922 38223 86978 38279
rect 87046 38223 87102 38279
rect 86674 38099 86730 38155
rect 86798 38099 86854 38155
rect 86922 38099 86978 38155
rect 87046 38099 87102 38155
rect 86674 37975 86730 38031
rect 86798 37975 86854 38031
rect 86922 37975 86978 38031
rect 87046 37975 87102 38031
rect 86674 37851 86730 37907
rect 86798 37851 86854 37907
rect 86922 37851 86978 37907
rect 87046 37851 87102 37907
rect 86674 37727 86730 37783
rect 86798 37727 86854 37783
rect 86922 37727 86978 37783
rect 87046 37727 87102 37783
rect 86674 37603 86730 37659
rect 86798 37603 86854 37659
rect 86922 37603 86978 37659
rect 87046 37603 87102 37659
rect 86674 37479 86730 37535
rect 86798 37479 86854 37535
rect 86922 37479 86978 37535
rect 87046 37479 87102 37535
rect 86674 37355 86730 37411
rect 86798 37355 86854 37411
rect 86922 37355 86978 37411
rect 87046 37355 87102 37411
rect 86674 37231 86730 37287
rect 86798 37231 86854 37287
rect 86922 37231 86978 37287
rect 87046 37231 87102 37287
rect 86674 37107 86730 37163
rect 86798 37107 86854 37163
rect 86922 37107 86978 37163
rect 87046 37107 87102 37163
rect 86550 33400 86606 33456
rect 86550 33276 86606 33332
rect 86550 33152 86606 33208
rect 86550 33028 86606 33084
rect 86550 32904 86606 32960
rect 86550 32780 86606 32836
rect 86550 32656 86606 32712
rect 86550 32532 86606 32588
rect 86674 33400 86730 33456
rect 86798 33400 86854 33456
rect 86922 33400 86978 33456
rect 87046 33400 87102 33456
rect 86674 33276 86730 33332
rect 86798 33276 86854 33332
rect 86922 33276 86978 33332
rect 87046 33276 87102 33332
rect 86674 33152 86730 33208
rect 86798 33152 86854 33208
rect 86922 33152 86978 33208
rect 87046 33152 87102 33208
rect 86674 33028 86730 33084
rect 86798 33028 86854 33084
rect 86922 33028 86978 33084
rect 87046 33028 87102 33084
rect 86674 32904 86730 32960
rect 86798 32904 86854 32960
rect 86922 32904 86978 32960
rect 87046 32904 87102 32960
rect 86674 32780 86730 32836
rect 86798 32780 86854 32836
rect 86922 32780 86978 32836
rect 87046 32780 87102 32836
rect 86674 32656 86730 32712
rect 86798 32656 86854 32712
rect 86922 32656 86978 32712
rect 87046 32656 87102 32712
rect 86674 32532 86730 32588
rect 86798 32532 86854 32588
rect 86922 32532 86978 32588
rect 87046 32532 87102 32588
rect 1068 31744 1124 31800
rect 1068 31620 1124 31676
rect 1068 31496 1124 31552
rect 1068 31372 1124 31428
rect 1068 31248 1124 31304
rect 1068 31124 1124 31180
rect 1068 31000 1124 31056
rect 1068 30876 1124 30932
rect 1192 31744 1248 31800
rect 1316 31744 1372 31800
rect 1440 31744 1496 31800
rect 1564 31744 1620 31800
rect 1192 31620 1248 31676
rect 1316 31620 1372 31676
rect 1440 31620 1496 31676
rect 1564 31620 1620 31676
rect 1192 31496 1248 31552
rect 1316 31496 1372 31552
rect 1440 31496 1496 31552
rect 1564 31496 1620 31552
rect 1192 31372 1248 31428
rect 1316 31372 1372 31428
rect 1440 31372 1496 31428
rect 1564 31372 1620 31428
rect 1192 31248 1248 31304
rect 1316 31248 1372 31304
rect 1440 31248 1496 31304
rect 1564 31248 1620 31304
rect 1192 31124 1248 31180
rect 1316 31124 1372 31180
rect 1440 31124 1496 31180
rect 1564 31124 1620 31180
rect 1192 31000 1248 31056
rect 1316 31000 1372 31056
rect 1440 31000 1496 31056
rect 1564 31000 1620 31056
rect 1192 30876 1248 30932
rect 1316 30876 1372 30932
rect 1440 30876 1496 30932
rect 1564 30876 1620 30932
rect 85750 31744 85806 31800
rect 85750 31620 85806 31676
rect 85750 31496 85806 31552
rect 85750 31372 85806 31428
rect 85750 31248 85806 31304
rect 85750 31124 85806 31180
rect 85750 31000 85806 31056
rect 85750 30876 85806 30932
rect 85874 31744 85930 31800
rect 85998 31744 86054 31800
rect 86122 31744 86178 31800
rect 86246 31744 86302 31800
rect 85874 31620 85930 31676
rect 85998 31620 86054 31676
rect 86122 31620 86178 31676
rect 86246 31620 86302 31676
rect 85874 31496 85930 31552
rect 85998 31496 86054 31552
rect 86122 31496 86178 31552
rect 86246 31496 86302 31552
rect 85874 31372 85930 31428
rect 85998 31372 86054 31428
rect 86122 31372 86178 31428
rect 86246 31372 86302 31428
rect 85874 31248 85930 31304
rect 85998 31248 86054 31304
rect 86122 31248 86178 31304
rect 86246 31248 86302 31304
rect 85874 31124 85930 31180
rect 85998 31124 86054 31180
rect 86122 31124 86178 31180
rect 86246 31124 86302 31180
rect 85874 31000 85930 31056
rect 85998 31000 86054 31056
rect 86122 31000 86178 31056
rect 86246 31000 86302 31056
rect 85874 30876 85930 30932
rect 85998 30876 86054 30932
rect 86122 30876 86178 30932
rect 86246 30876 86302 30932
rect 1930 20003 1986 20059
rect 2054 20003 2110 20059
rect 2178 20003 2234 20059
rect 2302 20003 2358 20059
rect 1930 19879 1986 19935
rect 2054 19879 2110 19935
rect 2178 19879 2234 19935
rect 2302 19879 2358 19935
rect 1930 19755 1986 19811
rect 2054 19755 2110 19811
rect 2178 19755 2234 19811
rect 2302 19755 2358 19811
rect 1930 19631 1986 19687
rect 2054 19631 2110 19687
rect 2178 19631 2234 19687
rect 2302 19631 2358 19687
rect 86612 20003 86668 20059
rect 86736 20003 86792 20059
rect 86860 20003 86916 20059
rect 86984 20003 87040 20059
rect 86612 19879 86668 19935
rect 86736 19879 86792 19935
rect 86860 19879 86916 19935
rect 86984 19879 87040 19935
rect 86612 19755 86668 19811
rect 86736 19755 86792 19811
rect 86860 19755 86916 19811
rect 86984 19755 87040 19811
rect 86612 19631 86668 19687
rect 86736 19631 86792 19687
rect 86860 19631 86916 19687
rect 86984 19631 87040 19687
rect 1130 18808 1186 18864
rect 1254 18808 1310 18864
rect 1378 18808 1434 18864
rect 1502 18808 1558 18864
rect 1130 18684 1186 18740
rect 1254 18684 1310 18740
rect 1378 18684 1434 18740
rect 1502 18684 1558 18740
rect 1130 18560 1186 18616
rect 1254 18560 1310 18616
rect 1378 18560 1434 18616
rect 1502 18560 1558 18616
rect 1130 18436 1186 18492
rect 1254 18436 1310 18492
rect 1378 18436 1434 18492
rect 1502 18436 1558 18492
rect 85812 18808 85868 18864
rect 85936 18808 85992 18864
rect 86060 18808 86116 18864
rect 86184 18808 86240 18864
rect 85812 18684 85868 18740
rect 85936 18684 85992 18740
rect 86060 18684 86116 18740
rect 86184 18684 86240 18740
rect 85812 18560 85868 18616
rect 85936 18560 85992 18616
rect 86060 18560 86116 18616
rect 86184 18560 86240 18616
rect 85812 18436 85868 18492
rect 85936 18436 85992 18492
rect 86060 18436 86116 18492
rect 86184 18436 86240 18492
rect 86612 17908 86668 17964
rect 86736 17908 86792 17964
rect 86860 17908 86916 17964
rect 86984 17908 87040 17964
rect 1930 17784 1986 17840
rect 2054 17784 2110 17840
rect 2178 17784 2234 17840
rect 2302 17784 2358 17840
rect 1930 17660 1986 17716
rect 2054 17660 2110 17716
rect 2178 17660 2234 17716
rect 2302 17660 2358 17716
rect 86612 17784 86668 17840
rect 86736 17784 86792 17840
rect 86860 17784 86916 17840
rect 86984 17784 87040 17840
rect 86612 17660 86668 17716
rect 86736 17660 86792 17716
rect 86860 17660 86916 17716
rect 86984 17660 87040 17716
rect 86612 17536 86668 17592
rect 86736 17536 86792 17592
rect 86860 17536 86916 17592
rect 86984 17536 87040 17592
rect 1130 17008 1186 17064
rect 1254 17008 1310 17064
rect 1378 17008 1434 17064
rect 1502 17008 1558 17064
rect 1130 16884 1186 16940
rect 1254 16884 1310 16940
rect 1378 16884 1434 16940
rect 1502 16884 1558 16940
rect 1130 16760 1186 16816
rect 1254 16760 1310 16816
rect 1378 16760 1434 16816
rect 1502 16760 1558 16816
rect 1130 16636 1186 16692
rect 1254 16636 1310 16692
rect 1378 16636 1434 16692
rect 1502 16636 1558 16692
rect 85812 17008 85868 17064
rect 85936 17008 85992 17064
rect 86060 17008 86116 17064
rect 86184 17008 86240 17064
rect 85812 16884 85868 16940
rect 85936 16884 85992 16940
rect 86060 16884 86116 16940
rect 86184 16884 86240 16940
rect 85812 16760 85868 16816
rect 85936 16760 85992 16816
rect 86060 16760 86116 16816
rect 86184 16760 86240 16816
rect 85812 16636 85868 16692
rect 85936 16636 85992 16692
rect 86060 16636 86116 16692
rect 86184 16636 86240 16692
rect 86612 16108 86668 16164
rect 86736 16108 86792 16164
rect 86860 16108 86916 16164
rect 86984 16108 87040 16164
rect 1930 15984 1986 16040
rect 2054 15984 2110 16040
rect 2178 15984 2234 16040
rect 2302 15984 2358 16040
rect 1930 15860 1986 15916
rect 2054 15860 2110 15916
rect 2178 15860 2234 15916
rect 2302 15860 2358 15916
rect 86612 15984 86668 16040
rect 86736 15984 86792 16040
rect 86860 15984 86916 16040
rect 86984 15984 87040 16040
rect 86612 15860 86668 15916
rect 86736 15860 86792 15916
rect 86860 15860 86916 15916
rect 86984 15860 87040 15916
rect 86612 15736 86668 15792
rect 86736 15736 86792 15792
rect 86860 15736 86916 15792
rect 86984 15736 87040 15792
rect 1130 15208 1186 15264
rect 1254 15208 1310 15264
rect 1378 15208 1434 15264
rect 1502 15208 1558 15264
rect 1130 15084 1186 15140
rect 1254 15084 1310 15140
rect 1378 15084 1434 15140
rect 1502 15084 1558 15140
rect 1130 14960 1186 15016
rect 1254 14960 1310 15016
rect 1378 14960 1434 15016
rect 1502 14960 1558 15016
rect 1130 14836 1186 14892
rect 1254 14836 1310 14892
rect 1378 14836 1434 14892
rect 1502 14836 1558 14892
rect 85812 15208 85868 15264
rect 85936 15208 85992 15264
rect 86060 15208 86116 15264
rect 86184 15208 86240 15264
rect 85812 15084 85868 15140
rect 85936 15084 85992 15140
rect 86060 15084 86116 15140
rect 86184 15084 86240 15140
rect 85812 14960 85868 15016
rect 85936 14960 85992 15016
rect 86060 14960 86116 15016
rect 86184 14960 86240 15016
rect 85812 14836 85868 14892
rect 85936 14836 85992 14892
rect 86060 14836 86116 14892
rect 86184 14836 86240 14892
rect 86612 14308 86668 14364
rect 86736 14308 86792 14364
rect 86860 14308 86916 14364
rect 86984 14308 87040 14364
rect 1930 14184 1986 14240
rect 2054 14184 2110 14240
rect 2178 14184 2234 14240
rect 2302 14184 2358 14240
rect 1930 14060 1986 14116
rect 2054 14060 2110 14116
rect 2178 14060 2234 14116
rect 2302 14060 2358 14116
rect 86612 14184 86668 14240
rect 86736 14184 86792 14240
rect 86860 14184 86916 14240
rect 86984 14184 87040 14240
rect 86612 14060 86668 14116
rect 86736 14060 86792 14116
rect 86860 14060 86916 14116
rect 86984 14060 87040 14116
rect 86612 13936 86668 13992
rect 86736 13936 86792 13992
rect 86860 13936 86916 13992
rect 86984 13936 87040 13992
rect 1130 13408 1186 13464
rect 1254 13408 1310 13464
rect 1378 13408 1434 13464
rect 1502 13408 1558 13464
rect 1130 13284 1186 13340
rect 1254 13284 1310 13340
rect 1378 13284 1434 13340
rect 1502 13284 1558 13340
rect 1130 13160 1186 13216
rect 1254 13160 1310 13216
rect 1378 13160 1434 13216
rect 1502 13160 1558 13216
rect 1130 13036 1186 13092
rect 1254 13036 1310 13092
rect 1378 13036 1434 13092
rect 1502 13036 1558 13092
rect 85812 13408 85868 13464
rect 85936 13408 85992 13464
rect 86060 13408 86116 13464
rect 86184 13408 86240 13464
rect 85812 13284 85868 13340
rect 85936 13284 85992 13340
rect 86060 13284 86116 13340
rect 86184 13284 86240 13340
rect 85812 13160 85868 13216
rect 85936 13160 85992 13216
rect 86060 13160 86116 13216
rect 86184 13160 86240 13216
rect 85812 13036 85868 13092
rect 85936 13036 85992 13092
rect 86060 13036 86116 13092
rect 86184 13036 86240 13092
rect 86612 12508 86668 12564
rect 86736 12508 86792 12564
rect 86860 12508 86916 12564
rect 86984 12508 87040 12564
rect 1930 12384 1986 12440
rect 2054 12384 2110 12440
rect 2178 12384 2234 12440
rect 2302 12384 2358 12440
rect 1930 12260 1986 12316
rect 2054 12260 2110 12316
rect 2178 12260 2234 12316
rect 2302 12260 2358 12316
rect 86612 12384 86668 12440
rect 86736 12384 86792 12440
rect 86860 12384 86916 12440
rect 86984 12384 87040 12440
rect 86612 12260 86668 12316
rect 86736 12260 86792 12316
rect 86860 12260 86916 12316
rect 86984 12260 87040 12316
rect 86612 12136 86668 12192
rect 86736 12136 86792 12192
rect 86860 12136 86916 12192
rect 86984 12136 87040 12192
rect 1130 11608 1186 11664
rect 1254 11608 1310 11664
rect 1378 11608 1434 11664
rect 1502 11608 1558 11664
rect 1130 11484 1186 11540
rect 1254 11484 1310 11540
rect 1378 11484 1434 11540
rect 1502 11484 1558 11540
rect 1130 11360 1186 11416
rect 1254 11360 1310 11416
rect 1378 11360 1434 11416
rect 1502 11360 1558 11416
rect 1130 11236 1186 11292
rect 1254 11236 1310 11292
rect 1378 11236 1434 11292
rect 1502 11236 1558 11292
rect 85812 11608 85868 11664
rect 85936 11608 85992 11664
rect 86060 11608 86116 11664
rect 86184 11608 86240 11664
rect 85812 11484 85868 11540
rect 85936 11484 85992 11540
rect 86060 11484 86116 11540
rect 86184 11484 86240 11540
rect 85812 11360 85868 11416
rect 85936 11360 85992 11416
rect 86060 11360 86116 11416
rect 86184 11360 86240 11416
rect 85812 11236 85868 11292
rect 85936 11236 85992 11292
rect 86060 11236 86116 11292
rect 86184 11236 86240 11292
rect 86612 10708 86668 10764
rect 86736 10708 86792 10764
rect 86860 10708 86916 10764
rect 86984 10708 87040 10764
rect 1930 10584 1986 10640
rect 2054 10584 2110 10640
rect 2178 10584 2234 10640
rect 2302 10584 2358 10640
rect 1930 10460 1986 10516
rect 2054 10460 2110 10516
rect 2178 10460 2234 10516
rect 2302 10460 2358 10516
rect 86612 10584 86668 10640
rect 86736 10584 86792 10640
rect 86860 10584 86916 10640
rect 86984 10584 87040 10640
rect 86612 10460 86668 10516
rect 86736 10460 86792 10516
rect 86860 10460 86916 10516
rect 86984 10460 87040 10516
rect 86612 10336 86668 10392
rect 86736 10336 86792 10392
rect 86860 10336 86916 10392
rect 86984 10336 87040 10392
rect 1130 9808 1186 9864
rect 1254 9808 1310 9864
rect 1378 9808 1434 9864
rect 1502 9808 1558 9864
rect 1130 9684 1186 9740
rect 1254 9684 1310 9740
rect 1378 9684 1434 9740
rect 1502 9684 1558 9740
rect 1130 9560 1186 9616
rect 1254 9560 1310 9616
rect 1378 9560 1434 9616
rect 1502 9560 1558 9616
rect 1130 9436 1186 9492
rect 1254 9436 1310 9492
rect 1378 9436 1434 9492
rect 1502 9436 1558 9492
rect 85812 9808 85868 9864
rect 85936 9808 85992 9864
rect 86060 9808 86116 9864
rect 86184 9808 86240 9864
rect 85812 9684 85868 9740
rect 85936 9684 85992 9740
rect 86060 9684 86116 9740
rect 86184 9684 86240 9740
rect 85812 9560 85868 9616
rect 85936 9560 85992 9616
rect 86060 9560 86116 9616
rect 86184 9560 86240 9616
rect 85812 9436 85868 9492
rect 85936 9436 85992 9492
rect 86060 9436 86116 9492
rect 86184 9436 86240 9492
rect 86612 8908 86668 8964
rect 86736 8908 86792 8964
rect 86860 8908 86916 8964
rect 86984 8908 87040 8964
rect 1930 8784 1986 8840
rect 2054 8784 2110 8840
rect 2178 8784 2234 8840
rect 2302 8784 2358 8840
rect 1930 8660 1986 8716
rect 2054 8660 2110 8716
rect 2178 8660 2234 8716
rect 2302 8660 2358 8716
rect 86612 8784 86668 8840
rect 86736 8784 86792 8840
rect 86860 8784 86916 8840
rect 86984 8784 87040 8840
rect 86612 8660 86668 8716
rect 86736 8660 86792 8716
rect 86860 8660 86916 8716
rect 86984 8660 87040 8716
rect 86612 8536 86668 8592
rect 86736 8536 86792 8592
rect 86860 8536 86916 8592
rect 86984 8536 87040 8592
rect 1130 8008 1186 8064
rect 1254 8008 1310 8064
rect 1378 8008 1434 8064
rect 1502 8008 1558 8064
rect 1130 7884 1186 7940
rect 1254 7884 1310 7940
rect 1378 7884 1434 7940
rect 1502 7884 1558 7940
rect 1130 7760 1186 7816
rect 1254 7760 1310 7816
rect 1378 7760 1434 7816
rect 1502 7760 1558 7816
rect 1130 7636 1186 7692
rect 1254 7636 1310 7692
rect 1378 7636 1434 7692
rect 1502 7636 1558 7692
rect 85812 8008 85868 8064
rect 85936 8008 85992 8064
rect 86060 8008 86116 8064
rect 86184 8008 86240 8064
rect 85812 7884 85868 7940
rect 85936 7884 85992 7940
rect 86060 7884 86116 7940
rect 86184 7884 86240 7940
rect 85812 7760 85868 7816
rect 85936 7760 85992 7816
rect 86060 7760 86116 7816
rect 86184 7760 86240 7816
rect 85812 7636 85868 7692
rect 85936 7636 85992 7692
rect 86060 7636 86116 7692
rect 86184 7636 86240 7692
rect 86612 7108 86668 7164
rect 86736 7108 86792 7164
rect 86860 7108 86916 7164
rect 86984 7108 87040 7164
rect 1930 6984 1986 7040
rect 2054 6984 2110 7040
rect 2178 6984 2234 7040
rect 2302 6984 2358 7040
rect 1930 6860 1986 6916
rect 2054 6860 2110 6916
rect 2178 6860 2234 6916
rect 2302 6860 2358 6916
rect 86612 6984 86668 7040
rect 86736 6984 86792 7040
rect 86860 6984 86916 7040
rect 86984 6984 87040 7040
rect 86612 6860 86668 6916
rect 86736 6860 86792 6916
rect 86860 6860 86916 6916
rect 86984 6860 87040 6916
rect 86612 6736 86668 6792
rect 86736 6736 86792 6792
rect 86860 6736 86916 6792
rect 86984 6736 87040 6792
rect 1130 6208 1186 6264
rect 1254 6208 1310 6264
rect 1378 6208 1434 6264
rect 1502 6208 1558 6264
rect 1130 6084 1186 6140
rect 1254 6084 1310 6140
rect 1378 6084 1434 6140
rect 1502 6084 1558 6140
rect 1130 5960 1186 6016
rect 1254 5960 1310 6016
rect 1378 5960 1434 6016
rect 1502 5960 1558 6016
rect 1130 5836 1186 5892
rect 1254 5836 1310 5892
rect 1378 5836 1434 5892
rect 1502 5836 1558 5892
rect 85812 6208 85868 6264
rect 85936 6208 85992 6264
rect 86060 6208 86116 6264
rect 86184 6208 86240 6264
rect 85812 6084 85868 6140
rect 85936 6084 85992 6140
rect 86060 6084 86116 6140
rect 86184 6084 86240 6140
rect 85812 5960 85868 6016
rect 85936 5960 85992 6016
rect 86060 5960 86116 6016
rect 86184 5960 86240 6016
rect 85812 5836 85868 5892
rect 85936 5836 85992 5892
rect 86060 5836 86116 5892
rect 86184 5836 86240 5892
rect 86612 5308 86668 5364
rect 86736 5308 86792 5364
rect 86860 5308 86916 5364
rect 86984 5308 87040 5364
rect 1930 5184 1986 5240
rect 2054 5184 2110 5240
rect 2178 5184 2234 5240
rect 2302 5184 2358 5240
rect 1930 5060 1986 5116
rect 2054 5060 2110 5116
rect 2178 5060 2234 5116
rect 2302 5060 2358 5116
rect 86612 5184 86668 5240
rect 86736 5184 86792 5240
rect 86860 5184 86916 5240
rect 86984 5184 87040 5240
rect 86612 5060 86668 5116
rect 86736 5060 86792 5116
rect 86860 5060 86916 5116
rect 86984 5060 87040 5116
rect 86612 4936 86668 4992
rect 86736 4936 86792 4992
rect 86860 4936 86916 4992
rect 86984 4936 87040 4992
rect 1130 4408 1186 4464
rect 1254 4408 1310 4464
rect 1378 4408 1434 4464
rect 1502 4408 1558 4464
rect 1130 4284 1186 4340
rect 1254 4284 1310 4340
rect 1378 4284 1434 4340
rect 1502 4284 1558 4340
rect 1130 4160 1186 4216
rect 1254 4160 1310 4216
rect 1378 4160 1434 4216
rect 1502 4160 1558 4216
rect 1130 4036 1186 4092
rect 1254 4036 1310 4092
rect 1378 4036 1434 4092
rect 1502 4036 1558 4092
rect 85812 4408 85868 4464
rect 85936 4408 85992 4464
rect 86060 4408 86116 4464
rect 86184 4408 86240 4464
rect 85812 4284 85868 4340
rect 85936 4284 85992 4340
rect 86060 4284 86116 4340
rect 86184 4284 86240 4340
rect 85812 4160 85868 4216
rect 85936 4160 85992 4216
rect 86060 4160 86116 4216
rect 86184 4160 86240 4216
rect 85812 4036 85868 4092
rect 85936 4036 85992 4092
rect 86060 4036 86116 4092
rect 86184 4036 86240 4092
rect 86612 3576 86668 3632
rect 86736 3576 86792 3632
rect 86860 3576 86916 3632
rect 86984 3576 87040 3632
rect 1930 3384 1986 3440
rect 2054 3384 2110 3440
rect 2178 3384 2234 3440
rect 2302 3384 2358 3440
rect 1930 3260 1986 3316
rect 2054 3260 2110 3316
rect 2178 3260 2234 3316
rect 2302 3260 2358 3316
rect 86612 3452 86668 3508
rect 86736 3452 86792 3508
rect 86860 3452 86916 3508
rect 86984 3452 87040 3508
rect 86612 3328 86668 3384
rect 86736 3328 86792 3384
rect 86860 3328 86916 3384
rect 86984 3328 87040 3384
rect 86612 3204 86668 3260
rect 86736 3204 86792 3260
rect 86860 3204 86916 3260
rect 86984 3204 87040 3260
<< metal4 >>
rect 1044 42689 1644 52528
rect 1044 42633 1068 42689
rect 1124 42633 1192 42689
rect 1248 42633 1316 42689
rect 1372 42633 1440 42689
rect 1496 42633 1564 42689
rect 1620 42633 1644 42689
rect 1044 42565 1644 42633
rect 1044 42509 1068 42565
rect 1124 42509 1192 42565
rect 1248 42509 1316 42565
rect 1372 42509 1440 42565
rect 1496 42509 1564 42565
rect 1620 42509 1644 42565
rect 1044 42441 1644 42509
rect 1044 42385 1068 42441
rect 1124 42385 1192 42441
rect 1248 42385 1316 42441
rect 1372 42385 1440 42441
rect 1496 42385 1564 42441
rect 1620 42385 1644 42441
rect 1044 42317 1644 42385
rect 1044 42261 1068 42317
rect 1124 42261 1192 42317
rect 1248 42261 1316 42317
rect 1372 42261 1440 42317
rect 1496 42261 1564 42317
rect 1620 42261 1644 42317
rect 1044 42193 1644 42261
rect 1044 42137 1068 42193
rect 1124 42137 1192 42193
rect 1248 42137 1316 42193
rect 1372 42137 1440 42193
rect 1496 42137 1564 42193
rect 1620 42137 1644 42193
rect 1044 42069 1644 42137
rect 1044 42013 1068 42069
rect 1124 42013 1192 42069
rect 1248 42013 1316 42069
rect 1372 42013 1440 42069
rect 1496 42013 1564 42069
rect 1620 42013 1644 42069
rect 1044 41945 1644 42013
rect 1044 41889 1068 41945
rect 1124 41889 1192 41945
rect 1248 41889 1316 41945
rect 1372 41889 1440 41945
rect 1496 41889 1564 41945
rect 1620 41889 1644 41945
rect 1044 41821 1644 41889
rect 1044 41765 1068 41821
rect 1124 41765 1192 41821
rect 1248 41765 1316 41821
rect 1372 41765 1440 41821
rect 1496 41765 1564 41821
rect 1620 41765 1644 41821
rect 1044 41697 1644 41765
rect 1044 41641 1068 41697
rect 1124 41641 1192 41697
rect 1248 41641 1316 41697
rect 1372 41641 1440 41697
rect 1496 41641 1564 41697
rect 1620 41641 1644 41697
rect 1044 41573 1644 41641
rect 1044 41517 1068 41573
rect 1124 41517 1192 41573
rect 1248 41517 1316 41573
rect 1372 41517 1440 41573
rect 1496 41517 1564 41573
rect 1620 41517 1644 41573
rect 1044 41449 1644 41517
rect 1044 41393 1068 41449
rect 1124 41393 1192 41449
rect 1248 41393 1316 41449
rect 1372 41393 1440 41449
rect 1496 41393 1564 41449
rect 1620 41393 1644 41449
rect 1044 41325 1644 41393
rect 1044 41269 1068 41325
rect 1124 41269 1192 41325
rect 1248 41269 1316 41325
rect 1372 41269 1440 41325
rect 1496 41269 1564 41325
rect 1620 41269 1644 41325
rect 1044 41201 1644 41269
rect 1044 41145 1068 41201
rect 1124 41145 1192 41201
rect 1248 41145 1316 41201
rect 1372 41145 1440 41201
rect 1496 41145 1564 41201
rect 1620 41145 1644 41201
rect 1044 41077 1644 41145
rect 1044 41021 1068 41077
rect 1124 41021 1192 41077
rect 1248 41021 1316 41077
rect 1372 41021 1440 41077
rect 1496 41021 1564 41077
rect 1620 41021 1644 41077
rect 1044 40953 1644 41021
rect 1044 40897 1068 40953
rect 1124 40897 1192 40953
rect 1248 40897 1316 40953
rect 1372 40897 1440 40953
rect 1496 40897 1564 40953
rect 1620 40897 1644 40953
rect 1044 40829 1644 40897
rect 1044 40773 1068 40829
rect 1124 40773 1192 40829
rect 1248 40773 1316 40829
rect 1372 40773 1440 40829
rect 1496 40773 1564 40829
rect 1620 40773 1644 40829
rect 1044 40705 1644 40773
rect 1044 40649 1068 40705
rect 1124 40649 1192 40705
rect 1248 40649 1316 40705
rect 1372 40649 1440 40705
rect 1496 40649 1564 40705
rect 1620 40649 1644 40705
rect 1044 31800 1644 40649
rect 1044 31744 1068 31800
rect 1124 31744 1192 31800
rect 1248 31744 1316 31800
rect 1372 31744 1440 31800
rect 1496 31744 1564 31800
rect 1620 31744 1644 31800
rect 1044 31676 1644 31744
rect 1044 31620 1068 31676
rect 1124 31620 1192 31676
rect 1248 31620 1316 31676
rect 1372 31620 1440 31676
rect 1496 31620 1564 31676
rect 1620 31620 1644 31676
rect 1044 31552 1644 31620
rect 1044 31496 1068 31552
rect 1124 31496 1192 31552
rect 1248 31496 1316 31552
rect 1372 31496 1440 31552
rect 1496 31496 1564 31552
rect 1620 31496 1644 31552
rect 1044 31428 1644 31496
rect 1044 31372 1068 31428
rect 1124 31372 1192 31428
rect 1248 31372 1316 31428
rect 1372 31372 1440 31428
rect 1496 31372 1564 31428
rect 1620 31372 1644 31428
rect 1044 31304 1644 31372
rect 1044 31248 1068 31304
rect 1124 31248 1192 31304
rect 1248 31248 1316 31304
rect 1372 31248 1440 31304
rect 1496 31248 1564 31304
rect 1620 31248 1644 31304
rect 1044 31180 1644 31248
rect 1044 31124 1068 31180
rect 1124 31124 1192 31180
rect 1248 31124 1316 31180
rect 1372 31124 1440 31180
rect 1496 31124 1564 31180
rect 1620 31124 1644 31180
rect 1044 31056 1644 31124
rect 1044 31000 1068 31056
rect 1124 31000 1192 31056
rect 1248 31000 1316 31056
rect 1372 31000 1440 31056
rect 1496 31000 1564 31056
rect 1620 31000 1644 31056
rect 1044 30932 1644 31000
rect 1044 30876 1068 30932
rect 1124 30876 1192 30932
rect 1248 30876 1316 30932
rect 1372 30876 1440 30932
rect 1496 30876 1564 30932
rect 1620 30876 1644 30932
rect 1044 18864 1644 30876
rect 1044 18808 1130 18864
rect 1186 18808 1254 18864
rect 1310 18808 1378 18864
rect 1434 18808 1502 18864
rect 1558 18808 1644 18864
rect 1044 18740 1644 18808
rect 1044 18684 1130 18740
rect 1186 18684 1254 18740
rect 1310 18684 1378 18740
rect 1434 18684 1502 18740
rect 1558 18684 1644 18740
rect 1044 18616 1644 18684
rect 1044 18560 1130 18616
rect 1186 18560 1254 18616
rect 1310 18560 1378 18616
rect 1434 18560 1502 18616
rect 1558 18560 1644 18616
rect 1044 18492 1644 18560
rect 1044 18436 1130 18492
rect 1186 18436 1254 18492
rect 1310 18436 1378 18492
rect 1434 18436 1502 18492
rect 1558 18436 1644 18492
rect 1044 17064 1644 18436
rect 1044 17008 1130 17064
rect 1186 17008 1254 17064
rect 1310 17008 1378 17064
rect 1434 17008 1502 17064
rect 1558 17008 1644 17064
rect 1044 16940 1644 17008
rect 1044 16884 1130 16940
rect 1186 16884 1254 16940
rect 1310 16884 1378 16940
rect 1434 16884 1502 16940
rect 1558 16884 1644 16940
rect 1044 16816 1644 16884
rect 1044 16760 1130 16816
rect 1186 16760 1254 16816
rect 1310 16760 1378 16816
rect 1434 16760 1502 16816
rect 1558 16760 1644 16816
rect 1044 16692 1644 16760
rect 1044 16636 1130 16692
rect 1186 16636 1254 16692
rect 1310 16636 1378 16692
rect 1434 16636 1502 16692
rect 1558 16636 1644 16692
rect 1044 15264 1644 16636
rect 1044 15208 1130 15264
rect 1186 15208 1254 15264
rect 1310 15208 1378 15264
rect 1434 15208 1502 15264
rect 1558 15208 1644 15264
rect 1044 15140 1644 15208
rect 1044 15084 1130 15140
rect 1186 15084 1254 15140
rect 1310 15084 1378 15140
rect 1434 15084 1502 15140
rect 1558 15084 1644 15140
rect 1044 15016 1644 15084
rect 1044 14960 1130 15016
rect 1186 14960 1254 15016
rect 1310 14960 1378 15016
rect 1434 14960 1502 15016
rect 1558 14960 1644 15016
rect 1044 14892 1644 14960
rect 1044 14836 1130 14892
rect 1186 14836 1254 14892
rect 1310 14836 1378 14892
rect 1434 14836 1502 14892
rect 1558 14836 1644 14892
rect 1044 13464 1644 14836
rect 1044 13408 1130 13464
rect 1186 13408 1254 13464
rect 1310 13408 1378 13464
rect 1434 13408 1502 13464
rect 1558 13408 1644 13464
rect 1044 13340 1644 13408
rect 1044 13284 1130 13340
rect 1186 13284 1254 13340
rect 1310 13284 1378 13340
rect 1434 13284 1502 13340
rect 1558 13284 1644 13340
rect 1044 13216 1644 13284
rect 1044 13160 1130 13216
rect 1186 13160 1254 13216
rect 1310 13160 1378 13216
rect 1434 13160 1502 13216
rect 1558 13160 1644 13216
rect 1044 13092 1644 13160
rect 1044 13036 1130 13092
rect 1186 13036 1254 13092
rect 1310 13036 1378 13092
rect 1434 13036 1502 13092
rect 1558 13036 1644 13092
rect 1044 11664 1644 13036
rect 1044 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1644 11664
rect 1044 11540 1644 11608
rect 1044 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1644 11540
rect 1044 11416 1644 11484
rect 1044 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1644 11416
rect 1044 11292 1644 11360
rect 1044 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1644 11292
rect 1044 9864 1644 11236
rect 1044 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1644 9864
rect 1044 9740 1644 9808
rect 1044 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1644 9740
rect 1044 9616 1644 9684
rect 1044 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1644 9616
rect 1044 9492 1644 9560
rect 1044 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1644 9492
rect 1044 8064 1644 9436
rect 1044 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1644 8064
rect 1044 7940 1644 8008
rect 1044 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1644 7940
rect 1044 7816 1644 7884
rect 1044 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1644 7816
rect 1044 7692 1644 7760
rect 1044 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1644 7692
rect 1044 6264 1644 7636
rect 1044 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1644 6264
rect 1044 6140 1644 6208
rect 1044 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1644 6140
rect 1044 6016 1644 6084
rect 1044 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1644 6016
rect 1044 5892 1644 5960
rect 1044 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1644 5892
rect 1044 4464 1644 5836
rect 1044 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1644 4464
rect 1044 4340 1644 4408
rect 1044 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1644 4340
rect 1044 4216 1644 4284
rect 1044 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1644 4216
rect 1044 4092 1644 4160
rect 1044 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1644 4092
rect 1044 3136 1644 4036
rect 1844 52225 2444 52528
rect 1844 52169 1901 52225
rect 1957 52169 2444 52225
rect 1844 52101 2444 52169
rect 1844 52045 1901 52101
rect 1957 52045 2444 52101
rect 1844 51977 2444 52045
rect 1844 51921 1901 51977
rect 1957 51921 2444 51977
rect 1844 51853 2444 51921
rect 1844 51797 1901 51853
rect 1957 51797 2444 51853
rect 1844 51729 2444 51797
rect 1844 51673 1901 51729
rect 1957 51673 2444 51729
rect 1844 51605 2444 51673
rect 1844 51549 1901 51605
rect 1957 51549 2444 51605
rect 1844 51481 2444 51549
rect 1844 51425 1901 51481
rect 1957 51425 2444 51481
rect 1844 51357 2444 51425
rect 1844 51301 1901 51357
rect 1957 51301 2444 51357
rect 1844 51233 2444 51301
rect 1844 51177 1901 51233
rect 1957 51177 2444 51233
rect 1844 51109 2444 51177
rect 1844 51053 1901 51109
rect 1957 51053 2444 51109
rect 1844 47701 2444 51053
rect 1844 47645 1930 47701
rect 1986 47645 2054 47701
rect 2110 47645 2178 47701
rect 2234 47645 2302 47701
rect 2358 47645 2444 47701
rect 1844 47577 2444 47645
rect 1844 47521 1930 47577
rect 1986 47521 2054 47577
rect 2110 47521 2178 47577
rect 2234 47521 2302 47577
rect 2358 47521 2444 47577
rect 1844 47453 2444 47521
rect 1844 47397 1930 47453
rect 1986 47397 2054 47453
rect 2110 47397 2178 47453
rect 2234 47397 2302 47453
rect 2358 47397 2444 47453
rect 1844 47329 2444 47397
rect 1844 47273 1930 47329
rect 1986 47273 2054 47329
rect 2110 47273 2178 47329
rect 2234 47273 2302 47329
rect 2358 47273 2444 47329
rect 1844 40387 2444 47273
rect 1844 40331 1868 40387
rect 1924 40331 1992 40387
rect 2048 40331 2116 40387
rect 2172 40331 2240 40387
rect 2296 40331 2364 40387
rect 2420 40331 2444 40387
rect 1844 40263 2444 40331
rect 1844 40207 1868 40263
rect 1924 40207 1992 40263
rect 2048 40207 2116 40263
rect 2172 40207 2240 40263
rect 2296 40207 2364 40263
rect 2420 40207 2444 40263
rect 1844 40139 2444 40207
rect 1844 40083 1868 40139
rect 1924 40083 1992 40139
rect 2048 40083 2116 40139
rect 2172 40083 2240 40139
rect 2296 40083 2364 40139
rect 2420 40083 2444 40139
rect 1844 40015 2444 40083
rect 1844 39959 1868 40015
rect 1924 39959 1992 40015
rect 2048 39959 2116 40015
rect 2172 39959 2240 40015
rect 2296 39959 2364 40015
rect 2420 39959 2444 40015
rect 1844 39891 2444 39959
rect 1844 39835 1868 39891
rect 1924 39835 1992 39891
rect 2048 39835 2116 39891
rect 2172 39835 2240 39891
rect 2296 39835 2364 39891
rect 2420 39835 2444 39891
rect 1844 39767 2444 39835
rect 1844 39711 1868 39767
rect 1924 39711 1992 39767
rect 2048 39711 2116 39767
rect 2172 39711 2240 39767
rect 2296 39711 2364 39767
rect 2420 39711 2444 39767
rect 1844 39643 2444 39711
rect 1844 39587 1868 39643
rect 1924 39587 1992 39643
rect 2048 39587 2116 39643
rect 2172 39587 2240 39643
rect 2296 39587 2364 39643
rect 2420 39587 2444 39643
rect 1844 39519 2444 39587
rect 1844 39463 1868 39519
rect 1924 39463 1992 39519
rect 2048 39463 2116 39519
rect 2172 39463 2240 39519
rect 2296 39463 2364 39519
rect 2420 39463 2444 39519
rect 1844 39395 2444 39463
rect 1844 39339 1868 39395
rect 1924 39339 1992 39395
rect 2048 39339 2116 39395
rect 2172 39339 2240 39395
rect 2296 39339 2364 39395
rect 2420 39339 2444 39395
rect 1844 39271 2444 39339
rect 1844 39215 1868 39271
rect 1924 39215 1992 39271
rect 2048 39215 2116 39271
rect 2172 39215 2240 39271
rect 2296 39215 2364 39271
rect 2420 39215 2444 39271
rect 1844 39147 2444 39215
rect 1844 39091 1868 39147
rect 1924 39091 1992 39147
rect 2048 39091 2116 39147
rect 2172 39091 2240 39147
rect 2296 39091 2364 39147
rect 2420 39091 2444 39147
rect 1844 39023 2444 39091
rect 1844 38967 1868 39023
rect 1924 38967 1992 39023
rect 2048 38967 2116 39023
rect 2172 38967 2240 39023
rect 2296 38967 2364 39023
rect 2420 38967 2444 39023
rect 1844 38899 2444 38967
rect 1844 38843 1868 38899
rect 1924 38843 1992 38899
rect 2048 38843 2116 38899
rect 2172 38843 2240 38899
rect 2296 38843 2364 38899
rect 2420 38843 2444 38899
rect 1844 38775 2444 38843
rect 1844 38719 1868 38775
rect 1924 38719 1992 38775
rect 2048 38719 2116 38775
rect 2172 38719 2240 38775
rect 2296 38719 2364 38775
rect 2420 38719 2444 38775
rect 1844 38651 2444 38719
rect 1844 38595 1868 38651
rect 1924 38595 1992 38651
rect 2048 38595 2116 38651
rect 2172 38595 2240 38651
rect 2296 38595 2364 38651
rect 2420 38595 2444 38651
rect 1844 38527 2444 38595
rect 1844 38471 1868 38527
rect 1924 38471 1992 38527
rect 2048 38471 2116 38527
rect 2172 38471 2240 38527
rect 2296 38471 2364 38527
rect 2420 38471 2444 38527
rect 1844 38403 2444 38471
rect 1844 38347 1868 38403
rect 1924 38347 1992 38403
rect 2048 38347 2116 38403
rect 2172 38347 2240 38403
rect 2296 38347 2364 38403
rect 2420 38347 2444 38403
rect 1844 38279 2444 38347
rect 1844 38223 1868 38279
rect 1924 38223 1992 38279
rect 2048 38223 2116 38279
rect 2172 38223 2240 38279
rect 2296 38223 2364 38279
rect 2420 38223 2444 38279
rect 1844 38155 2444 38223
rect 1844 38099 1868 38155
rect 1924 38099 1992 38155
rect 2048 38099 2116 38155
rect 2172 38099 2240 38155
rect 2296 38099 2364 38155
rect 2420 38099 2444 38155
rect 1844 38031 2444 38099
rect 1844 37975 1868 38031
rect 1924 37975 1992 38031
rect 2048 37975 2116 38031
rect 2172 37975 2240 38031
rect 2296 37975 2364 38031
rect 2420 37975 2444 38031
rect 1844 37907 2444 37975
rect 1844 37851 1868 37907
rect 1924 37851 1992 37907
rect 2048 37851 2116 37907
rect 2172 37851 2240 37907
rect 2296 37851 2364 37907
rect 2420 37851 2444 37907
rect 1844 37783 2444 37851
rect 1844 37727 1868 37783
rect 1924 37727 1992 37783
rect 2048 37727 2116 37783
rect 2172 37727 2240 37783
rect 2296 37727 2364 37783
rect 2420 37727 2444 37783
rect 1844 37659 2444 37727
rect 1844 37603 1868 37659
rect 1924 37603 1992 37659
rect 2048 37603 2116 37659
rect 2172 37603 2240 37659
rect 2296 37603 2364 37659
rect 2420 37603 2444 37659
rect 1844 37535 2444 37603
rect 1844 37479 1868 37535
rect 1924 37479 1992 37535
rect 2048 37479 2116 37535
rect 2172 37479 2240 37535
rect 2296 37479 2364 37535
rect 2420 37479 2444 37535
rect 1844 37411 2444 37479
rect 1844 37355 1868 37411
rect 1924 37355 1992 37411
rect 2048 37355 2116 37411
rect 2172 37355 2240 37411
rect 2296 37355 2364 37411
rect 2420 37355 2444 37411
rect 1844 37287 2444 37355
rect 1844 37231 1868 37287
rect 1924 37231 1992 37287
rect 2048 37231 2116 37287
rect 2172 37231 2240 37287
rect 2296 37231 2364 37287
rect 2420 37231 2444 37287
rect 1844 37163 2444 37231
rect 1844 37107 1868 37163
rect 1924 37107 1992 37163
rect 2048 37107 2116 37163
rect 2172 37107 2240 37163
rect 2296 37107 2364 37163
rect 2420 37107 2444 37163
rect 1844 20059 2444 37107
rect 1844 20003 1930 20059
rect 1986 20003 2054 20059
rect 2110 20003 2178 20059
rect 2234 20003 2302 20059
rect 2358 20003 2444 20059
rect 1844 19935 2444 20003
rect 1844 19879 1930 19935
rect 1986 19879 2054 19935
rect 2110 19879 2178 19935
rect 2234 19879 2302 19935
rect 2358 19879 2444 19935
rect 1844 19811 2444 19879
rect 1844 19755 1930 19811
rect 1986 19755 2054 19811
rect 2110 19755 2178 19811
rect 2234 19755 2302 19811
rect 2358 19755 2444 19811
rect 1844 19687 2444 19755
rect 1844 19631 1930 19687
rect 1986 19631 2054 19687
rect 2110 19631 2178 19687
rect 2234 19631 2302 19687
rect 2358 19631 2444 19687
rect 1844 17840 2444 19631
rect 1844 17784 1930 17840
rect 1986 17784 2054 17840
rect 2110 17784 2178 17840
rect 2234 17784 2302 17840
rect 2358 17784 2444 17840
rect 1844 17716 2444 17784
rect 1844 17660 1930 17716
rect 1986 17660 2054 17716
rect 2110 17660 2178 17716
rect 2234 17660 2302 17716
rect 2358 17660 2444 17716
rect 1844 16040 2444 17660
rect 1844 15984 1930 16040
rect 1986 15984 2054 16040
rect 2110 15984 2178 16040
rect 2234 15984 2302 16040
rect 2358 15984 2444 16040
rect 1844 15916 2444 15984
rect 1844 15860 1930 15916
rect 1986 15860 2054 15916
rect 2110 15860 2178 15916
rect 2234 15860 2302 15916
rect 2358 15860 2444 15916
rect 1844 14240 2444 15860
rect 1844 14184 1930 14240
rect 1986 14184 2054 14240
rect 2110 14184 2178 14240
rect 2234 14184 2302 14240
rect 2358 14184 2444 14240
rect 1844 14116 2444 14184
rect 1844 14060 1930 14116
rect 1986 14060 2054 14116
rect 2110 14060 2178 14116
rect 2234 14060 2302 14116
rect 2358 14060 2444 14116
rect 1844 12440 2444 14060
rect 1844 12384 1930 12440
rect 1986 12384 2054 12440
rect 2110 12384 2178 12440
rect 2234 12384 2302 12440
rect 2358 12384 2444 12440
rect 1844 12316 2444 12384
rect 1844 12260 1930 12316
rect 1986 12260 2054 12316
rect 2110 12260 2178 12316
rect 2234 12260 2302 12316
rect 2358 12260 2444 12316
rect 1844 10640 2444 12260
rect 1844 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2444 10640
rect 1844 10516 2444 10584
rect 1844 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2444 10516
rect 1844 8840 2444 10460
rect 1844 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2444 8840
rect 1844 8716 2444 8784
rect 1844 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2444 8716
rect 1844 7040 2444 8660
rect 1844 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2444 7040
rect 1844 6916 2444 6984
rect 1844 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2444 6916
rect 1844 5240 2444 6860
rect 1844 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2444 5240
rect 1844 5116 2444 5184
rect 1844 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2444 5116
rect 1844 3440 2444 5060
rect 1844 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2444 3440
rect 1844 3316 2444 3384
rect 1844 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2444 3316
rect 1844 3136 2444 3260
rect 85726 42689 86326 52528
rect 85726 42633 85750 42689
rect 85806 42633 85874 42689
rect 85930 42633 85998 42689
rect 86054 42633 86122 42689
rect 86178 42633 86246 42689
rect 86302 42633 86326 42689
rect 85726 42565 86326 42633
rect 85726 42509 85750 42565
rect 85806 42509 85874 42565
rect 85930 42509 85998 42565
rect 86054 42509 86122 42565
rect 86178 42509 86246 42565
rect 86302 42509 86326 42565
rect 85726 42441 86326 42509
rect 85726 42385 85750 42441
rect 85806 42385 85874 42441
rect 85930 42385 85998 42441
rect 86054 42385 86122 42441
rect 86178 42385 86246 42441
rect 86302 42385 86326 42441
rect 85726 42317 86326 42385
rect 85726 42261 85750 42317
rect 85806 42261 85874 42317
rect 85930 42261 85998 42317
rect 86054 42261 86122 42317
rect 86178 42261 86246 42317
rect 86302 42261 86326 42317
rect 85726 42193 86326 42261
rect 85726 42137 85750 42193
rect 85806 42137 85874 42193
rect 85930 42137 85998 42193
rect 86054 42137 86122 42193
rect 86178 42137 86246 42193
rect 86302 42137 86326 42193
rect 85726 42069 86326 42137
rect 85726 42013 85750 42069
rect 85806 42013 85874 42069
rect 85930 42013 85998 42069
rect 86054 42013 86122 42069
rect 86178 42013 86246 42069
rect 86302 42013 86326 42069
rect 85726 41945 86326 42013
rect 85726 41889 85750 41945
rect 85806 41889 85874 41945
rect 85930 41889 85998 41945
rect 86054 41889 86122 41945
rect 86178 41889 86246 41945
rect 86302 41889 86326 41945
rect 85726 41821 86326 41889
rect 85726 41765 85750 41821
rect 85806 41765 85874 41821
rect 85930 41765 85998 41821
rect 86054 41765 86122 41821
rect 86178 41765 86246 41821
rect 86302 41765 86326 41821
rect 85726 41697 86326 41765
rect 85726 41641 85750 41697
rect 85806 41641 85874 41697
rect 85930 41641 85998 41697
rect 86054 41641 86122 41697
rect 86178 41641 86246 41697
rect 86302 41641 86326 41697
rect 85726 41573 86326 41641
rect 85726 41517 85750 41573
rect 85806 41517 85874 41573
rect 85930 41517 85998 41573
rect 86054 41517 86122 41573
rect 86178 41517 86246 41573
rect 86302 41517 86326 41573
rect 85726 41449 86326 41517
rect 85726 41393 85750 41449
rect 85806 41393 85874 41449
rect 85930 41393 85998 41449
rect 86054 41393 86122 41449
rect 86178 41393 86246 41449
rect 86302 41393 86326 41449
rect 85726 41325 86326 41393
rect 85726 41269 85750 41325
rect 85806 41269 85874 41325
rect 85930 41269 85998 41325
rect 86054 41269 86122 41325
rect 86178 41269 86246 41325
rect 86302 41269 86326 41325
rect 85726 41201 86326 41269
rect 85726 41145 85750 41201
rect 85806 41145 85874 41201
rect 85930 41145 85998 41201
rect 86054 41145 86122 41201
rect 86178 41145 86246 41201
rect 86302 41145 86326 41201
rect 85726 41077 86326 41145
rect 85726 41021 85750 41077
rect 85806 41021 85874 41077
rect 85930 41021 85998 41077
rect 86054 41021 86122 41077
rect 86178 41021 86246 41077
rect 86302 41021 86326 41077
rect 85726 40953 86326 41021
rect 85726 40897 85750 40953
rect 85806 40897 85874 40953
rect 85930 40897 85998 40953
rect 86054 40897 86122 40953
rect 86178 40897 86246 40953
rect 86302 40897 86326 40953
rect 85726 40829 86326 40897
rect 85726 40773 85750 40829
rect 85806 40773 85874 40829
rect 85930 40773 85998 40829
rect 86054 40773 86122 40829
rect 86178 40773 86246 40829
rect 86302 40773 86326 40829
rect 85726 40705 86326 40773
rect 85726 40649 85750 40705
rect 85806 40649 85874 40705
rect 85930 40649 85998 40705
rect 86054 40649 86122 40705
rect 86178 40649 86246 40705
rect 86302 40649 86326 40705
rect 85726 31800 86326 40649
rect 85726 31744 85750 31800
rect 85806 31744 85874 31800
rect 85930 31744 85998 31800
rect 86054 31744 86122 31800
rect 86178 31744 86246 31800
rect 86302 31744 86326 31800
rect 85726 31676 86326 31744
rect 85726 31620 85750 31676
rect 85806 31620 85874 31676
rect 85930 31620 85998 31676
rect 86054 31620 86122 31676
rect 86178 31620 86246 31676
rect 86302 31620 86326 31676
rect 85726 31552 86326 31620
rect 85726 31496 85750 31552
rect 85806 31496 85874 31552
rect 85930 31496 85998 31552
rect 86054 31496 86122 31552
rect 86178 31496 86246 31552
rect 86302 31496 86326 31552
rect 85726 31428 86326 31496
rect 85726 31372 85750 31428
rect 85806 31372 85874 31428
rect 85930 31372 85998 31428
rect 86054 31372 86122 31428
rect 86178 31372 86246 31428
rect 86302 31372 86326 31428
rect 85726 31304 86326 31372
rect 85726 31248 85750 31304
rect 85806 31248 85874 31304
rect 85930 31248 85998 31304
rect 86054 31248 86122 31304
rect 86178 31248 86246 31304
rect 86302 31248 86326 31304
rect 85726 31180 86326 31248
rect 85726 31124 85750 31180
rect 85806 31124 85874 31180
rect 85930 31124 85998 31180
rect 86054 31124 86122 31180
rect 86178 31124 86246 31180
rect 86302 31124 86326 31180
rect 85726 31056 86326 31124
rect 85726 31000 85750 31056
rect 85806 31000 85874 31056
rect 85930 31000 85998 31056
rect 86054 31000 86122 31056
rect 86178 31000 86246 31056
rect 86302 31000 86326 31056
rect 85726 30932 86326 31000
rect 85726 30876 85750 30932
rect 85806 30876 85874 30932
rect 85930 30876 85998 30932
rect 86054 30876 86122 30932
rect 86178 30876 86246 30932
rect 86302 30876 86326 30932
rect 85726 18864 86326 30876
rect 85726 18808 85812 18864
rect 85868 18808 85936 18864
rect 85992 18808 86060 18864
rect 86116 18808 86184 18864
rect 86240 18808 86326 18864
rect 85726 18740 86326 18808
rect 85726 18684 85812 18740
rect 85868 18684 85936 18740
rect 85992 18684 86060 18740
rect 86116 18684 86184 18740
rect 86240 18684 86326 18740
rect 85726 18616 86326 18684
rect 85726 18560 85812 18616
rect 85868 18560 85936 18616
rect 85992 18560 86060 18616
rect 86116 18560 86184 18616
rect 86240 18560 86326 18616
rect 85726 18492 86326 18560
rect 85726 18436 85812 18492
rect 85868 18436 85936 18492
rect 85992 18436 86060 18492
rect 86116 18436 86184 18492
rect 86240 18436 86326 18492
rect 85726 17064 86326 18436
rect 85726 17008 85812 17064
rect 85868 17008 85936 17064
rect 85992 17008 86060 17064
rect 86116 17008 86184 17064
rect 86240 17008 86326 17064
rect 85726 16940 86326 17008
rect 85726 16884 85812 16940
rect 85868 16884 85936 16940
rect 85992 16884 86060 16940
rect 86116 16884 86184 16940
rect 86240 16884 86326 16940
rect 85726 16816 86326 16884
rect 85726 16760 85812 16816
rect 85868 16760 85936 16816
rect 85992 16760 86060 16816
rect 86116 16760 86184 16816
rect 86240 16760 86326 16816
rect 85726 16692 86326 16760
rect 85726 16636 85812 16692
rect 85868 16636 85936 16692
rect 85992 16636 86060 16692
rect 86116 16636 86184 16692
rect 86240 16636 86326 16692
rect 85726 15264 86326 16636
rect 85726 15208 85812 15264
rect 85868 15208 85936 15264
rect 85992 15208 86060 15264
rect 86116 15208 86184 15264
rect 86240 15208 86326 15264
rect 85726 15140 86326 15208
rect 85726 15084 85812 15140
rect 85868 15084 85936 15140
rect 85992 15084 86060 15140
rect 86116 15084 86184 15140
rect 86240 15084 86326 15140
rect 85726 15016 86326 15084
rect 85726 14960 85812 15016
rect 85868 14960 85936 15016
rect 85992 14960 86060 15016
rect 86116 14960 86184 15016
rect 86240 14960 86326 15016
rect 85726 14892 86326 14960
rect 85726 14836 85812 14892
rect 85868 14836 85936 14892
rect 85992 14836 86060 14892
rect 86116 14836 86184 14892
rect 86240 14836 86326 14892
rect 85726 13464 86326 14836
rect 85726 13408 85812 13464
rect 85868 13408 85936 13464
rect 85992 13408 86060 13464
rect 86116 13408 86184 13464
rect 86240 13408 86326 13464
rect 85726 13340 86326 13408
rect 85726 13284 85812 13340
rect 85868 13284 85936 13340
rect 85992 13284 86060 13340
rect 86116 13284 86184 13340
rect 86240 13284 86326 13340
rect 85726 13216 86326 13284
rect 85726 13160 85812 13216
rect 85868 13160 85936 13216
rect 85992 13160 86060 13216
rect 86116 13160 86184 13216
rect 86240 13160 86326 13216
rect 85726 13092 86326 13160
rect 85726 13036 85812 13092
rect 85868 13036 85936 13092
rect 85992 13036 86060 13092
rect 86116 13036 86184 13092
rect 86240 13036 86326 13092
rect 85726 11664 86326 13036
rect 85726 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86326 11664
rect 85726 11540 86326 11608
rect 85726 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86326 11540
rect 85726 11416 86326 11484
rect 85726 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86326 11416
rect 85726 11292 86326 11360
rect 85726 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86326 11292
rect 85726 9864 86326 11236
rect 85726 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86326 9864
rect 85726 9740 86326 9808
rect 85726 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86326 9740
rect 85726 9616 86326 9684
rect 85726 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86326 9616
rect 85726 9492 86326 9560
rect 85726 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86326 9492
rect 85726 8064 86326 9436
rect 85726 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86326 8064
rect 85726 7940 86326 8008
rect 85726 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86326 7940
rect 85726 7816 86326 7884
rect 85726 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86326 7816
rect 85726 7692 86326 7760
rect 85726 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86326 7692
rect 85726 6264 86326 7636
rect 85726 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86326 6264
rect 85726 6140 86326 6208
rect 85726 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86326 6140
rect 85726 6016 86326 6084
rect 85726 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86326 6016
rect 85726 5892 86326 5960
rect 85726 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86326 5892
rect 85726 4464 86326 5836
rect 85726 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86326 4464
rect 85726 4340 86326 4408
rect 85726 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86326 4340
rect 85726 4216 86326 4284
rect 85726 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86326 4216
rect 85726 4092 86326 4160
rect 85726 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86326 4092
rect 85726 3136 86326 4036
rect 86526 52225 87126 52528
rect 86526 52169 86550 52225
rect 86606 52169 86674 52225
rect 86730 52169 86798 52225
rect 86854 52169 86922 52225
rect 86978 52169 87046 52225
rect 87102 52169 87126 52225
rect 86526 52101 87126 52169
rect 86526 52045 86550 52101
rect 86606 52045 86674 52101
rect 86730 52045 86798 52101
rect 86854 52045 86922 52101
rect 86978 52045 87046 52101
rect 87102 52045 87126 52101
rect 86526 51977 87126 52045
rect 86526 51921 86550 51977
rect 86606 51921 86674 51977
rect 86730 51921 86798 51977
rect 86854 51921 86922 51977
rect 86978 51921 87046 51977
rect 87102 51921 87126 51977
rect 86526 51853 87126 51921
rect 86526 51797 86550 51853
rect 86606 51797 86674 51853
rect 86730 51797 86798 51853
rect 86854 51797 86922 51853
rect 86978 51797 87046 51853
rect 87102 51797 87126 51853
rect 86526 51729 87126 51797
rect 86526 51673 86550 51729
rect 86606 51673 86674 51729
rect 86730 51673 86798 51729
rect 86854 51673 86922 51729
rect 86978 51673 87046 51729
rect 87102 51673 87126 51729
rect 86526 51605 87126 51673
rect 86526 51549 86550 51605
rect 86606 51549 86674 51605
rect 86730 51549 86798 51605
rect 86854 51549 86922 51605
rect 86978 51549 87046 51605
rect 87102 51549 87126 51605
rect 86526 51481 87126 51549
rect 86526 51425 86550 51481
rect 86606 51425 86674 51481
rect 86730 51425 86798 51481
rect 86854 51425 86922 51481
rect 86978 51425 87046 51481
rect 87102 51425 87126 51481
rect 86526 51357 87126 51425
rect 86526 51301 86550 51357
rect 86606 51301 86674 51357
rect 86730 51301 86798 51357
rect 86854 51301 86922 51357
rect 86978 51301 87046 51357
rect 87102 51301 87126 51357
rect 86526 51233 87126 51301
rect 86526 51177 86550 51233
rect 86606 51177 86674 51233
rect 86730 51177 86798 51233
rect 86854 51177 86922 51233
rect 86978 51177 87046 51233
rect 87102 51177 87126 51233
rect 86526 51109 87126 51177
rect 86526 51053 86550 51109
rect 86606 51053 86674 51109
rect 86730 51053 86798 51109
rect 86854 51053 86922 51109
rect 86978 51053 87046 51109
rect 87102 51053 87126 51109
rect 86526 48991 87126 51053
rect 86526 48935 86550 48991
rect 86606 48935 86674 48991
rect 86730 48935 86798 48991
rect 86854 48935 86922 48991
rect 86978 48935 87046 48991
rect 87102 48935 87126 48991
rect 86526 48867 87126 48935
rect 86526 48811 86550 48867
rect 86606 48811 86674 48867
rect 86730 48811 86798 48867
rect 86854 48811 86922 48867
rect 86978 48811 87046 48867
rect 87102 48811 87126 48867
rect 86526 48743 87126 48811
rect 86526 48687 86550 48743
rect 86606 48687 86674 48743
rect 86730 48687 86798 48743
rect 86854 48687 86922 48743
rect 86978 48687 87046 48743
rect 87102 48687 87126 48743
rect 86526 48619 87126 48687
rect 86526 48563 86550 48619
rect 86606 48563 86674 48619
rect 86730 48563 86798 48619
rect 86854 48563 86922 48619
rect 86978 48563 87046 48619
rect 87102 48563 87126 48619
rect 86526 48495 87126 48563
rect 86526 48439 86550 48495
rect 86606 48439 86674 48495
rect 86730 48439 86798 48495
rect 86854 48439 86922 48495
rect 86978 48439 87046 48495
rect 87102 48439 87126 48495
rect 86526 48371 87126 48439
rect 86526 48315 86550 48371
rect 86606 48315 86674 48371
rect 86730 48315 86798 48371
rect 86854 48315 86922 48371
rect 86978 48315 87046 48371
rect 87102 48315 87126 48371
rect 86526 48247 87126 48315
rect 86526 48191 86550 48247
rect 86606 48191 86674 48247
rect 86730 48191 86798 48247
rect 86854 48191 86922 48247
rect 86978 48191 87046 48247
rect 87102 48191 87126 48247
rect 86526 48123 87126 48191
rect 86526 48067 86550 48123
rect 86606 48067 86674 48123
rect 86730 48067 86798 48123
rect 86854 48067 86922 48123
rect 86978 48067 87046 48123
rect 87102 48067 87126 48123
rect 86526 47999 87126 48067
rect 86526 47943 86550 47999
rect 86606 47943 86674 47999
rect 86730 47943 86798 47999
rect 86854 47943 86922 47999
rect 86978 47943 87046 47999
rect 87102 47943 87126 47999
rect 86526 47875 87126 47943
rect 86526 47819 86550 47875
rect 86606 47819 86674 47875
rect 86730 47819 86798 47875
rect 86854 47819 86922 47875
rect 86978 47819 87046 47875
rect 87102 47819 87126 47875
rect 86526 47751 87126 47819
rect 86526 47695 86550 47751
rect 86606 47695 86674 47751
rect 86730 47695 86798 47751
rect 86854 47695 86922 47751
rect 86978 47695 87046 47751
rect 87102 47695 87126 47751
rect 86526 47627 87126 47695
rect 86526 47571 86550 47627
rect 86606 47571 86674 47627
rect 86730 47571 86798 47627
rect 86854 47571 86922 47627
rect 86978 47571 87046 47627
rect 87102 47571 87126 47627
rect 86526 47503 87126 47571
rect 86526 47447 86550 47503
rect 86606 47447 86674 47503
rect 86730 47447 86798 47503
rect 86854 47447 86922 47503
rect 86978 47447 87046 47503
rect 87102 47447 87126 47503
rect 86526 47379 87126 47447
rect 86526 47323 86550 47379
rect 86606 47323 86674 47379
rect 86730 47323 86798 47379
rect 86854 47323 86922 47379
rect 86978 47323 87046 47379
rect 87102 47323 87126 47379
rect 86526 47255 87126 47323
rect 86526 47199 86550 47255
rect 86606 47199 86674 47255
rect 86730 47199 86798 47255
rect 86854 47199 86922 47255
rect 86978 47199 87046 47255
rect 87102 47199 87126 47255
rect 86526 40387 87126 47199
rect 86526 40331 86550 40387
rect 86606 40331 86674 40387
rect 86730 40331 86798 40387
rect 86854 40331 86922 40387
rect 86978 40331 87046 40387
rect 87102 40331 87126 40387
rect 86526 40263 87126 40331
rect 86526 40207 86550 40263
rect 86606 40207 86674 40263
rect 86730 40207 86798 40263
rect 86854 40207 86922 40263
rect 86978 40207 87046 40263
rect 87102 40207 87126 40263
rect 86526 40139 87126 40207
rect 86526 40083 86550 40139
rect 86606 40083 86674 40139
rect 86730 40083 86798 40139
rect 86854 40083 86922 40139
rect 86978 40083 87046 40139
rect 87102 40083 87126 40139
rect 86526 40015 87126 40083
rect 86526 39959 86550 40015
rect 86606 39959 86674 40015
rect 86730 39959 86798 40015
rect 86854 39959 86922 40015
rect 86978 39959 87046 40015
rect 87102 39959 87126 40015
rect 86526 39891 87126 39959
rect 86526 39835 86550 39891
rect 86606 39835 86674 39891
rect 86730 39835 86798 39891
rect 86854 39835 86922 39891
rect 86978 39835 87046 39891
rect 87102 39835 87126 39891
rect 86526 39767 87126 39835
rect 86526 39711 86550 39767
rect 86606 39711 86674 39767
rect 86730 39711 86798 39767
rect 86854 39711 86922 39767
rect 86978 39711 87046 39767
rect 87102 39711 87126 39767
rect 86526 39643 87126 39711
rect 86526 39587 86550 39643
rect 86606 39587 86674 39643
rect 86730 39587 86798 39643
rect 86854 39587 86922 39643
rect 86978 39587 87046 39643
rect 87102 39587 87126 39643
rect 86526 39519 87126 39587
rect 86526 39463 86550 39519
rect 86606 39463 86674 39519
rect 86730 39463 86798 39519
rect 86854 39463 86922 39519
rect 86978 39463 87046 39519
rect 87102 39463 87126 39519
rect 86526 39395 87126 39463
rect 86526 39339 86550 39395
rect 86606 39339 86674 39395
rect 86730 39339 86798 39395
rect 86854 39339 86922 39395
rect 86978 39339 87046 39395
rect 87102 39339 87126 39395
rect 86526 39271 87126 39339
rect 86526 39215 86550 39271
rect 86606 39215 86674 39271
rect 86730 39215 86798 39271
rect 86854 39215 86922 39271
rect 86978 39215 87046 39271
rect 87102 39215 87126 39271
rect 86526 39147 87126 39215
rect 86526 39091 86550 39147
rect 86606 39091 86674 39147
rect 86730 39091 86798 39147
rect 86854 39091 86922 39147
rect 86978 39091 87046 39147
rect 87102 39091 87126 39147
rect 86526 39023 87126 39091
rect 86526 38967 86550 39023
rect 86606 38967 86674 39023
rect 86730 38967 86798 39023
rect 86854 38967 86922 39023
rect 86978 38967 87046 39023
rect 87102 38967 87126 39023
rect 86526 38899 87126 38967
rect 86526 38843 86550 38899
rect 86606 38843 86674 38899
rect 86730 38843 86798 38899
rect 86854 38843 86922 38899
rect 86978 38843 87046 38899
rect 87102 38843 87126 38899
rect 86526 38775 87126 38843
rect 86526 38719 86550 38775
rect 86606 38719 86674 38775
rect 86730 38719 86798 38775
rect 86854 38719 86922 38775
rect 86978 38719 87046 38775
rect 87102 38719 87126 38775
rect 86526 38651 87126 38719
rect 86526 38595 86550 38651
rect 86606 38595 86674 38651
rect 86730 38595 86798 38651
rect 86854 38595 86922 38651
rect 86978 38595 87046 38651
rect 87102 38595 87126 38651
rect 86526 38527 87126 38595
rect 86526 38471 86550 38527
rect 86606 38471 86674 38527
rect 86730 38471 86798 38527
rect 86854 38471 86922 38527
rect 86978 38471 87046 38527
rect 87102 38471 87126 38527
rect 86526 38403 87126 38471
rect 86526 38347 86550 38403
rect 86606 38347 86674 38403
rect 86730 38347 86798 38403
rect 86854 38347 86922 38403
rect 86978 38347 87046 38403
rect 87102 38347 87126 38403
rect 86526 38279 87126 38347
rect 86526 38223 86550 38279
rect 86606 38223 86674 38279
rect 86730 38223 86798 38279
rect 86854 38223 86922 38279
rect 86978 38223 87046 38279
rect 87102 38223 87126 38279
rect 86526 38155 87126 38223
rect 86526 38099 86550 38155
rect 86606 38099 86674 38155
rect 86730 38099 86798 38155
rect 86854 38099 86922 38155
rect 86978 38099 87046 38155
rect 87102 38099 87126 38155
rect 86526 38031 87126 38099
rect 86526 37975 86550 38031
rect 86606 37975 86674 38031
rect 86730 37975 86798 38031
rect 86854 37975 86922 38031
rect 86978 37975 87046 38031
rect 87102 37975 87126 38031
rect 86526 37907 87126 37975
rect 86526 37851 86550 37907
rect 86606 37851 86674 37907
rect 86730 37851 86798 37907
rect 86854 37851 86922 37907
rect 86978 37851 87046 37907
rect 87102 37851 87126 37907
rect 86526 37783 87126 37851
rect 86526 37727 86550 37783
rect 86606 37727 86674 37783
rect 86730 37727 86798 37783
rect 86854 37727 86922 37783
rect 86978 37727 87046 37783
rect 87102 37727 87126 37783
rect 86526 37659 87126 37727
rect 86526 37603 86550 37659
rect 86606 37603 86674 37659
rect 86730 37603 86798 37659
rect 86854 37603 86922 37659
rect 86978 37603 87046 37659
rect 87102 37603 87126 37659
rect 86526 37535 87126 37603
rect 86526 37479 86550 37535
rect 86606 37479 86674 37535
rect 86730 37479 86798 37535
rect 86854 37479 86922 37535
rect 86978 37479 87046 37535
rect 87102 37479 87126 37535
rect 86526 37411 87126 37479
rect 86526 37355 86550 37411
rect 86606 37355 86674 37411
rect 86730 37355 86798 37411
rect 86854 37355 86922 37411
rect 86978 37355 87046 37411
rect 87102 37355 87126 37411
rect 86526 37287 87126 37355
rect 86526 37231 86550 37287
rect 86606 37231 86674 37287
rect 86730 37231 86798 37287
rect 86854 37231 86922 37287
rect 86978 37231 87046 37287
rect 87102 37231 87126 37287
rect 86526 37163 87126 37231
rect 86526 37107 86550 37163
rect 86606 37107 86674 37163
rect 86730 37107 86798 37163
rect 86854 37107 86922 37163
rect 86978 37107 87046 37163
rect 87102 37107 87126 37163
rect 86526 33456 87126 37107
rect 86526 33400 86550 33456
rect 86606 33400 86674 33456
rect 86730 33400 86798 33456
rect 86854 33400 86922 33456
rect 86978 33400 87046 33456
rect 87102 33400 87126 33456
rect 86526 33332 87126 33400
rect 86526 33276 86550 33332
rect 86606 33276 86674 33332
rect 86730 33276 86798 33332
rect 86854 33276 86922 33332
rect 86978 33276 87046 33332
rect 87102 33276 87126 33332
rect 86526 33208 87126 33276
rect 86526 33152 86550 33208
rect 86606 33152 86674 33208
rect 86730 33152 86798 33208
rect 86854 33152 86922 33208
rect 86978 33152 87046 33208
rect 87102 33152 87126 33208
rect 86526 33084 87126 33152
rect 86526 33028 86550 33084
rect 86606 33028 86674 33084
rect 86730 33028 86798 33084
rect 86854 33028 86922 33084
rect 86978 33028 87046 33084
rect 87102 33028 87126 33084
rect 86526 32960 87126 33028
rect 86526 32904 86550 32960
rect 86606 32904 86674 32960
rect 86730 32904 86798 32960
rect 86854 32904 86922 32960
rect 86978 32904 87046 32960
rect 87102 32904 87126 32960
rect 86526 32836 87126 32904
rect 86526 32780 86550 32836
rect 86606 32780 86674 32836
rect 86730 32780 86798 32836
rect 86854 32780 86922 32836
rect 86978 32780 87046 32836
rect 87102 32780 87126 32836
rect 86526 32712 87126 32780
rect 86526 32656 86550 32712
rect 86606 32656 86674 32712
rect 86730 32656 86798 32712
rect 86854 32656 86922 32712
rect 86978 32656 87046 32712
rect 87102 32656 87126 32712
rect 86526 32588 87126 32656
rect 86526 32532 86550 32588
rect 86606 32532 86674 32588
rect 86730 32532 86798 32588
rect 86854 32532 86922 32588
rect 86978 32532 87046 32588
rect 87102 32532 87126 32588
rect 86526 20059 87126 32532
rect 86526 20003 86612 20059
rect 86668 20003 86736 20059
rect 86792 20003 86860 20059
rect 86916 20003 86984 20059
rect 87040 20003 87126 20059
rect 86526 19935 87126 20003
rect 86526 19879 86612 19935
rect 86668 19879 86736 19935
rect 86792 19879 86860 19935
rect 86916 19879 86984 19935
rect 87040 19879 87126 19935
rect 86526 19811 87126 19879
rect 86526 19755 86612 19811
rect 86668 19755 86736 19811
rect 86792 19755 86860 19811
rect 86916 19755 86984 19811
rect 87040 19755 87126 19811
rect 86526 19687 87126 19755
rect 86526 19631 86612 19687
rect 86668 19631 86736 19687
rect 86792 19631 86860 19687
rect 86916 19631 86984 19687
rect 87040 19631 87126 19687
rect 86526 17964 87126 19631
rect 86526 17908 86612 17964
rect 86668 17908 86736 17964
rect 86792 17908 86860 17964
rect 86916 17908 86984 17964
rect 87040 17908 87126 17964
rect 86526 17840 87126 17908
rect 86526 17784 86612 17840
rect 86668 17784 86736 17840
rect 86792 17784 86860 17840
rect 86916 17784 86984 17840
rect 87040 17784 87126 17840
rect 86526 17716 87126 17784
rect 86526 17660 86612 17716
rect 86668 17660 86736 17716
rect 86792 17660 86860 17716
rect 86916 17660 86984 17716
rect 87040 17660 87126 17716
rect 86526 17592 87126 17660
rect 86526 17536 86612 17592
rect 86668 17536 86736 17592
rect 86792 17536 86860 17592
rect 86916 17536 86984 17592
rect 87040 17536 87126 17592
rect 86526 16164 87126 17536
rect 86526 16108 86612 16164
rect 86668 16108 86736 16164
rect 86792 16108 86860 16164
rect 86916 16108 86984 16164
rect 87040 16108 87126 16164
rect 86526 16040 87126 16108
rect 86526 15984 86612 16040
rect 86668 15984 86736 16040
rect 86792 15984 86860 16040
rect 86916 15984 86984 16040
rect 87040 15984 87126 16040
rect 86526 15916 87126 15984
rect 86526 15860 86612 15916
rect 86668 15860 86736 15916
rect 86792 15860 86860 15916
rect 86916 15860 86984 15916
rect 87040 15860 87126 15916
rect 86526 15792 87126 15860
rect 86526 15736 86612 15792
rect 86668 15736 86736 15792
rect 86792 15736 86860 15792
rect 86916 15736 86984 15792
rect 87040 15736 87126 15792
rect 86526 14364 87126 15736
rect 86526 14308 86612 14364
rect 86668 14308 86736 14364
rect 86792 14308 86860 14364
rect 86916 14308 86984 14364
rect 87040 14308 87126 14364
rect 86526 14240 87126 14308
rect 86526 14184 86612 14240
rect 86668 14184 86736 14240
rect 86792 14184 86860 14240
rect 86916 14184 86984 14240
rect 87040 14184 87126 14240
rect 86526 14116 87126 14184
rect 86526 14060 86612 14116
rect 86668 14060 86736 14116
rect 86792 14060 86860 14116
rect 86916 14060 86984 14116
rect 87040 14060 87126 14116
rect 86526 13992 87126 14060
rect 86526 13936 86612 13992
rect 86668 13936 86736 13992
rect 86792 13936 86860 13992
rect 86916 13936 86984 13992
rect 87040 13936 87126 13992
rect 86526 12564 87126 13936
rect 86526 12508 86612 12564
rect 86668 12508 86736 12564
rect 86792 12508 86860 12564
rect 86916 12508 86984 12564
rect 87040 12508 87126 12564
rect 86526 12440 87126 12508
rect 86526 12384 86612 12440
rect 86668 12384 86736 12440
rect 86792 12384 86860 12440
rect 86916 12384 86984 12440
rect 87040 12384 87126 12440
rect 86526 12316 87126 12384
rect 86526 12260 86612 12316
rect 86668 12260 86736 12316
rect 86792 12260 86860 12316
rect 86916 12260 86984 12316
rect 87040 12260 87126 12316
rect 86526 12192 87126 12260
rect 86526 12136 86612 12192
rect 86668 12136 86736 12192
rect 86792 12136 86860 12192
rect 86916 12136 86984 12192
rect 87040 12136 87126 12192
rect 86526 10764 87126 12136
rect 86526 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87126 10764
rect 86526 10640 87126 10708
rect 86526 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87126 10640
rect 86526 10516 87126 10584
rect 86526 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87126 10516
rect 86526 10392 87126 10460
rect 86526 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87126 10392
rect 86526 8964 87126 10336
rect 86526 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87126 8964
rect 86526 8840 87126 8908
rect 86526 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87126 8840
rect 86526 8716 87126 8784
rect 86526 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87126 8716
rect 86526 8592 87126 8660
rect 86526 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87126 8592
rect 86526 7164 87126 8536
rect 86526 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87126 7164
rect 86526 7040 87126 7108
rect 86526 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87126 7040
rect 86526 6916 87126 6984
rect 86526 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87126 6916
rect 86526 6792 87126 6860
rect 86526 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87126 6792
rect 86526 5364 87126 6736
rect 86526 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87126 5364
rect 86526 5240 87126 5308
rect 86526 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87126 5240
rect 86526 5116 87126 5184
rect 86526 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87126 5116
rect 86526 4992 87126 5060
rect 86526 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87126 4992
rect 86526 3632 87126 4936
rect 86526 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87126 3632
rect 86526 3508 87126 3576
rect 86526 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87126 3508
rect 86526 3384 87126 3452
rect 86526 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87126 3384
rect 86526 3260 87126 3328
rect 86526 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87126 3260
rect 86526 3136 87126 3204
use gf180mcu_fd_ip_sram__sram128x8m8wm1  RAM
timestamp 0
transform -1 0 87372 0 -1 54776
box 0 0 86372 53776
<< labels >>
flabel metal2 s 52944 55176 53056 55976 0 FreeSans 448 90 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 54644 55176 54756 55976 0 FreeSans 448 90 0 0 A[1]
port 1 nsew signal input
flabel metal2 s 56344 55176 56456 55976 0 FreeSans 448 90 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 30944 55176 31056 55976 0 FreeSans 448 90 0 0 A[3]
port 3 nsew signal input
flabel metal2 s 31944 55176 32056 55976 0 FreeSans 448 90 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 32744 55176 32856 55976 0 FreeSans 448 90 0 0 A[5]
port 5 nsew signal input
flabel metal2 s 33344 55176 33456 55976 0 FreeSans 448 90 0 0 A[6]
port 6 nsew signal input
flabel metal2 s 36844 55176 36956 55976 0 FreeSans 448 90 0 0 CEN
port 7 nsew signal input
flabel metal2 s 59244 55176 59356 55976 0 FreeSans 448 90 0 0 CLK
port 8 nsew signal input
flabel metal2 s 85344 55176 85456 55976 0 FreeSans 448 90 0 0 D[0]
port 9 nsew signal input
flabel metal2 s 74944 55176 75056 55976 0 FreeSans 448 90 0 0 D[1]
port 10 nsew signal input
flabel metal2 s 73744 55176 73856 55976 0 FreeSans 448 90 0 0 D[2]
port 11 nsew signal input
flabel metal2 s 63344 55176 63456 55976 0 FreeSans 448 90 0 0 D[3]
port 12 nsew signal input
flabel metal2 s 25744 55176 25856 55976 0 FreeSans 448 90 0 0 D[4]
port 13 nsew signal input
flabel metal2 s 15444 55176 15556 55976 0 FreeSans 448 90 0 0 D[5]
port 14 nsew signal input
flabel metal2 s 14144 55176 14256 55976 0 FreeSans 448 90 0 0 D[6]
port 15 nsew signal input
flabel metal2 s 3744 55176 3856 55976 0 FreeSans 448 90 0 0 D[7]
port 16 nsew signal input
flabel metal2 s 46568 55176 46680 55976 0 FreeSans 448 90 0 0 GWEN
port 17 nsew signal input
flabel metal2 s 83844 55176 83956 55976 0 FreeSans 448 90 0 0 Q[0]
port 18 nsew signal tristate
flabel metal2 s 75644 55176 75756 55976 0 FreeSans 448 90 0 0 Q[1]
port 19 nsew signal tristate
flabel metal2 s 73044 55176 73156 55976 0 FreeSans 448 90 0 0 Q[2]
port 20 nsew signal tristate
flabel metal2 s 64944 55176 65056 55976 0 FreeSans 448 90 0 0 Q[3]
port 21 nsew signal tristate
flabel metal2 s 24244 55176 24356 55976 0 FreeSans 448 90 0 0 Q[4]
port 22 nsew signal tristate
flabel metal2 s 16044 55176 16156 55976 0 FreeSans 448 90 0 0 Q[5]
port 23 nsew signal tristate
flabel metal2 s 13444 55176 13556 55976 0 FreeSans 448 90 0 0 Q[6]
port 24 nsew signal tristate
flabel metal2 s 5344 55176 5456 55976 0 FreeSans 448 90 0 0 Q[7]
port 25 nsew signal tristate
flabel metal4 s 1044 3136 1644 52528 0 FreeSans 2560 90 0 0 VDD
port 26 nsew power bidirectional
flabel metal4 s 85726 3136 86326 52528 0 FreeSans 2560 90 0 0 VDD
port 26 nsew power bidirectional
flabel metal4 s 1844 3136 2444 52528 0 FreeSans 2560 90 0 0 VSS
port 27 nsew ground bidirectional
flabel metal4 s 86526 3136 87126 52528 0 FreeSans 2560 90 0 0 VSS
port 27 nsew ground bidirectional
flabel metal2 s 84644 55176 84756 55976 0 FreeSans 448 90 0 0 WEN[0]
port 28 nsew signal input
flabel metal2 s 74544 55176 74656 55976 0 FreeSans 448 90 0 0 WEN[1]
port 29 nsew signal input
flabel metal2 s 74144 55176 74256 55976 0 FreeSans 448 90 0 0 WEN[2]
port 30 nsew signal input
flabel metal2 s 63744 55176 63856 55976 0 FreeSans 448 90 0 0 WEN[3]
port 31 nsew signal input
flabel metal2 s 25044 55176 25156 55976 0 FreeSans 448 90 0 0 WEN[4]
port 32 nsew signal input
flabel metal2 s 14994 55176 15106 55976 0 FreeSans 448 90 0 0 WEN[5]
port 33 nsew signal input
flabel metal2 s 14544 55176 14656 55976 0 FreeSans 448 90 0 0 WEN[6]
port 34 nsew signal input
flabel metal2 s 4444 55176 4556 55976 0 FreeSans 448 90 0 0 WEN[7]
port 35 nsew signal input
rlabel via3 86274 42661 86274 42661 0 VDD
rlabel via3 87074 52197 87074 52197 0 VSS
rlabel metal2 53032 54992 53032 54992 0 A[0]
rlabel metal2 54712 54992 54712 54992 0 A[1]
rlabel metal2 56392 54992 56392 54992 0 A[2]
rlabel metal2 30968 54992 30968 54992 0 A[3]
rlabel metal2 32032 54838 32032 54838 0 A[4]
rlabel metal2 32760 54992 32760 54992 0 A[5]
rlabel metal2 33432 54992 33432 54992 0 A[6]
rlabel metal2 36904 54992 36904 54992 0 CEN
rlabel metal2 59304 54992 59304 54992 0 CLK
rlabel metal2 85400 54992 85400 54992 0 D[0]
rlabel metal2 74984 54992 74984 54992 0 D[1]
rlabel metal2 73752 54992 73752 54992 0 D[2]
rlabel metal2 63448 54992 63448 54992 0 D[3]
rlabel metal2 25816 54992 25816 54992 0 D[4]
rlabel metal2 15512 54992 15512 54992 0 D[5]
rlabel metal2 14168 54992 14168 54992 0 D[6]
rlabel metal2 3808 54838 3808 54838 0 D[7]
rlabel metal2 46648 54992 46648 54992 0 GWEN
rlabel metal2 83944 54992 83944 54992 0 Q[0]
rlabel metal2 75656 54992 75656 54992 0 Q[1]
rlabel metal2 73080 54992 73080 54992 0 Q[2]
rlabel metal2 65016 54992 65016 54992 0 Q[3]
rlabel metal2 24248 54992 24248 54992 0 Q[4]
rlabel metal2 16072 54992 16072 54992 0 Q[5]
rlabel metal2 13496 54992 13496 54992 0 Q[6]
rlabel metal2 5432 54992 5432 54992 0 Q[7]
rlabel metal2 84728 54992 84728 54992 0 WEN[0]
rlabel metal2 74648 54992 74648 54992 0 WEN[1]
rlabel metal2 74200 54992 74200 54992 0 WEN[2]
rlabel metal2 63784 54992 63784 54992 0 WEN[3]
rlabel metal2 25144 54992 25144 54992 0 WEN[4]
rlabel metal2 15064 54992 15064 54992 0 WEN[5]
rlabel metal2 14616 54992 14616 54992 0 WEN[6]
rlabel metal2 4536 54992 4536 54992 0 WEN[7]
<< properties >>
string FIXED_BBOX 0 0 88972 55976
<< end >>
