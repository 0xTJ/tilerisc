VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO interp_tri
  CLASS BLOCK ;
  FOREIGN interp_tri ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 196.000 283.920 200.000 ;
    END
  END clk
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 41.685 15.380 43.285 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 113.220 15.380 114.820 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 184.755 15.380 186.355 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 256.290 15.380 257.890 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 77.450 15.380 79.050 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 148.985 15.380 150.585 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 220.520 15.380 222.120 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 292.055 15.380 293.655 184.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 4.000 113.680 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 4.000 102.480 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.320 4.000 96.880 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 4.000 80.080 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 4.000 68.880 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 62.720 4.000 63.280 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 4.000 46.480 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 4.000 35.280 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.920 4.000 18.480 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.320 4.000 12.880 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 4.000 169.680 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.520 4.000 164.080 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 4.000 147.280 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 4.000 136.080 ;
    END
  END wbs_dat_i[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END wbs_we_i
  PIN x_end[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 196.000 93.520 200.000 ;
    END
  END x_end[0]
  PIN x_end[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 196.000 82.320 200.000 ;
    END
  END x_end[1]
  PIN x_end[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 196.000 71.120 200.000 ;
    END
  END x_end[2]
  PIN x_end[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 196.000 59.920 200.000 ;
    END
  END x_end[3]
  PIN x_end[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 196.000 48.720 200.000 ;
    END
  END x_end[4]
  PIN x_end[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 196.000 37.520 200.000 ;
    END
  END x_end[5]
  PIN x_end[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 196.000 26.320 200.000 ;
    END
  END x_end[6]
  PIN x_end[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 196.000 15.120 200.000 ;
    END
  END x_end[7]
  PIN x_start[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 196.000 183.120 200.000 ;
    END
  END x_start[0]
  PIN x_start[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 196.000 171.920 200.000 ;
    END
  END x_start[1]
  PIN x_start[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 196.000 160.720 200.000 ;
    END
  END x_start[2]
  PIN x_start[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 196.000 149.520 200.000 ;
    END
  END x_start[3]
  PIN x_start[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 196.000 138.320 200.000 ;
    END
  END x_start[4]
  PIN x_start[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 196.000 127.120 200.000 ;
    END
  END x_start[5]
  PIN x_start[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 196.000 115.920 200.000 ;
    END
  END x_start[6]
  PIN x_start[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 196.000 104.720 200.000 ;
    END
  END x_start[7]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 196.000 272.720 200.000 ;
    END
  END y[0]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 196.000 261.520 200.000 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 196.000 250.320 200.000 ;
    END
  END y[2]
  PIN y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 196.000 239.120 200.000 ;
    END
  END y[3]
  PIN y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 196.000 227.920 200.000 ;
    END
  END y[4]
  PIN y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 196.000 216.720 200.000 ;
    END
  END y[5]
  PIN y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 196.000 205.520 200.000 ;
    END
  END y[6]
  PIN y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 196.000 194.320 200.000 ;
    END
  END y[7]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 293.655 184.540 ;
      LAYER Metal2 ;
        RECT 5.180 195.700 14.260 196.420 ;
        RECT 15.420 195.700 25.460 196.420 ;
        RECT 26.620 195.700 36.660 196.420 ;
        RECT 37.820 195.700 47.860 196.420 ;
        RECT 49.020 195.700 59.060 196.420 ;
        RECT 60.220 195.700 70.260 196.420 ;
        RECT 71.420 195.700 81.460 196.420 ;
        RECT 82.620 195.700 92.660 196.420 ;
        RECT 93.820 195.700 103.860 196.420 ;
        RECT 105.020 195.700 115.060 196.420 ;
        RECT 116.220 195.700 126.260 196.420 ;
        RECT 127.420 195.700 137.460 196.420 ;
        RECT 138.620 195.700 148.660 196.420 ;
        RECT 149.820 195.700 159.860 196.420 ;
        RECT 161.020 195.700 171.060 196.420 ;
        RECT 172.220 195.700 182.260 196.420 ;
        RECT 183.420 195.700 193.460 196.420 ;
        RECT 194.620 195.700 204.660 196.420 ;
        RECT 205.820 195.700 215.860 196.420 ;
        RECT 217.020 195.700 227.060 196.420 ;
        RECT 228.220 195.700 238.260 196.420 ;
        RECT 239.420 195.700 249.460 196.420 ;
        RECT 250.620 195.700 260.660 196.420 ;
        RECT 261.820 195.700 271.860 196.420 ;
        RECT 273.020 195.700 283.060 196.420 ;
        RECT 284.220 195.700 293.515 196.420 ;
        RECT 5.180 4.300 293.515 195.700 ;
        RECT 5.180 4.000 13.140 4.300 ;
        RECT 14.300 4.000 37.780 4.300 ;
        RECT 38.940 4.000 62.420 4.300 ;
        RECT 63.580 4.000 87.060 4.300 ;
        RECT 88.220 4.000 111.700 4.300 ;
        RECT 112.860 4.000 136.340 4.300 ;
        RECT 137.500 4.000 160.980 4.300 ;
        RECT 162.140 4.000 185.620 4.300 ;
        RECT 186.780 4.000 210.260 4.300 ;
        RECT 211.420 4.000 234.900 4.300 ;
        RECT 236.060 4.000 259.540 4.300 ;
        RECT 260.700 4.000 284.180 4.300 ;
        RECT 285.340 4.000 293.515 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 186.780 293.565 186.900 ;
        RECT 4.300 185.620 293.565 186.780 ;
        RECT 3.500 181.180 293.565 185.620 ;
        RECT 4.300 180.020 293.565 181.180 ;
        RECT 3.500 175.580 293.565 180.020 ;
        RECT 4.300 174.420 293.565 175.580 ;
        RECT 3.500 169.980 293.565 174.420 ;
        RECT 4.300 168.820 293.565 169.980 ;
        RECT 3.500 164.380 293.565 168.820 ;
        RECT 4.300 163.220 293.565 164.380 ;
        RECT 3.500 158.780 293.565 163.220 ;
        RECT 4.300 157.620 293.565 158.780 ;
        RECT 3.500 153.180 293.565 157.620 ;
        RECT 4.300 152.020 293.565 153.180 ;
        RECT 3.500 147.580 293.565 152.020 ;
        RECT 4.300 146.420 293.565 147.580 ;
        RECT 3.500 141.980 293.565 146.420 ;
        RECT 4.300 140.820 293.565 141.980 ;
        RECT 3.500 136.380 293.565 140.820 ;
        RECT 4.300 135.220 293.565 136.380 ;
        RECT 3.500 130.780 293.565 135.220 ;
        RECT 4.300 129.620 293.565 130.780 ;
        RECT 3.500 125.180 293.565 129.620 ;
        RECT 4.300 124.020 293.565 125.180 ;
        RECT 3.500 119.580 293.565 124.020 ;
        RECT 4.300 118.420 293.565 119.580 ;
        RECT 3.500 113.980 293.565 118.420 ;
        RECT 4.300 112.820 293.565 113.980 ;
        RECT 3.500 108.380 293.565 112.820 ;
        RECT 4.300 107.220 293.565 108.380 ;
        RECT 3.500 102.780 293.565 107.220 ;
        RECT 4.300 101.620 293.565 102.780 ;
        RECT 3.500 97.180 293.565 101.620 ;
        RECT 4.300 96.020 293.565 97.180 ;
        RECT 3.500 91.580 293.565 96.020 ;
        RECT 4.300 90.420 293.565 91.580 ;
        RECT 3.500 85.980 293.565 90.420 ;
        RECT 4.300 84.820 293.565 85.980 ;
        RECT 3.500 80.380 293.565 84.820 ;
        RECT 4.300 79.220 293.565 80.380 ;
        RECT 3.500 74.780 293.565 79.220 ;
        RECT 4.300 73.620 293.565 74.780 ;
        RECT 3.500 69.180 293.565 73.620 ;
        RECT 4.300 68.020 293.565 69.180 ;
        RECT 3.500 63.580 293.565 68.020 ;
        RECT 4.300 62.420 293.565 63.580 ;
        RECT 3.500 57.980 293.565 62.420 ;
        RECT 4.300 56.820 293.565 57.980 ;
        RECT 3.500 52.380 293.565 56.820 ;
        RECT 4.300 51.220 293.565 52.380 ;
        RECT 3.500 46.780 293.565 51.220 ;
        RECT 4.300 45.620 293.565 46.780 ;
        RECT 3.500 41.180 293.565 45.620 ;
        RECT 4.300 40.020 293.565 41.180 ;
        RECT 3.500 35.580 293.565 40.020 ;
        RECT 4.300 34.420 293.565 35.580 ;
        RECT 3.500 29.980 293.565 34.420 ;
        RECT 4.300 28.820 293.565 29.980 ;
        RECT 3.500 24.380 293.565 28.820 ;
        RECT 4.300 23.220 293.565 24.380 ;
        RECT 3.500 18.780 293.565 23.220 ;
        RECT 4.300 17.620 293.565 18.780 ;
        RECT 3.500 13.180 293.565 17.620 ;
        RECT 4.300 12.020 293.565 13.180 ;
        RECT 3.500 10.780 293.565 12.020 ;
      LAYER Metal4 ;
        RECT 10.220 21.370 41.385 172.950 ;
        RECT 43.585 21.370 77.150 172.950 ;
        RECT 79.350 21.370 112.920 172.950 ;
        RECT 115.120 21.370 148.685 172.950 ;
        RECT 150.885 21.370 184.455 172.950 ;
        RECT 186.655 21.370 220.220 172.950 ;
        RECT 222.420 21.370 255.990 172.950 ;
        RECT 258.190 21.370 284.900 172.950 ;
  END
END interp_tri
END LIBRARY

