// This is the unpowered netlist.
module interp_tri (clk,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_adr_i,
    wbs_dat_i,
    wbs_sel_i,
    x_end,
    x_start,
    y);
 input clk;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [3:2] wbs_adr_i;
 input [31:0] wbs_dat_i;
 input [3:0] wbs_sel_i;
 output [7:0] x_end;
 output [7:0] x_start;
 input [7:0] y;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire \a[0][0] ;
 wire \a[0][1] ;
 wire \a[0][2] ;
 wire \a[0][3] ;
 wire \a[0][4] ;
 wire \a[0][5] ;
 wire \a[0][6] ;
 wire \a[0][7] ;
 wire \a[1][0] ;
 wire \a[1][1] ;
 wire \a[1][2] ;
 wire \a[1][3] ;
 wire \a[1][4] ;
 wire \a[1][5] ;
 wire \a[1][6] ;
 wire \a[1][7] ;
 wire \b[0][0] ;
 wire \b[0][1] ;
 wire \b[0][2] ;
 wire \b[0][3] ;
 wire \b[0][4] ;
 wire \b[0][5] ;
 wire \b[0][6] ;
 wire \b[0][7] ;
 wire \b[1][0] ;
 wire \b[1][1] ;
 wire \b[1][2] ;
 wire \b[1][3] ;
 wire \b[1][4] ;
 wire \b[1][5] ;
 wire \b[1][6] ;
 wire \b[1][7] ;
 wire bflip;
 wire \c[0][0] ;
 wire \c[0][1] ;
 wire \c[0][2] ;
 wire \c[0][3] ;
 wire \c[0][4] ;
 wire \c[0][5] ;
 wire \c[0][6] ;
 wire \c[0][7] ;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \delta_t[0] ;
 wire \delta_t[1] ;
 wire \delta_t[2] ;
 wire \delta_t[3] ;
 wire \delta_t[4] ;
 wire \delta_t[5] ;
 wire \delta_t[6] ;
 wire \delta_t[7] ;
 wire \delta_t[8] ;
 wire \delta_t[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \t_reg[0] ;
 wire \t_reg[1] ;
 wire \t_reg[2] ;
 wire \t_reg[3] ;
 wire \t_reg[4] ;
 wire \t_reg[5] ;
 wire \t_reg[6] ;
 wire \t_reg[7] ;
 wire \t_reg[8] ;
 wire \t_reg[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__I (.I(\a[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1391__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1391__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1395__I (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__A3 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__I (.I(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__B2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__I (.I(\a[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__A1 (.I(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A2 (.I(\a[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__I (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__I (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__I (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A2 (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A2 (.I(\a[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(\a[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A1 (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A1 (.I(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A1 (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__A2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A3 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A1 (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A1 (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__I (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__B2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A1 (.I(\a[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__I (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(\b[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__I (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__I (.I(\a[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__I (.I(\a[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(\b[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A1 (.I(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__B (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(\a[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I (.I(\b[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__I (.I(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A3 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(\a[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A3 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I (.I(\c[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I (.I(\c[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__I (.I(\c[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A3 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__I (.I(\c[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__I (.I(\c[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A1 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__B2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__I (.I(\c[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(\c[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(\c[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__I (.I(\c[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A1 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(\c[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(\c[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__I (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A2 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(\c[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(\c[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(\c[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A1 (.I(\c[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A2 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A2 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(\c[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(\c[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A1 (.I(\c[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A1 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__I (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__I (.I(\c[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__I (.I(\c[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__B (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A3 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__I (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__B (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A1 (.I(\c[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A1 (.I(\c[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A3 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A4 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__C (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__C (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__C (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__C (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__C (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__C (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__C (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__C (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__C (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__C (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A3 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__C (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__I (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__B (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__B (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__B (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A1 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__B (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(wbs_sel_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(wbs_sel_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(wbs_sel_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(y[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(y[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(y[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(y[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(y[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(y[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(y[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(y[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(wbs_adr_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(wbs_adr_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer2_I (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1357_ (.A1(net27),
    .A2(net5),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1358_ (.I(_0551_),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1359_ (.I(\a[0][0] ),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1360_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1361_ (.I(\a[0][1] ),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1362_ (.I(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1363_ (.I(\a[0][0] ),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1364_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1365_ (.I0(\a[1][2] ),
    .I1(\b[1][2] ),
    .S(bflip),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1366_ (.A1(net31),
    .A2(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1367_ (.I0(\a[1][1] ),
    .I1(\b[1][1] ),
    .S(bflip),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1368_ (.A1(net30),
    .A2(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1369_ (.I(bflip),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1370_ (.I0(\a[1][6] ),
    .I1(\b[1][6] ),
    .S(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1371_ (.A1(_0563_),
    .A2(net35),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1372_ (.I0(\a[1][5] ),
    .I1(\b[1][5] ),
    .S(_0562_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1373_ (.A1(net34),
    .A2(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1374_ (.A1(_0559_),
    .A2(_0561_),
    .A3(_0564_),
    .A4(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1375_ (.I(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1376_ (.I0(\a[1][4] ),
    .I1(\b[1][4] ),
    .S(_0562_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1377_ (.A1(net33),
    .A2(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1378_ (.I0(\a[1][7] ),
    .I1(\b[1][7] ),
    .S(_0562_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1379_ (.A1(net36),
    .A2(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1380_ (.I(bflip),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1381_ (.I0(\a[1][0] ),
    .I1(\b[1][0] ),
    .S(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1382_ (.A1(_0574_),
    .A2(net29),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1383_ (.I0(\a[1][3] ),
    .I1(\b[1][3] ),
    .S(_0573_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1384_ (.A1(_0576_),
    .A2(net32),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1385_ (.A1(_0570_),
    .A2(_0572_),
    .A3(_0575_),
    .A4(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1386_ (.I(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1387_ (.I(\t_reg[5] ),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1388_ (.A1(_0568_),
    .A2(_0579_),
    .B(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1389_ (.A1(_0581_),
    .A2(\delta_t[6] ),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1390_ (.I(\delta_t[4] ),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1391_ (.A1(_0567_),
    .A2(_0578_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1392_ (.A1(_0584_),
    .A2(\t_reg[3] ),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1393_ (.I(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1394_ (.A1(_0586_),
    .A2(_0583_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1395_ (.I(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1396_ (.I(\delta_t[2] ),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _1397_ (.A1(_0559_),
    .A2(_0561_),
    .A3(_0564_),
    .A4(_0566_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _1398_ (.A1(_0570_),
    .A2(_0572_),
    .A3(_0575_),
    .A4(_0577_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1399_ (.A1(_0590_),
    .A2(_0591_),
    .B(\t_reg[1] ),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1400_ (.A1(_0590_),
    .A2(_0591_),
    .B(\delta_t[1] ),
    .C(\t_reg[0] ),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1401_ (.A1(_0589_),
    .A2(_0592_),
    .B(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1402_ (.A1(_0590_),
    .A2(_0591_),
    .B(\t_reg[2] ),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1403_ (.I(\delta_t[3] ),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1404_ (.A1(_0589_),
    .A2(_0592_),
    .B1(_0595_),
    .B2(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1405_ (.A1(_0596_),
    .A2(_0595_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1406_ (.A1(\delta_t[4] ),
    .A2(_0585_),
    .B1(_0594_),
    .B2(_0597_),
    .C(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1407_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1408_ (.I(\t_reg[4] ),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1409_ (.A1(_0568_),
    .A2(_0579_),
    .B(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1410_ (.A1(\delta_t[5] ),
    .A2(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1411_ (.I(\delta_t[5] ),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1412_ (.I(_0602_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1413_ (.A1(_0604_),
    .A2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1414_ (.A1(_0588_),
    .A2(_0600_),
    .A3(_0603_),
    .B(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1415_ (.A1(net94),
    .A2(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1416_ (.I(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1417_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1418_ (.A1(_0588_),
    .A2(_0600_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1419_ (.A1(\delta_t[5] ),
    .A2(_0602_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1420_ (.A1(_0611_),
    .A2(net80),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1421_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1422_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1423_ (.A1(_0555_),
    .A2(_0557_),
    .A3(_0610_),
    .A4(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1424_ (.I(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1425_ (.I(\a[0][2] ),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1426_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1427_ (.A1(_0619_),
    .A2(_0614_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1428_ (.I(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1429_ (.I(\delta_t[7] ),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1430_ (.I(\t_reg[6] ),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1431_ (.A1(_0568_),
    .A2(_0579_),
    .B(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1432_ (.A1(_0622_),
    .A2(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1433_ (.A1(_0582_),
    .A2(_0612_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1434_ (.A1(\delta_t[6] ),
    .A2(_0581_),
    .B1(_0602_),
    .B2(\delta_t[5] ),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1435_ (.I(_0581_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1436_ (.A1(\delta_t[6] ),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _1437_ (.A1(net77),
    .A2(net83),
    .A3(_0626_),
    .B1(_0627_),
    .B2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1438_ (.A1(_0625_),
    .A2(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1439_ (.I(net78),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1440_ (.I(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1441_ (.A1(_0557_),
    .A2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1442_ (.A1(_0555_),
    .A2(_0610_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1443_ (.A1(_0621_),
    .A2(_0634_),
    .A3(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1444_ (.A1(_0617_),
    .A2(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1445_ (.I(\b[0][2] ),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1446_ (.I(_0615_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1447_ (.A1(_0638_),
    .A2(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1448_ (.I(\b[0][1] ),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1449_ (.I(_0610_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1450_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1451_ (.A1(_0641_),
    .A2(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1452_ (.I(\b[0][0] ),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1453_ (.I(_0633_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1454_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1455_ (.A1(_0645_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1456_ (.A1(_0640_),
    .A2(_0644_),
    .A3(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1457_ (.I(_0641_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1458_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1459_ (.I(_0642_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1460_ (.I(_0652_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1461_ (.I(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1462_ (.I(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1463_ (.I(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1464_ (.I(_0639_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1465_ (.I(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1466_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1467_ (.I(_0645_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1468_ (.A1(_0651_),
    .A2(_0656_),
    .B(_0659_),
    .C(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1469_ (.A1(_0649_),
    .A2(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1470_ (.A1(_0637_),
    .A2(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1471_ (.I(_0659_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1472_ (.A1(_0660_),
    .A2(_0654_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1473_ (.A1(_0651_),
    .A2(_0664_),
    .B(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1474_ (.A1(_0660_),
    .A2(_0664_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1475_ (.A1(_0651_),
    .A2(_0656_),
    .B(_0666_),
    .C(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1476_ (.A1(_0649_),
    .A2(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1477_ (.A1(_0617_),
    .A2(_0636_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1478_ (.I(\a[0][3] ),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1479_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1480_ (.I(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1481_ (.A1(_0673_),
    .A2(_0615_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1482_ (.A1(_0634_),
    .A2(_0635_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1483_ (.A1(_0634_),
    .A2(_0635_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1484_ (.A1(_0621_),
    .A2(_0675_),
    .B(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1485_ (.A1(_0618_),
    .A2(_0608_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1486_ (.I(\delta_t[8] ),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1487_ (.I(\t_reg[7] ),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1488_ (.A1(_0568_),
    .A2(_0579_),
    .B(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1489_ (.A1(_0679_),
    .A2(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1490_ (.I(_0624_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1491_ (.A1(_0622_),
    .A2(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1492_ (.A1(_0625_),
    .A2(_0630_),
    .B(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1493_ (.A1(_0682_),
    .A2(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1494_ (.I(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1495_ (.A1(_0556_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1496_ (.A1(_0554_),
    .A2(_0632_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1497_ (.A1(_0678_),
    .A2(_0688_),
    .A3(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1498_ (.A1(_0674_),
    .A2(_0677_),
    .A3(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1499_ (.A1(_0670_),
    .A2(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1500_ (.I(_0657_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1501_ (.A1(_0650_),
    .A2(_0693_),
    .A3(_0649_),
    .A4(_0665_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1502_ (.I(\b[0][3] ),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1503_ (.I(_0615_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1504_ (.A1(_0695_),
    .A2(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1505_ (.A1(_0644_),
    .A2(_0648_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1506_ (.A1(_0644_),
    .A2(_0648_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1507_ (.A1(_0640_),
    .A2(_0698_),
    .B(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1508_ (.A1(_0638_),
    .A2(_0643_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1509_ (.I(_0687_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1510_ (.I(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1511_ (.A1(\b[0][0] ),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1512_ (.I(_0646_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1513_ (.A1(_0641_),
    .A2(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1514_ (.A1(_0701_),
    .A2(_0704_),
    .A3(_0706_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1515_ (.A1(_0697_),
    .A2(_0700_),
    .A3(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1516_ (.A1(_0694_),
    .A2(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1517_ (.A1(_0692_),
    .A2(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1518_ (.A1(_0663_),
    .A2(_0669_),
    .A3(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1519_ (.A1(_0637_),
    .A2(_0662_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1520_ (.I(_0555_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1521_ (.A1(_0557_),
    .A2(_0656_),
    .B1(_0664_),
    .B2(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1522_ (.A1(_0617_),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1523_ (.I(_0557_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1524_ (.I(_0664_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1525_ (.A1(_0716_),
    .A2(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1526_ (.A1(_0667_),
    .A2(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1527_ (.A1(_0666_),
    .A2(_0667_),
    .B(_0668_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1528_ (.A1(_0715_),
    .A2(_0719_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1529_ (.A1(_0720_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1530_ (.A1(_0715_),
    .A2(_0719_),
    .B(_0722_),
    .C(_0663_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1531_ (.A1(_0711_),
    .A2(_0712_),
    .A3(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1532_ (.A1(_0663_),
    .A2(_0669_),
    .B(_0710_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1533_ (.A1(_0670_),
    .A2(_0691_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1534_ (.I(\a[0][4] ),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1535_ (.I(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1536_ (.A1(_0728_),
    .A2(_0672_),
    .A3(_0608_),
    .A4(_0613_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1537_ (.A1(_0672_),
    .A2(_0609_),
    .B1(_0613_),
    .B2(_0728_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1538_ (.A1(_0729_),
    .A2(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1539_ (.I(_0678_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1540_ (.A1(\delta_t[8] ),
    .A2(_0681_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1541_ (.A1(net88),
    .A2(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1542_ (.I(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1543_ (.A1(_0553_),
    .A2(_0735_),
    .B(_0689_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1544_ (.I(_0552_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1545_ (.A1(_0737_),
    .A2(_0735_),
    .A3(_0689_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1546_ (.A1(_0732_),
    .A2(_0736_),
    .B(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1547_ (.A1(\a[0][2] ),
    .A2(_0631_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1548_ (.A1(_0686_),
    .A2(\a[0][1] ),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1549_ (.A1(net98),
    .A2(_0612_),
    .A3(_0625_),
    .A4(_0733_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1550_ (.A1(_0588_),
    .A2(_0600_),
    .A3(_0742_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1551_ (.I(\delta_t[8] ),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1552_ (.I(_0681_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1553_ (.A1(_0744_),
    .A2(_0745_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1554_ (.I(\delta_t[7] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1555_ (.A1(_0747_),
    .A2(_0624_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1556_ (.A1(_0629_),
    .A2(_0748_),
    .A3(_0627_),
    .A4(_0682_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1557_ (.A1(_0744_),
    .A2(_0681_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1558_ (.A1(_0684_),
    .A2(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1559_ (.A1(_0746_),
    .A2(_0749_),
    .A3(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1560_ (.A1(_0743_),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1561_ (.I0(_0573_),
    .I1(\t_reg[8] ),
    .S(_0584_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1562_ (.A1(\delta_t[9] ),
    .A2(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1563_ (.I(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1564_ (.A1(_0753_),
    .A2(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1565_ (.A1(_0552_),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1566_ (.A1(_0740_),
    .A2(_0741_),
    .A3(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1567_ (.A1(_0731_),
    .A2(_0739_),
    .A3(net87),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1568_ (.A1(_0677_),
    .A2(_0690_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1569_ (.A1(_0677_),
    .A2(_0690_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1570_ (.A1(_0674_),
    .A2(_0761_),
    .B(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1571_ (.A1(_0726_),
    .A2(_0760_),
    .A3(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1572_ (.A1(_0700_),
    .A2(_0707_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1573_ (.A1(_0700_),
    .A2(_0707_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1574_ (.A1(_0697_),
    .A2(_0765_),
    .B(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1575_ (.A1(\b[0][3] ),
    .A2(_0652_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1576_ (.A1(\b[0][4] ),
    .A2(_0696_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1577_ (.A1(_0768_),
    .A2(_0769_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1578_ (.A1(_0704_),
    .A2(_0706_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1579_ (.A1(_0704_),
    .A2(_0706_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1580_ (.A1(_0701_),
    .A2(_0771_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1581_ (.A1(\b[0][2] ),
    .A2(_0646_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1582_ (.A1(_0753_),
    .A2(_0755_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1583_ (.I(_0775_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1584_ (.I(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1585_ (.A1(\b[0][0] ),
    .A2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1586_ (.A1(\b[0][1] ),
    .A2(_0702_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1587_ (.A1(_0778_),
    .A2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1588_ (.A1(_0774_),
    .A2(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1589_ (.A1(_0773_),
    .A2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1590_ (.A1(_0770_),
    .A2(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1591_ (.A1(_0764_),
    .A2(_0767_),
    .A3(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1592_ (.A1(_0694_),
    .A2(_0708_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1593_ (.A1(_0692_),
    .A2(_0709_),
    .B(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1594_ (.A1(_0784_),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1595_ (.A1(_0725_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1596_ (.A1(_0724_),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1597_ (.A1(_0553_),
    .A2(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1598_ (.A1(_0784_),
    .A2(_0786_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1599_ (.A1(_0725_),
    .A2(_0787_),
    .B1(_0788_),
    .B2(_0724_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1600_ (.I(\b[0][4] ),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1601_ (.I(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1602_ (.A1(_0794_),
    .A2(_0659_),
    .A3(_0768_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1603_ (.A1(_0760_),
    .A2(_0763_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1604_ (.A1(_0760_),
    .A2(_0763_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1605_ (.A1(_0726_),
    .A2(_0796_),
    .B(net84),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1606_ (.I(_0731_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1607_ (.A1(_0759_),
    .A2(_0739_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1608_ (.A1(_0739_),
    .A2(_0759_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1609_ (.A1(_0799_),
    .A2(_0800_),
    .B(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(_0613_),
    .A2(\a[0][5] ),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1611_ (.A1(_0608_),
    .A2(\a[0][4] ),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1612_ (.A1(_0671_),
    .A2(net79),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1613_ (.A1(_0803_),
    .A2(_0804_),
    .A3(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1614_ (.I(\a[0][1] ),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1615_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1616_ (.A1(_0808_),
    .A2(_0734_),
    .B1(_0757_),
    .B2(_0737_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1617_ (.A1(_0807_),
    .A2(_0737_),
    .A3(_0734_),
    .A4(_0757_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1618_ (.A1(_0740_),
    .A2(_0809_),
    .B(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1619_ (.A1(_0618_),
    .A2(_0686_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1620_ (.A1(_0554_),
    .A2(_0775_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1621_ (.I(_0584_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1622_ (.A1(\delta_t[9] ),
    .A2(_0754_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1623_ (.A1(_0588_),
    .A2(_0600_),
    .A3(_0742_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1624_ (.A1(_0746_),
    .A2(_0749_),
    .A3(_0751_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1625_ (.A1(_0816_),
    .A2(_0817_),
    .B(_0755_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1626_ (.A1(\t_reg[9] ),
    .A2(_0814_),
    .B1(_0815_),
    .B2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1627_ (.I(_0815_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1628_ (.A1(_0743_),
    .A2(_0752_),
    .B(_0756_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1629_ (.A1(\t_reg[9] ),
    .A2(_0584_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1630_ (.A1(_0820_),
    .A2(_0821_),
    .A3(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1631_ (.A1(_0819_),
    .A2(_0823_),
    .B(\a[0][0] ),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1632_ (.A1(_0812_),
    .A2(_0813_),
    .A3(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1633_ (.A1(_0806_),
    .A2(_0811_),
    .A3(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1634_ (.A1(_0729_),
    .A2(_0802_),
    .A3(net97),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1635_ (.I(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1636_ (.A1(_0795_),
    .A2(_0798_),
    .A3(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1637_ (.A1(_0770_),
    .A2(_0782_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1638_ (.A1(_0773_),
    .A2(_0781_),
    .B(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1639_ (.A1(_0778_),
    .A2(_0779_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1640_ (.A1(_0774_),
    .A2(_0780_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1641_ (.A1(_0832_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1642_ (.I(_0703_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1643_ (.A1(_0638_),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1644_ (.A1(_0641_),
    .A2(_0776_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1645_ (.A1(_0820_),
    .A2(_0821_),
    .B(_0822_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1646_ (.A1(\t_reg[9] ),
    .A2(_0814_),
    .A3(_0815_),
    .A4(_0818_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1647_ (.A1(_0838_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1648_ (.I(_0840_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1649_ (.A1(\b[0][0] ),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1650_ (.A1(_0837_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1651_ (.A1(_0836_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1652_ (.A1(_0834_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1653_ (.A1(\b[0][5] ),
    .A2(_0696_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1654_ (.A1(\b[0][4] ),
    .A2(_0642_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1655_ (.A1(\b[0][3] ),
    .A2(_0705_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1656_ (.A1(_0847_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1657_ (.A1(_0846_),
    .A2(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1658_ (.A1(_0845_),
    .A2(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1659_ (.A1(_0831_),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1660_ (.A1(_0829_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1661_ (.A1(_0767_),
    .A2(_0783_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1662_ (.A1(_0767_),
    .A2(_0783_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1663_ (.A1(_0764_),
    .A2(_0854_),
    .B(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1664_ (.A1(_0853_),
    .A2(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1665_ (.A1(_0791_),
    .A2(_0792_),
    .A3(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1666_ (.A1(_0713_),
    .A2(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1667_ (.A1(_0790_),
    .A2(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1668_ (.I(_0860_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1669_ (.A1(_0713_),
    .A2(_0858_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1670_ (.A1(_0790_),
    .A2(_0859_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1671_ (.A1(_0861_),
    .A2(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1672_ (.I(_0619_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1673_ (.I(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1674_ (.A1(_0853_),
    .A2(_0856_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1675_ (.A1(_0791_),
    .A2(_0857_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1676_ (.A1(_0791_),
    .A2(_0857_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1677_ (.A1(_0792_),
    .A2(_0867_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1678_ (.A1(_0798_),
    .A2(_0828_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1679_ (.A1(_0794_),
    .A2(_0717_),
    .A3(_0768_),
    .A4(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1680_ (.A1(_0831_),
    .A2(_0851_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1681_ (.A1(_0829_),
    .A2(_0852_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1682_ (.A1(_0872_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1683_ (.A1(_0847_),
    .A2(_0848_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1684_ (.A1(_0846_),
    .A2(_0849_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1685_ (.A1(_0875_),
    .A2(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1686_ (.A1(\b[0][6] ),
    .A2(_0693_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1687_ (.A1(_0726_),
    .A2(_0796_),
    .A3(_0828_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1688_ (.A1(_0797_),
    .A2(_0827_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1689_ (.A1(net86),
    .A2(_0826_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1690_ (.A1(net96),
    .A2(net95),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1691_ (.A1(_0729_),
    .A2(_0881_),
    .B(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1692_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1693_ (.A1(_0804_),
    .A2(_0805_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1694_ (.A1(_0804_),
    .A2(_0805_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1695_ (.A1(_0803_),
    .A2(_0885_),
    .B(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1696_ (.I(\a[0][6] ),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1697_ (.A1(_0888_),
    .A2(_0614_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1698_ (.A1(_0887_),
    .A2(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1699_ (.A1(_0811_),
    .A2(_0825_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1700_ (.A1(net99),
    .A2(_0825_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1701_ (.A1(net85),
    .A2(_0891_),
    .B(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1702_ (.A1(\a[0][5] ),
    .A2(_0609_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1703_ (.A1(_0727_),
    .A2(_0671_),
    .A3(_0632_),
    .A4(_0687_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1704_ (.I(\a[0][3] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1705_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1706_ (.A1(_0727_),
    .A2(_0632_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1707_ (.A1(_0897_),
    .A2(_0734_),
    .B(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1708_ (.A1(_0895_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1709_ (.A1(_0894_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1710_ (.A1(_0813_),
    .A2(_0824_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1711_ (.A1(_0813_),
    .A2(_0824_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1712_ (.A1(_0812_),
    .A2(_0902_),
    .B(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1713_ (.A1(_0808_),
    .A2(_0737_),
    .B1(_0838_),
    .B2(_0839_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1714_ (.I(_0819_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1715_ (.I(_0823_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1716_ (.A1(_0906_),
    .A2(_0907_),
    .B(_0555_),
    .C(_0556_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1717_ (.A1(_0905_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1718_ (.A1(_0619_),
    .A2(_0776_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1719_ (.A1(_0909_),
    .A2(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1720_ (.A1(_0901_),
    .A2(_0904_),
    .A3(_0911_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1721_ (.A1(_0890_),
    .A2(_0893_),
    .A3(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1722_ (.I(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1723_ (.A1(net90),
    .A2(_0884_),
    .A3(_0914_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1724_ (.A1(_0878_),
    .A2(_0879_),
    .A3(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1725_ (.A1(_0834_),
    .A2(_0844_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1726_ (.A1(_0845_),
    .A2(_0850_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1727_ (.A1(_0917_),
    .A2(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1728_ (.A1(_0836_),
    .A2(_0843_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1729_ (.A1(_0837_),
    .A2(_0842_),
    .B(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1730_ (.I(_0841_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1731_ (.I(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1732_ (.A1(_0650_),
    .A2(_0645_),
    .B(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1733_ (.A1(_0650_),
    .A2(_0645_),
    .A3(_0922_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1734_ (.A1(_0924_),
    .A2(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1735_ (.I(_0638_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1736_ (.I(_0777_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1737_ (.A1(_0927_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1738_ (.A1(_0926_),
    .A2(_0929_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1739_ (.A1(\b[0][5] ),
    .A2(_0653_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1740_ (.I(_0647_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1741_ (.A1(\b[0][4] ),
    .A2(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1742_ (.I(_0835_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1743_ (.A1(_0695_),
    .A2(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1744_ (.A1(_0933_),
    .A2(_0935_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1745_ (.A1(_0933_),
    .A2(_0935_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1746_ (.A1(_0936_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1747_ (.A1(_0931_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1748_ (.A1(_0921_),
    .A2(_0930_),
    .A3(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1749_ (.A1(_0919_),
    .A2(_0940_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1750_ (.A1(_0877_),
    .A2(_0916_),
    .A3(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1751_ (.A1(_0871_),
    .A2(_0874_),
    .A3(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1752_ (.A1(_0866_),
    .A2(_0869_),
    .A3(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1753_ (.A1(_0865_),
    .A2(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1754_ (.A1(_0863_),
    .A2(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1755_ (.I(_0946_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1756_ (.A1(_0865_),
    .A2(_0944_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1757_ (.A1(_0863_),
    .A2(_0945_),
    .B(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1758_ (.A1(_0866_),
    .A2(_0943_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1759_ (.A1(_0866_),
    .A2(_0943_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1760_ (.A1(_0869_),
    .A2(_0949_),
    .B(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1761_ (.A1(_0879_),
    .A2(_0915_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1762_ (.A1(_0878_),
    .A2(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1763_ (.A1(_0877_),
    .A2(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1764_ (.A1(_0874_),
    .A2(_0942_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1765_ (.A1(_0874_),
    .A2(_0942_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1766_ (.A1(_0871_),
    .A2(_0955_),
    .B(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1767_ (.A1(_0877_),
    .A2(_0916_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1768_ (.A1(_0919_),
    .A2(_0940_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1769_ (.A1(_0958_),
    .A2(_0941_),
    .B(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1770_ (.A1(_0921_),
    .A2(_0930_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1771_ (.A1(_0921_),
    .A2(_0930_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1772_ (.A1(_0961_),
    .A2(_0939_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1773_ (.A1(_0926_),
    .A2(_0929_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1774_ (.A1(_0927_),
    .A2(_0923_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1775_ (.A1(_0926_),
    .A2(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1776_ (.A1(_0927_),
    .A2(_0925_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1777_ (.A1(_0925_),
    .A2(_0964_),
    .A3(_0966_),
    .B(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1778_ (.I(_0932_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1779_ (.A1(\b[0][5] ),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1780_ (.A1(_0793_),
    .A2(_0934_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1781_ (.I(_0695_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1782_ (.I(_0928_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1783_ (.A1(_0972_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1784_ (.A1(_0970_),
    .A2(_0971_),
    .A3(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1785_ (.A1(_0968_),
    .A2(_0975_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1786_ (.A1(_0963_),
    .A2(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1787_ (.I(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1788_ (.A1(_0878_),
    .A2(_0952_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1789_ (.A1(_0931_),
    .A2(_0938_),
    .B(_0936_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1790_ (.A1(_0884_),
    .A2(_0914_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1791_ (.A1(_0884_),
    .A2(_0914_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1792_ (.A1(_0880_),
    .A2(_0883_),
    .A3(_0913_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _1793_ (.A1(net91),
    .A2(_0981_),
    .A3(_0982_),
    .B1(_0983_),
    .B2(_0879_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1794_ (.I(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1795_ (.I(_0888_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1796_ (.A1(_0986_),
    .A2(_0639_),
    .A3(_0887_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1797_ (.A1(_0893_),
    .A2(_0912_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1798_ (.A1(_0893_),
    .A2(_0912_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1799_ (.A1(_0890_),
    .A2(_0988_),
    .B(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1800_ (.A1(_0894_),
    .A2(_0900_),
    .B(_0895_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1801_ (.A1(\a[0][6] ),
    .A2(_0609_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1802_ (.A1(_0991_),
    .A2(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1803_ (.A1(\a[0][7] ),
    .A2(_0614_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1804_ (.A1(_0993_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1805_ (.A1(_0904_),
    .A2(_0911_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1806_ (.A1(_0904_),
    .A2(_0911_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1807_ (.A1(_0901_),
    .A2(_0996_),
    .B(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1808_ (.I(\a[0][5] ),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1809_ (.A1(_0999_),
    .A2(_0633_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1810_ (.A1(_0728_),
    .A2(_0702_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1811_ (.I(_0672_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1812_ (.A1(_1002_),
    .A2(_0775_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1813_ (.A1(_1000_),
    .A2(_1001_),
    .A3(_1003_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1814_ (.A1(_0906_),
    .A2(_0907_),
    .B(_0619_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1815_ (.A1(_0905_),
    .A2(_0908_),
    .A3(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1816_ (.A1(_0905_),
    .A2(_0908_),
    .B(_1005_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1817_ (.A1(_0554_),
    .A2(_0556_),
    .B1(_0906_),
    .B2(_0907_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1818_ (.A1(_1008_),
    .A2(_0910_),
    .B(_0908_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1819_ (.A1(_0838_),
    .A2(_0839_),
    .B(_0807_),
    .C(_0552_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1820_ (.A1(_0864_),
    .A2(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1821_ (.A1(_1006_),
    .A2(_1007_),
    .A3(_1009_),
    .B(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1822_ (.A1(_1004_),
    .A2(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1823_ (.A1(_0995_),
    .A2(_0998_),
    .A3(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1824_ (.A1(_0987_),
    .A2(_0990_),
    .A3(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1825_ (.A1(_1015_),
    .A2(_0981_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1826_ (.A1(\b[0][6] ),
    .A2(_0654_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1827_ (.A1(\b[0][7] ),
    .A2(_0658_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1828_ (.A1(_1017_),
    .A2(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1829_ (.A1(_0985_),
    .A2(_1016_),
    .A3(_1019_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1830_ (.A1(_0979_),
    .A2(_0980_),
    .A3(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1831_ (.A1(_0960_),
    .A2(_0978_),
    .A3(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1832_ (.A1(_0954_),
    .A2(_0957_),
    .A3(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1833_ (.A1(_0951_),
    .A2(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1834_ (.A1(_0897_),
    .A2(_1024_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1835_ (.A1(_0948_),
    .A2(_1025_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1836_ (.I(_1026_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1837_ (.A1(_0673_),
    .A2(_1024_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1838_ (.A1(_0948_),
    .A2(_1025_),
    .B(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1839_ (.I(_0728_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1840_ (.A1(_0954_),
    .A2(_1022_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1841_ (.A1(_0951_),
    .A2(_1023_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1842_ (.A1(_0957_),
    .A2(_1030_),
    .B(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1843_ (.A1(_0978_),
    .A2(_1021_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1844_ (.A1(_0954_),
    .A2(_1022_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1845_ (.A1(_0960_),
    .A2(_1033_),
    .B(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1846_ (.A1(_0980_),
    .A2(_1020_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1847_ (.A1(_0980_),
    .A2(_1020_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1848_ (.A1(_0979_),
    .A2(_1036_),
    .B(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1849_ (.A1(_0979_),
    .A2(_0980_),
    .A3(_1020_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1850_ (.A1(_0963_),
    .A2(_0976_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1851_ (.A1(_0978_),
    .A2(_1039_),
    .B(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1852_ (.I(_0967_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1853_ (.A1(_0968_),
    .A2(_0975_),
    .B(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1854_ (.A1(_0924_),
    .A2(_0965_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1855_ (.A1(_0967_),
    .A2(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1856_ (.I(\b[0][5] ),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1857_ (.I(_0934_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1858_ (.A1(_1046_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1859_ (.A1(_0793_),
    .A2(_0928_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1860_ (.A1(_0695_),
    .A2(_0923_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1861_ (.A1(_1049_),
    .A2(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1862_ (.A1(_1048_),
    .A2(_1051_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1863_ (.A1(_1045_),
    .A2(_1052_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1864_ (.A1(_1043_),
    .A2(_1053_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1865_ (.I(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1866_ (.A1(_0985_),
    .A2(_1016_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1867_ (.I(_1019_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1868_ (.A1(_1017_),
    .A2(_1018_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1869_ (.A1(_1056_),
    .A2(_1057_),
    .B(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1870_ (.A1(_0971_),
    .A2(_0974_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1871_ (.A1(_0971_),
    .A2(_0974_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1872_ (.A1(_0970_),
    .A2(_1060_),
    .B(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1873_ (.A1(_0884_),
    .A2(_0914_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1874_ (.A1(_1063_),
    .A2(_1015_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1875_ (.A1(_1063_),
    .A2(_1015_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1876_ (.A1(_0984_),
    .A2(_1064_),
    .B(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1877_ (.A1(_0990_),
    .A2(_1014_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1878_ (.A1(_0990_),
    .A2(_1014_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1879_ (.A1(_0987_),
    .A2(_1067_),
    .B(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1880_ (.A1(_0986_),
    .A2(_0652_),
    .A3(_0991_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1881_ (.I(\a[0][7] ),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1882_ (.A1(_1071_),
    .A2(_0696_),
    .A3(_0993_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1883_ (.A1(_1070_),
    .A2(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1884_ (.A1(_0998_),
    .A2(_1013_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1885_ (.A1(_0998_),
    .A2(_1013_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1886_ (.A1(_0995_),
    .A2(_1074_),
    .B(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1887_ (.A1(_1004_),
    .A2(_1012_),
    .B(_1011_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1888_ (.A1(_0618_),
    .A2(_1010_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1889_ (.A1(_1008_),
    .A2(_1005_),
    .B(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1890_ (.I(_1079_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1891_ (.A1(_0999_),
    .A2(_0687_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _1892_ (.I(\a[0][4] ),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1893_ (.A1(_1082_),
    .A2(_0757_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1894_ (.I(_0840_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1895_ (.A1(_1002_),
    .A2(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1896_ (.A1(_1081_),
    .A2(_1083_),
    .A3(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1897_ (.A1(_1080_),
    .A2(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1898_ (.A1(_1077_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1899_ (.A1(_1001_),
    .A2(_1003_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1900_ (.A1(_1001_),
    .A2(_1003_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1901_ (.A1(_1000_),
    .A2(_1089_),
    .B(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1902_ (.A1(_0986_),
    .A2(_0633_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1903_ (.A1(_1091_),
    .A2(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1904_ (.A1(_1071_),
    .A2(_0610_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1905_ (.A1(_1093_),
    .A2(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1906_ (.A1(_1088_),
    .A2(_1095_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1907_ (.A1(_1073_),
    .A2(_1076_),
    .A3(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1908_ (.A1(_1069_),
    .A2(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(\b[0][7] ),
    .A2(_0655_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1910_ (.I(_0969_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1911_ (.A1(\b[0][6] ),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1912_ (.A1(_1099_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1913_ (.A1(_1066_),
    .A2(_1098_),
    .A3(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1914_ (.A1(_1059_),
    .A2(_1062_),
    .A3(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1915_ (.A1(_1041_),
    .A2(_1055_),
    .A3(_1104_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1916_ (.A1(_1038_),
    .A2(_1105_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1917_ (.A1(_1035_),
    .A2(_1106_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1918_ (.A1(_1029_),
    .A2(_1032_),
    .A3(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1919_ (.A1(_1028_),
    .A2(_1108_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1920_ (.I(_1109_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1921_ (.A1(_1032_),
    .A2(_1107_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1922_ (.A1(_1029_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1923_ (.A1(_1028_),
    .A2(_1108_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1924_ (.I(_0999_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1925_ (.A1(_1035_),
    .A2(_1106_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1926_ (.A1(_1032_),
    .A2(_1107_),
    .B(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1927_ (.A1(_1055_),
    .A2(_1104_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1928_ (.A1(_1041_),
    .A2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1929_ (.A1(_1038_),
    .A2(_1105_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1930_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1931_ (.I(_1062_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1932_ (.A1(_1120_),
    .A2(_1103_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1933_ (.A1(_1120_),
    .A2(_1103_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1934_ (.A1(_1059_),
    .A2(_1121_),
    .A3(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1935_ (.A1(_1121_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1936_ (.A1(_1043_),
    .A2(_1053_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1937_ (.A1(_1055_),
    .A2(_1104_),
    .B(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1938_ (.I(_1045_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1939_ (.A1(_1127_),
    .A2(_1052_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1940_ (.A1(_1042_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1941_ (.I(_0923_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1942_ (.A1(_0793_),
    .A2(_0972_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1943_ (.I(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1944_ (.I(_1130_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1945_ (.A1(_0794_),
    .A2(_0972_),
    .A3(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1946_ (.A1(_1132_),
    .A2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1947_ (.I(_0973_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1948_ (.I(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1949_ (.A1(_1046_),
    .A2(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1950_ (.A1(_1135_),
    .A2(_1138_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1951_ (.A1(_1127_),
    .A2(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1952_ (.A1(_1129_),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1953_ (.A1(_1066_),
    .A2(_1098_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1954_ (.A1(_1099_),
    .A2(_1101_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1955_ (.A1(_1142_),
    .A2(_1102_),
    .B(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1956_ (.A1(_1049_),
    .A2(_1050_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1957_ (.A1(_1048_),
    .A2(_1051_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1958_ (.A1(_1145_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1959_ (.A1(_1069_),
    .A2(_1097_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1960_ (.A1(_1069_),
    .A2(_1097_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1961_ (.A1(_1066_),
    .A2(_1148_),
    .B(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1962_ (.I(_1096_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1963_ (.A1(_1076_),
    .A2(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1964_ (.A1(_1076_),
    .A2(_1151_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1965_ (.A1(_1073_),
    .A2(_1152_),
    .B(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1966_ (.I(_0986_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1967_ (.A1(_1155_),
    .A2(_0932_),
    .A3(_1091_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1968_ (.A1(_1093_),
    .A2(_1094_),
    .B(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1969_ (.A1(_1077_),
    .A2(_1087_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1970_ (.A1(_1088_),
    .A2(_1095_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1971_ (.A1(_1158_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1972_ (.A1(_1080_),
    .A2(_1086_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1973_ (.A1(_1011_),
    .A2(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1974_ (.A1(_0727_),
    .A2(_0671_),
    .B(_0840_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1975_ (.A1(_0838_),
    .A2(_0839_),
    .B(_1082_),
    .C(_0896_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1976_ (.A1(_1163_),
    .A2(_1164_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1977_ (.A1(_0999_),
    .A2(_0775_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1978_ (.A1(_1165_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1979_ (.A1(_1079_),
    .A2(_1167_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1980_ (.A1(_1162_),
    .A2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1981_ (.A1(_1002_),
    .A2(_1084_),
    .B(_1083_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1982_ (.A1(_1002_),
    .A2(_1084_),
    .A3(_1083_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1983_ (.A1(_1081_),
    .A2(_1170_),
    .B(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1984_ (.A1(_0888_),
    .A2(_0702_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1985_ (.A1(_1172_),
    .A2(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1986_ (.A1(\a[0][7] ),
    .A2(_0646_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1987_ (.A1(_1174_),
    .A2(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1988_ (.A1(_1169_),
    .A2(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1989_ (.A1(_1160_),
    .A2(_1177_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1990_ (.A1(_1157_),
    .A2(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1991_ (.A1(_1154_),
    .A2(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1992_ (.I(\b[0][7] ),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1993_ (.A1(_1181_),
    .A2(_1100_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1994_ (.I(\b[0][6] ),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1995_ (.I(_1047_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1996_ (.A1(_1183_),
    .A2(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1997_ (.A1(_1182_),
    .A2(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1998_ (.A1(_1150_),
    .A2(_1180_),
    .A3(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1999_ (.A1(_1144_),
    .A2(_1147_),
    .A3(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2000_ (.A1(_1126_),
    .A2(_1141_),
    .A3(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2001_ (.A1(_1124_),
    .A2(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2002_ (.A1(_1119_),
    .A2(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2003_ (.A1(_1113_),
    .A2(_1115_),
    .A3(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2004_ (.A1(_1111_),
    .A2(_1112_),
    .B(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2005_ (.A1(_1111_),
    .A2(_1112_),
    .A3(_1192_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2006_ (.A1(_1193_),
    .A2(_1194_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2007_ (.A1(_1115_),
    .A2(_1191_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2008_ (.A1(_1113_),
    .A2(_1195_),
    .B(_1193_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2009_ (.I(_1155_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2010_ (.A1(_1119_),
    .A2(_1190_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2011_ (.A1(_1119_),
    .A2(_1190_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2012_ (.A1(_1115_),
    .A2(_1198_),
    .B(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2013_ (.A1(_1141_),
    .A2(_1188_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2014_ (.A1(_1126_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2015_ (.A1(_1124_),
    .A2(_1189_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2016_ (.A1(_1202_),
    .A2(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2017_ (.A1(_1150_),
    .A2(_1180_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2018_ (.A1(_1205_),
    .A2(_1186_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2019_ (.A1(_1147_),
    .A2(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2020_ (.A1(_1147_),
    .A2(_1187_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2021_ (.A1(_1144_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2022_ (.A1(_1207_),
    .A2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2023_ (.A1(_1129_),
    .A2(_1140_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2024_ (.A1(_1141_),
    .A2(_1188_),
    .B(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2025_ (.I(_1186_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2026_ (.A1(_1182_),
    .A2(_1185_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2027_ (.A1(_1205_),
    .A2(_1213_),
    .B(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2028_ (.A1(_1131_),
    .A2(_1138_),
    .B(_1134_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2029_ (.I(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2030_ (.A1(_1154_),
    .A2(_1179_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2031_ (.A1(_1154_),
    .A2(_1179_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2032_ (.A1(_1150_),
    .A2(_1218_),
    .B(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2033_ (.A1(_1160_),
    .A2(_1177_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2034_ (.A1(_1157_),
    .A2(_1178_),
    .B(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2035_ (.A1(_1155_),
    .A2(_0934_),
    .A3(_1172_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2036_ (.A1(_1174_),
    .A2(_1175_),
    .B(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2037_ (.A1(_1162_),
    .A2(_1168_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2038_ (.A1(_1169_),
    .A2(_1176_),
    .B(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2039_ (.A1(_1080_),
    .A2(_1167_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2040_ (.A1(_1011_),
    .A2(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2041_ (.A1(_1113_),
    .A2(_1084_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2042_ (.A1(_1165_),
    .A2(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2043_ (.A1(_1080_),
    .A2(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2044_ (.A1(_1228_),
    .A2(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2045_ (.A1(_1029_),
    .A2(_0673_),
    .A3(_0841_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2046_ (.A1(_1163_),
    .A2(_1166_),
    .B(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2047_ (.A1(_0888_),
    .A2(_0776_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2048_ (.A1(_1234_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2049_ (.A1(\a[0][7] ),
    .A2(_0703_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2050_ (.A1(_1236_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2051_ (.A1(_1232_),
    .A2(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2052_ (.A1(_1226_),
    .A2(_1239_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2053_ (.A1(_1224_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2054_ (.A1(_1222_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2055_ (.A1(_1181_),
    .A2(_1184_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2056_ (.I(_1136_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2057_ (.A1(_1183_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2058_ (.A1(_1243_),
    .A2(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2059_ (.A1(_1220_),
    .A2(_1242_),
    .A3(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2060_ (.A1(_1215_),
    .A2(_1217_),
    .A3(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2061_ (.A1(_1127_),
    .A2(_1139_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2062_ (.A1(_1042_),
    .A2(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2063_ (.A1(_1046_),
    .A2(_1133_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2064_ (.A1(_1135_),
    .A2(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2065_ (.A1(_1127_),
    .A2(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2066_ (.A1(_1250_),
    .A2(_1253_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2067_ (.A1(_1248_),
    .A2(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2068_ (.A1(_1210_),
    .A2(_1212_),
    .A3(_1255_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2069_ (.A1(_1204_),
    .A2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2070_ (.A1(_1200_),
    .A2(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2071_ (.A1(_1197_),
    .A2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2072_ (.A1(_1196_),
    .A2(_1259_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2073_ (.I(_1260_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2074_ (.I(_1071_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2075_ (.A1(_1202_),
    .A2(_1203_),
    .B(_1256_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2076_ (.A1(_1200_),
    .A2(_1257_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2077_ (.A1(_1261_),
    .A2(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2078_ (.A1(_1212_),
    .A2(_1255_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2079_ (.A1(_1210_),
    .A2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2080_ (.A1(_1212_),
    .A2(_1255_),
    .B(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2081_ (.A1(_1222_),
    .A2(_1241_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2082_ (.A1(_1220_),
    .A2(_1242_),
    .B(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2083_ (.A1(_1226_),
    .A2(_1239_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2084_ (.A1(_1224_),
    .A2(_1240_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2085_ (.A1(_1270_),
    .A2(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2086_ (.A1(_1261_),
    .A2(_1244_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2087_ (.A1(_1272_),
    .A2(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2088_ (.A1(_1163_),
    .A2(_1229_),
    .B(_1233_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2089_ (.A1(_1197_),
    .A2(_1133_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2090_ (.A1(_1155_),
    .A2(_1137_),
    .A3(_1234_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2091_ (.A1(_1071_),
    .A2(_1184_),
    .A3(_1236_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2092_ (.A1(_1277_),
    .A2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2093_ (.A1(_1276_),
    .A2(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2094_ (.A1(_1275_),
    .A2(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2095_ (.A1(_1228_),
    .A2(_1231_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2096_ (.A1(_1232_),
    .A2(_1238_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2097_ (.A1(_1282_),
    .A2(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2098_ (.I(_1133_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2099_ (.A1(_0864_),
    .A2(_1285_),
    .B(_0905_),
    .C(_1230_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2100_ (.A1(_1078_),
    .A2(_1230_),
    .B(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2101_ (.A1(_1281_),
    .A2(_1284_),
    .A3(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2102_ (.A1(_1269_),
    .A2(_1274_),
    .A3(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2103_ (.A1(_1220_),
    .A2(_1242_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2104_ (.A1(_1243_),
    .A2(_1245_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2105_ (.A1(_1243_),
    .A2(_1245_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2106_ (.A1(_1290_),
    .A2(_1291_),
    .B(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2107_ (.A1(_1250_),
    .A2(_1253_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2108_ (.A1(_1248_),
    .A2(_1254_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(_1294_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2110_ (.A1(_1183_),
    .A2(_1285_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2111_ (.A1(_1181_),
    .A2(_1244_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2112_ (.A1(_1131_),
    .A2(_1251_),
    .B(_1134_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2113_ (.A1(_1217_),
    .A2(_1247_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2114_ (.A1(_1215_),
    .A2(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2115_ (.A1(_1217_),
    .A2(_1247_),
    .B(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2116_ (.A1(_1298_),
    .A2(_1299_),
    .A3(_1302_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2117_ (.I0(_1044_),
    .I1(_1042_),
    .S(_1252_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2118_ (.A1(_1297_),
    .A2(_1303_),
    .A3(_1304_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2119_ (.A1(_1293_),
    .A2(_1296_),
    .A3(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2120_ (.A1(_1267_),
    .A2(_1289_),
    .A3(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2121_ (.A1(_1197_),
    .A2(_1258_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2122_ (.A1(_1196_),
    .A2(_1259_),
    .B(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2123_ (.A1(_1264_),
    .A2(_1307_),
    .A3(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2124_ (.I(_1310_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2125_ (.A1(_0553_),
    .A2(_0789_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2126_ (.I(_1311_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2127_ (.I(_0814_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2128_ (.A1(\delta_t[0] ),
    .A2(\t_reg[0] ),
    .A3(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2129_ (.I(\delta_t[1] ),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2130_ (.A1(_1314_),
    .A2(_0592_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2131_ (.A1(_1313_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2132_ (.I(_1316_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2133_ (.A1(\delta_t[1] ),
    .A2(\t_reg[1] ),
    .A3(_1312_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2134_ (.A1(\delta_t[0] ),
    .A2(\t_reg[0] ),
    .A3(_0814_),
    .A4(_1315_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2135_ (.A1(_1317_),
    .A2(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2136_ (.A1(\delta_t[2] ),
    .A2(_0595_),
    .A3(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2137_ (.I(_1320_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2138_ (.A1(_0589_),
    .A2(_0595_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2139_ (.A1(\delta_t[2] ),
    .A2(\t_reg[2] ),
    .A3(_1312_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2140_ (.A1(_1319_),
    .A2(_1321_),
    .B(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2141_ (.A1(\delta_t[3] ),
    .A2(_0586_),
    .A3(_1323_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2142_ (.I(_1324_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2143_ (.I(_0583_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2144_ (.A1(\delta_t[3] ),
    .A2(_0586_),
    .B(_1323_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2145_ (.I(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2146_ (.A1(\delta_t[3] ),
    .A2(_0586_),
    .B(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2147_ (.A1(_1325_),
    .A2(_0605_),
    .A3(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2148_ (.I(_1329_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2149_ (.I(_0604_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2150_ (.A1(_0583_),
    .A2(_0605_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2151_ (.A1(_1328_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2152_ (.A1(_0583_),
    .A2(_0605_),
    .B(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2153_ (.A1(_1330_),
    .A2(_0628_),
    .A3(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2154_ (.I(_1334_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2155_ (.I(\delta_t[6] ),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2156_ (.A1(_0604_),
    .A2(_0628_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2157_ (.A1(_1333_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2158_ (.A1(_0604_),
    .A2(_0628_),
    .B(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2159_ (.A1(_1335_),
    .A2(_0683_),
    .A3(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2160_ (.I(_1339_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2161_ (.A1(_1335_),
    .A2(_0683_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2162_ (.A1(_1338_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2163_ (.A1(_1335_),
    .A2(_0683_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2164_ (.A1(_0747_),
    .A2(_0745_),
    .A3(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2165_ (.I(_1343_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2166_ (.A1(_0744_),
    .A2(_0754_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2167_ (.A1(_0622_),
    .A2(_0745_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2168_ (.A1(_0622_),
    .A2(_0745_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2169_ (.A1(_1342_),
    .A2(_1345_),
    .B(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2170_ (.A1(_1344_),
    .A2(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2171_ (.I(_1348_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2172_ (.I(\delta_t[9] ),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2173_ (.A1(_0744_),
    .A2(_0754_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2174_ (.A1(_1344_),
    .A2(_1347_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2175_ (.A1(_1350_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2176_ (.A1(_1349_),
    .A2(_0822_),
    .A3(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2177_ (.I(_1353_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2178_ (.A1(\t_reg[0] ),
    .A2(_1312_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2179_ (.A1(\delta_t[0] ),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2180_ (.I(_1355_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2181_ (.I(\c[0][0] ),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2182_ (.A1(_1356_),
    .A2(_0969_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2183_ (.I(\c[0][1] ),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2184_ (.A1(_0078_),
    .A2(_0653_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2185_ (.I(\c[0][2] ),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2186_ (.A1(_0080_),
    .A2(_0657_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2187_ (.A1(_0079_),
    .A2(_0081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2188_ (.A1(_0077_),
    .A2(_0082_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2189_ (.I(_0078_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2190_ (.I(_1356_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2191_ (.A1(_0084_),
    .A2(_0085_),
    .A3(_0655_),
    .A4(_0659_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2192_ (.A1(_0083_),
    .A2(_0086_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2193_ (.A1(_0616_),
    .A2(_0636_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2194_ (.A1(_0083_),
    .A2(_0086_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2195_ (.A1(_0088_),
    .A2(_0089_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2196_ (.A1(_0087_),
    .A2(_0090_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2197_ (.A1(_0077_),
    .A2(_0082_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2198_ (.A1(_0079_),
    .A2(_0081_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2199_ (.I(\c[0][0] ),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2200_ (.A1(_0094_),
    .A2(_0735_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2201_ (.A1(_0078_),
    .A2(_0932_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2202_ (.I(\c[0][2] ),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2203_ (.A1(_0097_),
    .A2(_0643_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2204_ (.I(\c[0][3] ),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2205_ (.A1(_0099_),
    .A2(_0639_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2206_ (.A1(_0096_),
    .A2(_0098_),
    .A3(_0100_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2207_ (.A1(_0093_),
    .A2(_0095_),
    .A3(_0101_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2208_ (.A1(_0092_),
    .A2(_0102_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2209_ (.A1(_0692_),
    .A2(_0103_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2210_ (.A1(_0091_),
    .A2(_0104_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2211_ (.A1(_0088_),
    .A2(_0089_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2212_ (.A1(_0085_),
    .A2(_0656_),
    .B1(_0717_),
    .B2(_0084_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2213_ (.A1(_0715_),
    .A2(_0107_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2214_ (.A1(_0094_),
    .A2(_0716_),
    .A3(_0717_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2215_ (.I(_0086_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2216_ (.A1(_0110_),
    .A2(_0107_),
    .B(_0715_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2217_ (.A1(_0108_),
    .A2(_0109_),
    .B(_0111_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2218_ (.A1(_0090_),
    .A2(_0106_),
    .A3(_0112_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2219_ (.A1(_0091_),
    .A2(_0104_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2220_ (.A1(_0105_),
    .A2(_0113_),
    .B(_0114_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2221_ (.A1(_0092_),
    .A2(_0102_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2222_ (.A1(_0692_),
    .A2(_0103_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2223_ (.A1(_0116_),
    .A2(_0117_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2224_ (.A1(_0093_),
    .A2(_0101_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2225_ (.A1(_0093_),
    .A2(_0101_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2226_ (.A1(_0095_),
    .A2(_0119_),
    .B(_0120_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2227_ (.I(\c[0][4] ),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2228_ (.A1(_0122_),
    .A2(_1356_),
    .A3(_0657_),
    .A4(_0973_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2229_ (.A1(_0122_),
    .A2(_0658_),
    .B1(_0973_),
    .B2(_1356_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2230_ (.A1(_0123_),
    .A2(_0124_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2231_ (.A1(_0098_),
    .A2(_0100_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2232_ (.A1(_0098_),
    .A2(_0100_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2233_ (.A1(_0096_),
    .A2(_0126_),
    .B(_0127_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2234_ (.A1(\c[0][1] ),
    .A2(_0835_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2235_ (.I(\c[0][3] ),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2236_ (.A1(_0130_),
    .A2(\c[0][2] ),
    .A3(_0642_),
    .A4(_0705_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2237_ (.A1(_0130_),
    .A2(_0643_),
    .B1(_0705_),
    .B2(_0097_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2238_ (.A1(_0131_),
    .A2(_0132_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2239_ (.A1(_0129_),
    .A2(_0133_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2240_ (.A1(_0128_),
    .A2(_0134_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2241_ (.A1(_0125_),
    .A2(_0135_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2242_ (.A1(_0121_),
    .A2(_0136_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2243_ (.A1(_0764_),
    .A2(_0137_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2244_ (.A1(_0115_),
    .A2(_0118_),
    .A3(_0138_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2245_ (.A1(_0716_),
    .A2(_0139_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2246_ (.A1(_0118_),
    .A2(_0138_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2247_ (.A1(_0118_),
    .A2(_0138_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2248_ (.A1(_0115_),
    .A2(_0141_),
    .B(_0142_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2249_ (.A1(_0764_),
    .A2(_0137_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2250_ (.A1(_0121_),
    .A2(_0136_),
    .B(_0144_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2251_ (.A1(_0798_),
    .A2(_0828_),
    .A3(_0123_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2252_ (.A1(_0128_),
    .A2(_0134_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2253_ (.A1(_0125_),
    .A2(_0135_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2254_ (.A1(_0147_),
    .A2(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2255_ (.A1(_0129_),
    .A2(_0133_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2256_ (.A1(_0131_),
    .A2(_0150_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2257_ (.A1(_0099_),
    .A2(_0647_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2258_ (.A1(_0097_),
    .A2(_0835_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2259_ (.A1(_0078_),
    .A2(_0928_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2260_ (.A1(_0152_),
    .A2(_0153_),
    .A3(_0154_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2261_ (.A1(_0151_),
    .A2(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2262_ (.I(\c[0][5] ),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2263_ (.A1(_0157_),
    .A2(_0658_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2264_ (.A1(\c[0][0] ),
    .A2(_0922_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2265_ (.A1(\c[0][4] ),
    .A2(_0652_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2266_ (.A1(_0159_),
    .A2(_0160_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2267_ (.A1(_0158_),
    .A2(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2268_ (.A1(_0156_),
    .A2(_0162_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2269_ (.A1(_0149_),
    .A2(_0163_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2270_ (.A1(_0145_),
    .A2(_0146_),
    .A3(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2271_ (.A1(_0143_),
    .A2(_0165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2272_ (.A1(_0808_),
    .A2(_0166_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2273_ (.A1(_0140_),
    .A2(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2274_ (.I(_0168_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2275_ (.A1(_0140_),
    .A2(_0167_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2276_ (.A1(_0713_),
    .A2(_0166_),
    .B(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2277_ (.A1(_0870_),
    .A2(_0123_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2278_ (.A1(_0149_),
    .A2(_0163_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2279_ (.A1(_0146_),
    .A2(_0164_),
    .B(_0172_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2280_ (.I(_0159_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2281_ (.A1(_0174_),
    .A2(_0160_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2282_ (.A1(_0158_),
    .A2(_0161_),
    .B(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2283_ (.A1(\c[0][6] ),
    .A2(_0693_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2284_ (.A1(_0879_),
    .A2(_0983_),
    .A3(_0177_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2285_ (.A1(_0151_),
    .A2(_0155_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2286_ (.A1(_0156_),
    .A2(_0162_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2287_ (.A1(_0179_),
    .A2(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2288_ (.A1(_0152_),
    .A2(_0153_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2289_ (.A1(_0152_),
    .A2(_0153_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2290_ (.A1(_0182_),
    .A2(_0154_),
    .B(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2291_ (.A1(\c[0][1] ),
    .A2(_0841_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2292_ (.I(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2293_ (.A1(_0130_),
    .A2(_0703_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2294_ (.A1(_0080_),
    .A2(_0777_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2295_ (.A1(_0186_),
    .A2(_0187_),
    .A3(_0188_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2296_ (.A1(_0184_),
    .A2(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(\c[0][5] ),
    .A2(_0653_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2298_ (.A1(\c[0][4] ),
    .A2(_0647_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2299_ (.A1(_0159_),
    .A2(_0192_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2300_ (.A1(_0191_),
    .A2(_0193_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2301_ (.A1(_0190_),
    .A2(_0194_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2302_ (.I(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2303_ (.A1(_0181_),
    .A2(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2304_ (.A1(_0176_),
    .A2(_0178_),
    .A3(_0197_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2305_ (.A1(_0171_),
    .A2(_0173_),
    .A3(_0198_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2306_ (.A1(_0146_),
    .A2(_0164_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2307_ (.A1(_0143_),
    .A2(_0165_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2308_ (.A1(_0145_),
    .A2(_0200_),
    .B(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2309_ (.A1(_0199_),
    .A2(_0202_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2310_ (.A1(_0864_),
    .A2(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2311_ (.A1(_0170_),
    .A2(_0204_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2312_ (.I(_0205_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2313_ (.A1(_0170_),
    .A2(_0204_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2314_ (.A1(_0865_),
    .A2(_0203_),
    .B(_0206_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2315_ (.A1(_0199_),
    .A2(_0202_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2316_ (.A1(_0176_),
    .A2(_0178_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2317_ (.A1(_0173_),
    .A2(_0198_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2318_ (.A1(_0173_),
    .A2(_0198_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2319_ (.A1(_0171_),
    .A2(_0210_),
    .B(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2320_ (.A1(_0176_),
    .A2(_0178_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2321_ (.A1(_0181_),
    .A2(_0196_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2322_ (.A1(_0213_),
    .A2(_0197_),
    .B(_0214_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2323_ (.A1(_0184_),
    .A2(_0189_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2324_ (.A1(_0190_),
    .A2(_0194_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2325_ (.A1(_0187_),
    .A2(_0188_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2326_ (.A1(_0187_),
    .A2(_0188_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2327_ (.A1(_0186_),
    .A2(_0218_),
    .B(_0219_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2328_ (.A1(_0130_),
    .A2(_0777_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2329_ (.A1(_0097_),
    .A2(_0922_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2330_ (.A1(_0221_),
    .A2(_0222_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2331_ (.A1(_0186_),
    .A2(_0223_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2332_ (.A1(_0220_),
    .A2(_0224_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2333_ (.A1(_0220_),
    .A2(_0224_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2334_ (.A1(_0225_),
    .A2(_0226_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2335_ (.A1(\c[0][5] ),
    .A2(_0969_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2336_ (.A1(_0122_),
    .A2(_1047_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2337_ (.A1(_0174_),
    .A2(_0228_),
    .A3(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2338_ (.A1(_0227_),
    .A2(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2339_ (.A1(_0216_),
    .A2(_0217_),
    .B(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2340_ (.A1(_0216_),
    .A2(_0217_),
    .A3(_0231_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2341_ (.A1(_0232_),
    .A2(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2342_ (.A1(_0952_),
    .A2(_0177_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2343_ (.I(_0174_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2344_ (.A1(_0191_),
    .A2(_0193_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2345_ (.A1(_0236_),
    .A2(_0192_),
    .B(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2346_ (.A1(\c[0][6] ),
    .A2(_0654_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2347_ (.A1(\c[0][7] ),
    .A2(_0693_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2348_ (.A1(_0239_),
    .A2(_0240_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2349_ (.A1(_0985_),
    .A2(_1016_),
    .A3(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2350_ (.A1(_0235_),
    .A2(_0238_),
    .A3(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2351_ (.A1(_0215_),
    .A2(_0234_),
    .A3(_0243_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2352_ (.A1(_0209_),
    .A2(_0212_),
    .A3(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2353_ (.A1(_0208_),
    .A2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2354_ (.A1(_0897_),
    .A2(_0246_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2355_ (.A1(_0207_),
    .A2(_0247_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2356_ (.I(_0248_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2357_ (.A1(_0673_),
    .A2(_0246_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2358_ (.A1(_0207_),
    .A2(_0247_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2359_ (.A1(_0209_),
    .A2(_0244_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2360_ (.A1(_0199_),
    .A2(_0202_),
    .A3(_0245_),
    .B1(_0251_),
    .B2(_0212_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2361_ (.A1(_0234_),
    .A2(_0243_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2362_ (.A1(_0176_),
    .A2(net82),
    .A3(_0244_),
    .B1(_0253_),
    .B2(net76),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2363_ (.A1(_0238_),
    .A2(_0242_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2364_ (.A1(_0238_),
    .A2(_0242_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2365_ (.A1(_0235_),
    .A2(_0255_),
    .B(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2366_ (.A1(_0234_),
    .A2(_0243_),
    .B(_0232_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2367_ (.A1(_0227_),
    .A2(_0230_),
    .B(_0225_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2368_ (.I(_0099_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2369_ (.A1(_0260_),
    .A2(_0084_),
    .A3(_0222_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2370_ (.A1(_0099_),
    .A2(_0080_),
    .B(_1130_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2371_ (.A1(_0260_),
    .A2(_0222_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2372_ (.A1(_0185_),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2373_ (.A1(_0260_),
    .A2(_1137_),
    .A3(_0222_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2374_ (.A1(_0185_),
    .A2(_0223_),
    .B(_0264_),
    .C(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2375_ (.A1(_0261_),
    .A2(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2376_ (.I(_0157_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2377_ (.A1(_0268_),
    .A2(net93),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2378_ (.I(_0122_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2379_ (.A1(_0270_),
    .A2(_1136_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2380_ (.A1(_0174_),
    .A2(_0271_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2381_ (.A1(_0269_),
    .A2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2382_ (.A1(_0267_),
    .A2(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2383_ (.A1(_0259_),
    .A2(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2384_ (.A1(_0985_),
    .A2(_1016_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2385_ (.A1(_0239_),
    .A2(_0240_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2386_ (.A1(_0276_),
    .A2(_0241_),
    .B(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2387_ (.I(_0228_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2388_ (.A1(_0236_),
    .A2(_0229_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2389_ (.A1(_0236_),
    .A2(_0229_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2390_ (.A1(_0279_),
    .A2(_0280_),
    .B(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2391_ (.I(\c[0][7] ),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2392_ (.A1(_0283_),
    .A2(_0655_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2393_ (.I(\c[0][6] ),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2394_ (.A1(_0285_),
    .A2(_1100_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2395_ (.A1(_0284_),
    .A2(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2396_ (.A1(_1066_),
    .A2(_1098_),
    .A3(_0287_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2397_ (.A1(_0278_),
    .A2(_0282_),
    .A3(_0288_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2398_ (.A1(_0258_),
    .A2(_0275_),
    .A3(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2399_ (.A1(_0254_),
    .A2(_0257_),
    .A3(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2400_ (.A1(_1029_),
    .A2(_0252_),
    .A3(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2401_ (.A1(_0249_),
    .A2(_0250_),
    .B(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2402_ (.A1(_0249_),
    .A2(_0250_),
    .A3(_0292_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2403_ (.A1(_0293_),
    .A2(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2404_ (.I(_0295_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2405_ (.I(_1113_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2406_ (.A1(_0252_),
    .A2(_0291_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2407_ (.A1(_0252_),
    .A2(_0291_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2408_ (.A1(_1082_),
    .A2(_0297_),
    .A3(_0298_),
    .B(_0293_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2409_ (.A1(_0257_),
    .A2(_0290_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2410_ (.A1(net81),
    .A2(_0300_),
    .B(_0297_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2411_ (.A1(_0275_),
    .A2(_0289_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2412_ (.A1(_0257_),
    .A2(_0290_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2413_ (.A1(_0258_),
    .A2(_0302_),
    .B(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2414_ (.I(_0282_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2415_ (.A1(_0282_),
    .A2(_0288_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2416_ (.A1(_0278_),
    .A2(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2417_ (.A1(_0305_),
    .A2(_0288_),
    .B(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2418_ (.A1(_0259_),
    .A2(_0274_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2419_ (.A1(_0275_),
    .A2(_0289_),
    .B(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2420_ (.A1(_0267_),
    .A2(_0273_),
    .B(_0261_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2421_ (.A1(_0185_),
    .A2(_0262_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2422_ (.A1(_0261_),
    .A2(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2423_ (.A1(_0157_),
    .A2(_1136_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2424_ (.A1(_0270_),
    .A2(_0085_),
    .A3(_1130_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2425_ (.A1(_0270_),
    .A2(_0085_),
    .B1(_0906_),
    .B2(_0907_),
    .C(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2426_ (.A1(_0314_),
    .A2(_0316_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2427_ (.A1(_0313_),
    .A2(_0317_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2428_ (.A1(_0311_),
    .A2(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2429_ (.I(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2430_ (.A1(_0284_),
    .A2(_0286_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2431_ (.A1(_1142_),
    .A2(_0287_),
    .B(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2432_ (.A1(_0236_),
    .A2(_0271_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2433_ (.A1(_0269_),
    .A2(_0272_),
    .B(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2434_ (.A1(\c[0][7] ),
    .A2(_1100_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(\c[0][6] ),
    .A2(_1047_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2436_ (.A1(_0325_),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2437_ (.A1(_1150_),
    .A2(_1180_),
    .A3(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2438_ (.A1(_0322_),
    .A2(_0324_),
    .A3(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2439_ (.A1(_0310_),
    .A2(_0320_),
    .A3(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2440_ (.A1(_0308_),
    .A2(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2441_ (.A1(_0301_),
    .A2(_0304_),
    .A3(_0331_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2442_ (.A1(_0296_),
    .A2(_0299_),
    .A3(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2443_ (.I(_0333_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(_1197_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2445_ (.A1(_0296_),
    .A2(_0332_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2446_ (.A1(_0332_),
    .A2(_0296_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2447_ (.A1(_0299_),
    .A2(_0335_),
    .B(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2448_ (.A1(_0304_),
    .A2(_0331_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2449_ (.A1(_0304_),
    .A2(_0331_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2450_ (.A1(_0301_),
    .A2(_0338_),
    .B(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2451_ (.A1(_0319_),
    .A2(_0329_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2452_ (.A1(_0310_),
    .A2(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2453_ (.A1(_0308_),
    .A2(_0330_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2454_ (.A1(_0342_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2455_ (.A1(_1205_),
    .A2(_0327_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2456_ (.A1(_0324_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2457_ (.A1(_0324_),
    .A2(_0328_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2458_ (.A1(_0322_),
    .A2(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2459_ (.A1(_0346_),
    .A2(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2460_ (.A1(_0311_),
    .A2(_0318_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2461_ (.A1(_0320_),
    .A2(_0329_),
    .B(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2462_ (.A1(_0325_),
    .A2(_0326_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2463_ (.A1(_0325_),
    .A2(_0326_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2464_ (.A1(_1205_),
    .A2(_0352_),
    .B(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2465_ (.I(_0316_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2466_ (.A1(_0314_),
    .A2(_0355_),
    .B(_0315_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2467_ (.A1(_0283_),
    .A2(_1184_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2468_ (.A1(_0285_),
    .A2(_1137_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2469_ (.A1(_0357_),
    .A2(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2470_ (.A1(_1220_),
    .A2(_1242_),
    .A3(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2471_ (.A1(_0354_),
    .A2(_0356_),
    .A3(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2472_ (.I(_0261_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2473_ (.A1(_0313_),
    .A2(_0317_),
    .B(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2474_ (.A1(_0157_),
    .A2(_1285_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2475_ (.A1(_0355_),
    .A2(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2476_ (.A1(_0268_),
    .A2(_0355_),
    .B(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2477_ (.A1(_0313_),
    .A2(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2478_ (.A1(_0363_),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2479_ (.A1(_0351_),
    .A2(_0361_),
    .A3(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2480_ (.A1(_0349_),
    .A2(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2481_ (.A1(_0344_),
    .A2(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2482_ (.A1(_0340_),
    .A2(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2483_ (.A1(_0334_),
    .A2(_0337_),
    .A3(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2484_ (.I(_0373_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2485_ (.A1(_0334_),
    .A2(_0372_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(_0334_),
    .A2(_0372_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2487_ (.A1(_0337_),
    .A2(_0374_),
    .B(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2488_ (.A1(_0340_),
    .A2(_0371_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2489_ (.A1(_0344_),
    .A2(_0370_),
    .B(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2490_ (.A1(_0361_),
    .A2(_0368_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2491_ (.A1(_0351_),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2492_ (.A1(_0349_),
    .A2(_0369_),
    .B(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2493_ (.A1(_0283_),
    .A2(_1244_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2494_ (.A1(_0357_),
    .A2(_0358_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2495_ (.A1(_0357_),
    .A2(_0358_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2496_ (.A1(_1290_),
    .A2(_0383_),
    .B(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2497_ (.A1(_0382_),
    .A2(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2498_ (.A1(_0285_),
    .A2(_1285_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2499_ (.I(_0363_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(_0388_),
    .A2(_0367_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2501_ (.A1(_0361_),
    .A2(_0368_),
    .B(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2502_ (.A1(_0356_),
    .A2(_0360_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2503_ (.A1(_0356_),
    .A2(_0360_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2504_ (.A1(_0354_),
    .A2(_0391_),
    .B(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2505_ (.A1(_0268_),
    .A2(_0355_),
    .B(_0315_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2506_ (.A1(_0312_),
    .A2(_0366_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2507_ (.A1(_0362_),
    .A2(_0366_),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2508_ (.A1(_0394_),
    .A2(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2509_ (.A1(_1289_),
    .A2(_0393_),
    .A3(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2510_ (.A1(_0387_),
    .A2(_0390_),
    .A3(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2511_ (.A1(_0381_),
    .A2(_0386_),
    .A3(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2512_ (.A1(_1261_),
    .A2(_0378_),
    .A3(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2513_ (.A1(_0376_),
    .A2(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2514_ (.I(_0402_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2515_ (.A1(_0716_),
    .A2(_0139_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2516_ (.I(_0403_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2517_ (.I(net4),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2518_ (.I(net3),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2519_ (.A1(net28),
    .A2(net37),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2520_ (.A1(_0404_),
    .A2(_0405_),
    .A3(net25),
    .A4(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2521_ (.A1(net22),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2522_ (.I(net2),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2523_ (.I(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2524_ (.A1(_0679_),
    .A2(_0407_),
    .B(_0408_),
    .C(_0410_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2525_ (.A1(net23),
    .A2(_0407_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2526_ (.A1(_1349_),
    .A2(_0407_),
    .B(_0411_),
    .C(_0410_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2527_ (.A1(net4),
    .A2(net3),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2528_ (.A1(net24),
    .A2(_0406_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2529_ (.I(_0413_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2530_ (.A1(_0412_),
    .A2(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2531_ (.I(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2532_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2533_ (.A1(\delta_t[0] ),
    .A2(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2534_ (.I(_0413_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2535_ (.A1(_0412_),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2536_ (.A1(net6),
    .A2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2537_ (.I(_0409_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2538_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2539_ (.A1(_0418_),
    .A2(_0421_),
    .B(_0423_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2540_ (.I(_0416_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2541_ (.I(_0415_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2542_ (.A1(net11),
    .A2(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2543_ (.A1(_1314_),
    .A2(_0424_),
    .B(_0426_),
    .C(_0410_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2544_ (.A1(net16),
    .A2(_0425_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2545_ (.I(net2),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2546_ (.I(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2547_ (.A1(_0589_),
    .A2(_0424_),
    .B(_0427_),
    .C(_0429_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2548_ (.A1(net17),
    .A2(_0425_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2549_ (.A1(_0596_),
    .A2(_0424_),
    .B(_0430_),
    .C(_0429_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2550_ (.A1(net18),
    .A2(_0425_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2551_ (.A1(_1325_),
    .A2(_0424_),
    .B(_0431_),
    .C(_0429_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2552_ (.A1(net19),
    .A2(_0416_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2553_ (.A1(_1330_),
    .A2(_0417_),
    .B(_0432_),
    .C(_0429_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2554_ (.A1(_1335_),
    .A2(_0417_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2555_ (.A1(net20),
    .A2(_0420_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2556_ (.A1(_0433_),
    .A2(_0434_),
    .B(_0423_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2557_ (.A1(net21),
    .A2(_0416_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2558_ (.I(_0409_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2559_ (.A1(_0747_),
    .A2(_0417_),
    .B(_0435_),
    .C(_0436_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2560_ (.I(net7),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2561_ (.A1(net26),
    .A2(_0406_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2562_ (.I(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2563_ (.A1(_0412_),
    .A2(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2564_ (.A1(_0573_),
    .A2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2565_ (.A1(_0437_),
    .A2(_0440_),
    .B(_0441_),
    .C(_0436_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2566_ (.I(net3),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2567_ (.A1(net4),
    .A2(_0442_),
    .A3(_0414_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2568_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2569_ (.I(_0443_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2570_ (.A1(net6),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2571_ (.A1(_0553_),
    .A2(_0444_),
    .B(_0446_),
    .C(_0436_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2572_ (.A1(net11),
    .A2(_0445_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2573_ (.A1(_0808_),
    .A2(_0444_),
    .B(_0447_),
    .C(_0436_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2574_ (.I(_0443_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2575_ (.A1(_0865_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2576_ (.A1(_0404_),
    .A2(_0405_),
    .A3(_0419_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2577_ (.A1(net16),
    .A2(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2578_ (.A1(_0449_),
    .A2(_0451_),
    .B(_0423_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2579_ (.A1(net17),
    .A2(_0445_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2580_ (.I(_0409_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2581_ (.A1(_0897_),
    .A2(_0444_),
    .B(_0452_),
    .C(_0453_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2582_ (.A1(net18),
    .A2(_0445_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2583_ (.A1(_1082_),
    .A2(_0444_),
    .B(_0454_),
    .C(_0453_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2584_ (.A1(net19),
    .A2(_0443_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2585_ (.A1(_0296_),
    .A2(_0448_),
    .B(_0455_),
    .C(_0453_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2586_ (.A1(_0334_),
    .A2(_0448_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2587_ (.A1(net20),
    .A2(_0450_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2588_ (.A1(_0456_),
    .A2(_0457_),
    .B(_0423_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2589_ (.A1(_1261_),
    .A2(_0448_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2590_ (.A1(net21),
    .A2(_0450_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2591_ (.I(net2),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2592_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2593_ (.A1(_0458_),
    .A2(_0459_),
    .B(_0461_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2594_ (.A1(_0404_),
    .A2(_0442_),
    .A3(_0438_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2595_ (.I(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2596_ (.A1(\a[1][0] ),
    .A2(_0462_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2597_ (.A1(_0437_),
    .A2(_0463_),
    .B(_0464_),
    .C(_0453_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2598_ (.A1(_0404_),
    .A2(_0442_),
    .A3(_0439_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2599_ (.I(_0465_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2600_ (.A1(\a[1][1] ),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2601_ (.A1(net8),
    .A2(_0463_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2602_ (.A1(_0467_),
    .A2(_0468_),
    .B(_0461_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2603_ (.A1(\a[1][2] ),
    .A2(_0466_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2604_ (.A1(net9),
    .A2(_0463_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2605_ (.A1(_0469_),
    .A2(_0470_),
    .B(_0461_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2606_ (.A1(\a[1][3] ),
    .A2(_0466_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2607_ (.A1(net10),
    .A2(_0463_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2608_ (.A1(_0471_),
    .A2(_0472_),
    .B(_0461_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2609_ (.A1(\a[1][4] ),
    .A2(_0466_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2610_ (.I(_0462_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2611_ (.A1(net12),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2612_ (.I(_0460_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2613_ (.A1(_0473_),
    .A2(_0475_),
    .B(_0476_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2614_ (.A1(\a[1][5] ),
    .A2(_0465_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2615_ (.A1(net13),
    .A2(_0474_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2616_ (.A1(_0477_),
    .A2(_0478_),
    .B(_0476_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2617_ (.A1(\a[1][6] ),
    .A2(_0465_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2618_ (.A1(net14),
    .A2(_0474_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2619_ (.A1(_0479_),
    .A2(_0480_),
    .B(_0476_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2620_ (.A1(\a[1][7] ),
    .A2(_0465_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(net15),
    .A2(_0474_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2622_ (.A1(_0481_),
    .A2(_0482_),
    .B(_0476_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2623_ (.I(net4),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2624_ (.A1(_0483_),
    .A2(_0442_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2625_ (.A1(_0414_),
    .A2(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2626_ (.I(_0485_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2627_ (.A1(_0660_),
    .A2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2628_ (.A1(_0419_),
    .A2(_0484_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2629_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2630_ (.A1(net6),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2631_ (.I(_0460_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2632_ (.A1(_0487_),
    .A2(_0490_),
    .B(_0491_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2633_ (.A1(_0651_),
    .A2(_0486_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2634_ (.A1(net11),
    .A2(_0489_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2635_ (.A1(_0492_),
    .A2(_0493_),
    .B(_0491_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2636_ (.A1(_0927_),
    .A2(_0486_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2637_ (.A1(net16),
    .A2(_0489_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2638_ (.A1(_0494_),
    .A2(_0495_),
    .B(_0491_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_0972_),
    .A2(_0486_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2640_ (.A1(net17),
    .A2(_0489_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2641_ (.A1(_0496_),
    .A2(_0497_),
    .B(_0491_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2642_ (.I(_0485_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2643_ (.A1(_0794_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2644_ (.I(_0488_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2645_ (.A1(net18),
    .A2(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2646_ (.I(_0460_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2647_ (.A1(_0499_),
    .A2(_0501_),
    .B(_0502_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2648_ (.A1(_1046_),
    .A2(_0498_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2649_ (.A1(net19),
    .A2(_0500_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2650_ (.A1(_0503_),
    .A2(_0504_),
    .B(_0502_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2651_ (.A1(_1183_),
    .A2(_0498_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2652_ (.A1(net20),
    .A2(_0500_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2653_ (.A1(_0505_),
    .A2(_0506_),
    .B(_0502_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2654_ (.A1(_1181_),
    .A2(_0498_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2655_ (.A1(net21),
    .A2(_0500_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2656_ (.A1(_0507_),
    .A2(_0508_),
    .B(_0502_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2657_ (.A1(_0439_),
    .A2(_0484_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2658_ (.I(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2659_ (.A1(\b[1][0] ),
    .A2(_0509_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2660_ (.A1(_0437_),
    .A2(_0510_),
    .B(_0511_),
    .C(_0422_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2661_ (.A1(_0439_),
    .A2(_0484_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2662_ (.I(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2663_ (.A1(\b[1][1] ),
    .A2(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2664_ (.A1(net8),
    .A2(_0510_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2665_ (.I(_0428_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2666_ (.A1(_0514_),
    .A2(_0515_),
    .B(_0516_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2667_ (.A1(\b[1][2] ),
    .A2(_0513_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2668_ (.A1(net9),
    .A2(_0510_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2669_ (.A1(_0517_),
    .A2(_0518_),
    .B(_0516_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2670_ (.A1(\b[1][3] ),
    .A2(_0513_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2671_ (.A1(net10),
    .A2(_0510_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2672_ (.A1(_0519_),
    .A2(_0520_),
    .B(_0516_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(\b[1][4] ),
    .A2(_0513_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2674_ (.I(_0509_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2675_ (.A1(net12),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2676_ (.A1(_0521_),
    .A2(_0523_),
    .B(_0516_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2677_ (.A1(\b[1][5] ),
    .A2(_0512_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2678_ (.A1(net13),
    .A2(_0522_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2679_ (.I(_0428_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2680_ (.A1(_0524_),
    .A2(_0525_),
    .B(_0526_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2681_ (.A1(\b[1][6] ),
    .A2(_0512_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2682_ (.A1(net14),
    .A2(_0522_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2683_ (.A1(_0527_),
    .A2(_0528_),
    .B(_0526_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2684_ (.A1(\b[1][7] ),
    .A2(_0512_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(net15),
    .A2(_0522_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2686_ (.A1(_0529_),
    .A2(_0530_),
    .B(_0526_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2687_ (.A1(_0483_),
    .A2(_0405_),
    .A3(_0414_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2688_ (.I(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2689_ (.A1(net6),
    .A2(_0531_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2690_ (.A1(_0094_),
    .A2(_0532_),
    .B(_0533_),
    .C(_0422_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2691_ (.A1(_0084_),
    .A2(_0532_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2692_ (.A1(_0483_),
    .A2(_0405_),
    .A3(_0419_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2693_ (.I(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2694_ (.A1(net11),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2695_ (.A1(_0534_),
    .A2(_0537_),
    .B(_0526_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2696_ (.A1(_0080_),
    .A2(_0532_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2697_ (.A1(net16),
    .A2(_0536_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2698_ (.I(_0428_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2699_ (.A1(_0538_),
    .A2(_0539_),
    .B(_0540_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2700_ (.I(_0531_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2701_ (.A1(_0260_),
    .A2(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2702_ (.A1(net17),
    .A2(_0536_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2703_ (.A1(_0542_),
    .A2(_0543_),
    .B(_0540_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2704_ (.A1(_0270_),
    .A2(_0541_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2705_ (.A1(net18),
    .A2(_0536_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2706_ (.A1(_0544_),
    .A2(_0545_),
    .B(_0540_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2707_ (.A1(net19),
    .A2(_0531_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2708_ (.A1(_0268_),
    .A2(_0532_),
    .B(_0546_),
    .C(_0422_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2709_ (.A1(_0285_),
    .A2(_0541_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2710_ (.A1(net20),
    .A2(_0535_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2711_ (.A1(_0547_),
    .A2(_0548_),
    .B(_0540_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2712_ (.A1(_0283_),
    .A2(_0541_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2713_ (.A1(net21),
    .A2(_0535_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2714_ (.A1(_0549_),
    .A2(_0550_),
    .B(_0410_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2715_ (.D(_0026_),
    .CLK(net54),
    .Q(\delta_t[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2716_ (.D(_0027_),
    .CLK(net55),
    .Q(\delta_t[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2717_ (.D(_0000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2718_ (.D(_0001_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2719_ (.D(_0002_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2720_ (.D(_0003_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2721_ (.D(_0004_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2722_ (.D(_0005_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2723_ (.D(_0006_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2724_ (.D(_0007_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2725_ (.D(_0008_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2726_ (.D(_0009_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2727_ (.D(_0010_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2728_ (.D(_0011_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2729_ (.D(_0012_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2730_ (.D(_0013_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2731_ (.D(_0014_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2732_ (.D(_0015_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2733_ (.D(_0016_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2734_ (.D(_0017_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2735_ (.D(_0018_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2736_ (.D(_0019_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2737_ (.D(_0020_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2738_ (.D(_0021_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2739_ (.D(_0022_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2740_ (.D(_0023_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2741_ (.D(_0024_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2742_ (.D(_0025_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2743_ (.D(_0028_),
    .CLK(net58),
    .Q(\delta_t[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2744_ (.D(_0029_),
    .CLK(net56),
    .Q(\delta_t[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2745_ (.D(_0030_),
    .CLK(net54),
    .Q(\delta_t[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2746_ (.D(_0031_),
    .CLK(net54),
    .Q(\delta_t[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2747_ (.D(_0032_),
    .CLK(net54),
    .Q(\delta_t[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2748_ (.D(_0033_),
    .CLK(net55),
    .Q(\delta_t[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2749_ (.D(_0034_),
    .CLK(net57),
    .Q(\delta_t[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2750_ (.D(_0035_),
    .CLK(net55),
    .Q(\delta_t[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2751_ (.D(_0036_),
    .CLK(net61),
    .Q(bflip));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2752_ (.D(_0037_),
    .CLK(net57),
    .Q(\a[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2753_ (.D(_0038_),
    .CLK(net57),
    .Q(\a[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2754_ (.D(_0039_),
    .CLK(net58),
    .Q(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2755_ (.D(_0040_),
    .CLK(net57),
    .Q(\a[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2756_ (.D(_0041_),
    .CLK(net59),
    .Q(\a[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2757_ (.D(_0042_),
    .CLK(net58),
    .Q(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2758_ (.D(_0043_),
    .CLK(net59),
    .Q(\a[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2759_ (.D(_0044_),
    .CLK(net58),
    .Q(\a[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2760_ (.D(_0045_),
    .CLK(net56),
    .Q(\a[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2761_ (.D(_0046_),
    .CLK(net62),
    .Q(\a[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2762_ (.D(_0047_),
    .CLK(net64),
    .Q(\a[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2763_ (.D(_0048_),
    .CLK(net61),
    .Q(\a[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2764_ (.D(_0049_),
    .CLK(net64),
    .Q(\a[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2765_ (.D(_0050_),
    .CLK(net66),
    .Q(\a[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2766_ (.D(_0051_),
    .CLK(net65),
    .Q(\a[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2767_ (.D(_0052_),
    .CLK(net66),
    .Q(\a[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2768_ (.D(_0053_),
    .CLK(net73),
    .Q(\b[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2769_ (.D(_0054_),
    .CLK(net73),
    .Q(\b[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2770_ (.D(_0055_),
    .CLK(net73),
    .Q(\b[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2771_ (.D(_0056_),
    .CLK(net73),
    .Q(\b[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2772_ (.D(_0057_),
    .CLK(net63),
    .Q(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2773_ (.D(_0058_),
    .CLK(net69),
    .Q(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2774_ (.D(_0059_),
    .CLK(net70),
    .Q(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2775_ (.D(_0060_),
    .CLK(net67),
    .Q(\b[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2776_ (.D(_0061_),
    .CLK(net61),
    .Q(\b[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2777_ (.D(_0062_),
    .CLK(net62),
    .Q(\b[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2778_ (.D(_0063_),
    .CLK(net64),
    .Q(\b[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2779_ (.D(_0064_),
    .CLK(net61),
    .Q(\b[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2780_ (.D(_0065_),
    .CLK(net64),
    .Q(\b[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2781_ (.D(_0066_),
    .CLK(net65),
    .Q(\b[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2782_ (.D(_0067_),
    .CLK(net65),
    .Q(\b[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2783_ (.D(_0068_),
    .CLK(net67),
    .Q(\b[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2784_ (.D(_0069_),
    .CLK(net74),
    .Q(\c[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2785_ (.D(_0070_),
    .CLK(net63),
    .Q(\c[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2786_ (.D(_0071_),
    .CLK(net69),
    .Q(\c[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2787_ (.D(_0072_),
    .CLK(net69),
    .Q(\c[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2788_ (.D(_0073_),
    .CLK(net70),
    .Q(\c[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2789_ (.D(_0074_),
    .CLK(net74),
    .Q(\c[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2790_ (.D(_0075_),
    .CLK(net69),
    .Q(\c[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2791_ (.D(_0076_),
    .CLK(net68),
    .Q(\c[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout54 (.I(net56),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout56 (.I(net60),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout57 (.I(net59),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout59 (.I(net60),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout60 (.I(net72),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout61 (.I(net63),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout62 (.I(net63),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout63 (.I(net68),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout64 (.I(net66),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout66 (.I(net68),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout68 (.I(net71),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout70 (.I(net71),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout72 (.I(net75),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout73 (.I(net75),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout75 (.I(net1),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(wb_clk_i),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(wbs_dat_i[19]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(wbs_dat_i[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(wbs_dat_i[20]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(wbs_dat_i[21]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(wbs_dat_i[22]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(wbs_dat_i[23]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(wbs_dat_i[2]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input17 (.I(wbs_dat_i[3]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(wbs_dat_i[4]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input19 (.I(wbs_dat_i[5]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(wb_rst_i),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input20 (.I(wbs_dat_i[6]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input21 (.I(wbs_dat_i[7]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(wbs_dat_i[8]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(wbs_dat_i[9]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(wbs_sel_i[0]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input25 (.I(wbs_sel_i[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(wbs_sel_i[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(wbs_stb_i),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(wbs_we_i),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(y[0]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input3 (.I(wbs_adr_i[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(y[1]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(y[2]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(y[3]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(y[4]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(y[5]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(y[6]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(y[7]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input4 (.I(wbs_adr_i[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(wbs_cyc_i),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input6 (.I(wbs_dat_i[0]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(wbs_dat_i[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(wbs_dat_i[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(wbs_dat_i[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output37 (.I(net37),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(x_end[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output39 (.I(net39),
    .Z(x_end[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output40 (.I(net40),
    .Z(x_end[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output41 (.I(net41),
    .Z(x_end[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output42 (.I(net42),
    .Z(x_end[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output43 (.I(net43),
    .Z(x_end[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output44 (.I(net44),
    .Z(x_end[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(x_end[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(x_start[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output47 (.I(net47),
    .Z(x_start[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output48 (.I(net48),
    .Z(x_start[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output49 (.I(net49),
    .Z(x_start[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output50 (.I(net50),
    .Z(x_start[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(x_start[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output52 (.I(net52),
    .Z(x_start[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output53 (.I(net53),
    .Z(x_start[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer1 (.I(_0215_),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(_0806_),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(net92),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(net100),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer13 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer14 (.I(_0685_),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(_0880_),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(net90),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer17 (.I(_0802_),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer18 (.I(_0735_),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer19 (.I(net98),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer2 (.I(_0587_),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer20 (.I(_0826_),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer21 (.I(_0802_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer22 (.I(_0826_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer23 (.I(_0582_),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer24 (.I(_0811_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer25 (.I(_0759_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(_0631_),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(net78),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_0612_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(_0254_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(_0178_),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer8 (.I(_0599_),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(_0797_),
    .Z(net84));
endmodule

