VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpu_core
  CLASS BLOCK ;
  FOREIGN gpu_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 4000.000 ;
  PIN ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1952.160 4.000 1952.720 ;
    END
  END ack
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2520.000 4.000 2520.560 ;
    END
  END clk
  PIN cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1975.680 4.000 1976.240 ;
    END
  END cyc
  PIN dat_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2456.160 2500.000 2456.720 ;
    END
  END dat_in[0]
  PIN dat_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1575.840 2500.000 1576.400 ;
    END
  END dat_in[10]
  PIN dat_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1552.320 2500.000 1552.880 ;
    END
  END dat_in[11]
  PIN dat_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1632.960 2500.000 1633.520 ;
    END
  END dat_in[12]
  PIN dat_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1619.520 2500.000 1620.080 ;
    END
  END dat_in[13]
  PIN dat_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1629.600 2500.000 1630.160 ;
    END
  END dat_in[14]
  PIN dat_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1626.240 2500.000 1626.800 ;
    END
  END dat_in[15]
  PIN dat_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2352.000 4.000 2352.560 ;
    END
  END dat_in[16]
  PIN dat_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2304.960 2500.000 2305.520 ;
    END
  END dat_in[17]
  PIN dat_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2308.320 2500.000 2308.880 ;
    END
  END dat_in[18]
  PIN dat_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2288.160 4.000 2288.720 ;
    END
  END dat_in[19]
  PIN dat_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2442.720 2500.000 2443.280 ;
    END
  END dat_in[1]
  PIN dat_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2116.800 2500.000 2117.360 ;
    END
  END dat_in[20]
  PIN dat_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2103.360 2500.000 2103.920 ;
    END
  END dat_in[21]
  PIN dat_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2073.120 2500.000 2073.680 ;
    END
  END dat_in[22]
  PIN dat_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2056.320 2500.000 2056.880 ;
    END
  END dat_in[23]
  PIN dat_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1817.760 2500.000 1818.320 ;
    END
  END dat_in[24]
  PIN dat_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1757.280 2500.000 1757.840 ;
    END
  END dat_in[25]
  PIN dat_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1760.640 2500.000 1761.200 ;
    END
  END dat_in[26]
  PIN dat_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1753.920 2500.000 1754.480 ;
    END
  END dat_in[27]
  PIN dat_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1837.920 2500.000 1838.480 ;
    END
  END dat_in[28]
  PIN dat_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1794.240 2500.000 1794.800 ;
    END
  END dat_in[29]
  PIN dat_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2439.360 2500.000 2439.920 ;
    END
  END dat_in[2]
  PIN dat_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1777.440 2500.000 1778.000 ;
    END
  END dat_in[30]
  PIN dat_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1911.840 2500.000 1912.400 ;
    END
  END dat_in[31]
  PIN dat_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2439.360 4.000 2439.920 ;
    END
  END dat_in[32]
  PIN dat_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2432.640 4.000 2433.200 ;
    END
  END dat_in[33]
  PIN dat_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2429.280 4.000 2429.840 ;
    END
  END dat_in[34]
  PIN dat_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2456.160 4.000 2456.720 ;
    END
  END dat_in[35]
  PIN dat_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2204.160 4.000 2204.720 ;
    END
  END dat_in[36]
  PIN dat_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2200.800 4.000 2201.360 ;
    END
  END dat_in[37]
  PIN dat_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2180.640 4.000 2181.200 ;
    END
  END dat_in[38]
  PIN dat_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2184.000 4.000 2184.560 ;
    END
  END dat_in[39]
  PIN dat_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2436.000 2500.000 2436.560 ;
    END
  END dat_in[3]
  PIN dat_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1629.600 4.000 1630.160 ;
    END
  END dat_in[40]
  PIN dat_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1599.360 4.000 1599.920 ;
    END
  END dat_in[41]
  PIN dat_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1579.200 4.000 1579.760 ;
    END
  END dat_in[42]
  PIN dat_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1585.920 4.000 1586.480 ;
    END
  END dat_in[43]
  PIN dat_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1716.960 4.000 1717.520 ;
    END
  END dat_in[44]
  PIN dat_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1686.720 4.000 1687.280 ;
    END
  END dat_in[45]
  PIN dat_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1700.160 4.000 1700.720 ;
    END
  END dat_in[46]
  PIN dat_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1683.360 4.000 1683.920 ;
    END
  END dat_in[47]
  PIN dat_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2315.040 4.000 2315.600 ;
    END
  END dat_in[48]
  PIN dat_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2378.880 4.000 2379.440 ;
    END
  END dat_in[49]
  PIN dat_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2200.800 2500.000 2201.360 ;
    END
  END dat_in[4]
  PIN dat_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2392.320 4.000 2392.880 ;
    END
  END dat_in[50]
  PIN dat_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2348.640 4.000 2349.200 ;
    END
  END dat_in[51]
  PIN dat_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2106.720 4.000 2107.280 ;
    END
  END dat_in[52]
  PIN dat_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2093.280 4.000 2093.840 ;
    END
  END dat_in[53]
  PIN dat_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2116.800 4.000 2117.360 ;
    END
  END dat_in[54]
  PIN dat_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2103.360 4.000 2103.920 ;
    END
  END dat_in[55]
  PIN dat_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1780.800 4.000 1781.360 ;
    END
  END dat_in[56]
  PIN dat_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1770.720 4.000 1771.280 ;
    END
  END dat_in[57]
  PIN dat_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1764.000 4.000 1764.560 ;
    END
  END dat_in[58]
  PIN dat_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1784.160 4.000 1784.720 ;
    END
  END dat_in[59]
  PIN dat_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2177.280 2500.000 2177.840 ;
    END
  END dat_in[5]
  PIN dat_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1787.520 4.000 1788.080 ;
    END
  END dat_in[60]
  PIN dat_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1790.880 4.000 1791.440 ;
    END
  END dat_in[61]
  PIN dat_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1807.680 4.000 1808.240 ;
    END
  END dat_in[62]
  PIN dat_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1804.320 4.000 1804.880 ;
    END
  END dat_in[63]
  PIN dat_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2167.200 2500.000 2167.760 ;
    END
  END dat_in[6]
  PIN dat_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2157.120 2500.000 2157.680 ;
    END
  END dat_in[7]
  PIN dat_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1535.520 2500.000 1536.080 ;
    END
  END dat_in[8]
  PIN dat_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1538.880 2500.000 1539.440 ;
    END
  END dat_in[9]
  PIN dat_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2251.200 2500.000 2251.760 ;
    END
  END dat_out[0]
  PIN dat_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1690.080 2500.000 1690.640 ;
    END
  END dat_out[10]
  PIN dat_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1696.800 2500.000 1697.360 ;
    END
  END dat_out[11]
  PIN dat_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1693.440 2500.000 1694.000 ;
    END
  END dat_out[12]
  PIN dat_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1703.520 2500.000 1704.080 ;
    END
  END dat_out[13]
  PIN dat_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1700.160 2500.000 1700.720 ;
    END
  END dat_out[14]
  PIN dat_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1770.720 2500.000 1771.280 ;
    END
  END dat_out[15]
  PIN dat_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2261.280 4.000 2261.840 ;
    END
  END dat_out[16]
  PIN dat_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2294.880 4.000 2295.440 ;
    END
  END dat_out[17]
  PIN dat_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2298.240 4.000 2298.800 ;
    END
  END dat_out[18]
  PIN dat_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2291.520 4.000 2292.080 ;
    END
  END dat_out[19]
  PIN dat_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2375.520 2500.000 2376.080 ;
    END
  END dat_out[1]
  PIN dat_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2140.320 4.000 2140.880 ;
    END
  END dat_out[20]
  PIN dat_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2110.080 4.000 2110.640 ;
    END
  END dat_out[21]
  PIN dat_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2096.640 4.000 2097.200 ;
    END
  END dat_out[22]
  PIN dat_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2069.760 4.000 2070.320 ;
    END
  END dat_out[23]
  PIN dat_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1851.360 2500.000 1851.920 ;
    END
  END dat_out[24]
  PIN dat_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1817.760 4.000 1818.320 ;
    END
  END dat_out[25]
  PIN dat_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1848.000 2500.000 1848.560 ;
    END
  END dat_out[26]
  PIN dat_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1811.040 4.000 1811.600 ;
    END
  END dat_out[27]
  PIN dat_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1881.600 2500.000 1882.160 ;
    END
  END dat_out[28]
  PIN dat_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1895.040 4.000 1895.600 ;
    END
  END dat_out[29]
  PIN dat_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2402.400 2500.000 2402.960 ;
    END
  END dat_out[2]
  PIN dat_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1911.840 4.000 1912.400 ;
    END
  END dat_out[30]
  PIN dat_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1925.280 4.000 1925.840 ;
    END
  END dat_out[31]
  PIN dat_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2257.920 2500.000 2258.480 ;
    END
  END dat_out[32]
  PIN dat_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2395.680 2500.000 2396.240 ;
    END
  END dat_out[33]
  PIN dat_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2449.440 2500.000 2450.000 ;
    END
  END dat_out[34]
  PIN dat_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2446.080 2500.000 2446.640 ;
    END
  END dat_out[35]
  PIN dat_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2244.480 2500.000 2245.040 ;
    END
  END dat_out[36]
  PIN dat_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2036.160 2500.000 2036.720 ;
    END
  END dat_out[37]
  PIN dat_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2029.440 2500.000 2030.000 ;
    END
  END dat_out[38]
  PIN dat_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2019.360 2500.000 2019.920 ;
    END
  END dat_out[39]
  PIN dat_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2399.040 2500.000 2399.600 ;
    END
  END dat_out[3]
  PIN dat_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1955.520 2500.000 1956.080 ;
    END
  END dat_out[40]
  PIN dat_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1928.640 2500.000 1929.200 ;
    END
  END dat_out[41]
  PIN dat_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1915.200 2500.000 1915.760 ;
    END
  END dat_out[42]
  PIN dat_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1921.920 2500.000 1922.480 ;
    END
  END dat_out[43]
  PIN dat_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1932.000 2500.000 1932.560 ;
    END
  END dat_out[44]
  PIN dat_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1945.440 2500.000 1946.000 ;
    END
  END dat_out[45]
  PIN dat_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1958.880 2500.000 1959.440 ;
    END
  END dat_out[46]
  PIN dat_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 1962.240 2500.000 1962.800 ;
    END
  END dat_out[47]
  PIN dat_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2405.760 4.000 2406.320 ;
    END
  END dat_out[48]
  PIN dat_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2382.240 4.000 2382.800 ;
    END
  END dat_out[49]
  PIN dat_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2241.120 2500.000 2241.680 ;
    END
  END dat_out[4]
  PIN dat_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2415.840 4.000 2416.400 ;
    END
  END dat_out[50]
  PIN dat_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2399.040 4.000 2399.600 ;
    END
  END dat_out[51]
  PIN dat_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2157.120 4.000 2157.680 ;
    END
  END dat_out[52]
  PIN dat_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2100.000 4.000 2100.560 ;
    END
  END dat_out[53]
  PIN dat_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2163.840 4.000 2164.400 ;
    END
  END dat_out[54]
  PIN dat_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2113.440 4.000 2114.000 ;
    END
  END dat_out[55]
  PIN dat_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1814.400 4.000 1814.960 ;
    END
  END dat_out[56]
  PIN dat_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1797.600 4.000 1798.160 ;
    END
  END dat_out[57]
  PIN dat_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1800.960 4.000 1801.520 ;
    END
  END dat_out[58]
  PIN dat_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1794.240 4.000 1794.800 ;
    END
  END dat_out[59]
  PIN dat_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2052.960 2500.000 2053.520 ;
    END
  END dat_out[5]
  PIN dat_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1774.080 4.000 1774.640 ;
    END
  END dat_out[60]
  PIN dat_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1841.280 4.000 1841.840 ;
    END
  END dat_out[61]
  PIN dat_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1834.560 4.000 1835.120 ;
    END
  END dat_out[62]
  PIN dat_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1844.640 4.000 1845.200 ;
    END
  END dat_out[63]
  PIN dat_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2042.880 2500.000 2043.440 ;
    END
  END dat_out[6]
  PIN dat_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2022.720 2500.000 2023.280 ;
    END
  END dat_out[7]
  PIN dat_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 2496.000 2016.000 2500.000 2016.560 ;
    END
  END dat_out[8]
  PIN dat_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1690.080 4.000 1690.640 ;
    END
  END dat_out[9]
  PIN mat_idx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1962.240 4.000 1962.800 ;
    END
  END mat_idx[0]
  PIN mat_idx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1958.880 4.000 1959.440 ;
    END
  END mat_idx[1]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 3983.020 ;
    END
  END vdd
  PIN vector_idx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2022.720 4.000 2023.280 ;
    END
  END vector_idx[0]
  PIN vector_idx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2016.000 4.000 2016.560 ;
    END
  END vector_idx[1]
  PIN vector_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2019.360 4.000 2019.920 ;
    END
  END vector_type[0]
  PIN vector_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2012.640 4.000 2013.200 ;
    END
  END vector_type[1]
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 3983.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 3983.020 ;
    END
  END vss
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1979.040 4.000 1979.600 ;
    END
  END we
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2493.120 3983.020 ;
      LAYER Metal2 ;
        RECT 8.540 15.490 2491.860 3982.910 ;
      LAYER Metal3 ;
        RECT 4.000 2520.860 2496.000 3982.860 ;
        RECT 4.300 2519.700 2496.000 2520.860 ;
        RECT 4.000 2457.020 2496.000 2519.700 ;
        RECT 4.300 2455.860 2495.700 2457.020 ;
        RECT 4.000 2450.300 2496.000 2455.860 ;
        RECT 4.000 2449.140 2495.700 2450.300 ;
        RECT 4.000 2446.940 2496.000 2449.140 ;
        RECT 4.000 2445.780 2495.700 2446.940 ;
        RECT 4.000 2443.580 2496.000 2445.780 ;
        RECT 4.000 2442.420 2495.700 2443.580 ;
        RECT 4.000 2440.220 2496.000 2442.420 ;
        RECT 4.300 2439.060 2495.700 2440.220 ;
        RECT 4.000 2436.860 2496.000 2439.060 ;
        RECT 4.000 2435.700 2495.700 2436.860 ;
        RECT 4.000 2433.500 2496.000 2435.700 ;
        RECT 4.300 2432.340 2496.000 2433.500 ;
        RECT 4.000 2430.140 2496.000 2432.340 ;
        RECT 4.300 2428.980 2496.000 2430.140 ;
        RECT 4.000 2416.700 2496.000 2428.980 ;
        RECT 4.300 2415.540 2496.000 2416.700 ;
        RECT 4.000 2406.620 2496.000 2415.540 ;
        RECT 4.300 2405.460 2496.000 2406.620 ;
        RECT 4.000 2403.260 2496.000 2405.460 ;
        RECT 4.000 2402.100 2495.700 2403.260 ;
        RECT 4.000 2399.900 2496.000 2402.100 ;
        RECT 4.300 2398.740 2495.700 2399.900 ;
        RECT 4.000 2396.540 2496.000 2398.740 ;
        RECT 4.000 2395.380 2495.700 2396.540 ;
        RECT 4.000 2393.180 2496.000 2395.380 ;
        RECT 4.300 2392.020 2496.000 2393.180 ;
        RECT 4.000 2383.100 2496.000 2392.020 ;
        RECT 4.300 2381.940 2496.000 2383.100 ;
        RECT 4.000 2379.740 2496.000 2381.940 ;
        RECT 4.300 2378.580 2496.000 2379.740 ;
        RECT 4.000 2376.380 2496.000 2378.580 ;
        RECT 4.000 2375.220 2495.700 2376.380 ;
        RECT 4.000 2352.860 2496.000 2375.220 ;
        RECT 4.300 2351.700 2496.000 2352.860 ;
        RECT 4.000 2349.500 2496.000 2351.700 ;
        RECT 4.300 2348.340 2496.000 2349.500 ;
        RECT 4.000 2315.900 2496.000 2348.340 ;
        RECT 4.300 2314.740 2496.000 2315.900 ;
        RECT 4.000 2309.180 2496.000 2314.740 ;
        RECT 4.000 2308.020 2495.700 2309.180 ;
        RECT 4.000 2305.820 2496.000 2308.020 ;
        RECT 4.000 2304.660 2495.700 2305.820 ;
        RECT 4.000 2299.100 2496.000 2304.660 ;
        RECT 4.300 2297.940 2496.000 2299.100 ;
        RECT 4.000 2295.740 2496.000 2297.940 ;
        RECT 4.300 2294.580 2496.000 2295.740 ;
        RECT 4.000 2292.380 2496.000 2294.580 ;
        RECT 4.300 2291.220 2496.000 2292.380 ;
        RECT 4.000 2289.020 2496.000 2291.220 ;
        RECT 4.300 2287.860 2496.000 2289.020 ;
        RECT 4.000 2262.140 2496.000 2287.860 ;
        RECT 4.300 2260.980 2496.000 2262.140 ;
        RECT 4.000 2258.780 2496.000 2260.980 ;
        RECT 4.000 2257.620 2495.700 2258.780 ;
        RECT 4.000 2252.060 2496.000 2257.620 ;
        RECT 4.000 2250.900 2495.700 2252.060 ;
        RECT 4.000 2245.340 2496.000 2250.900 ;
        RECT 4.000 2244.180 2495.700 2245.340 ;
        RECT 4.000 2241.980 2496.000 2244.180 ;
        RECT 4.000 2240.820 2495.700 2241.980 ;
        RECT 4.000 2205.020 2496.000 2240.820 ;
        RECT 4.300 2203.860 2496.000 2205.020 ;
        RECT 4.000 2201.660 2496.000 2203.860 ;
        RECT 4.300 2200.500 2495.700 2201.660 ;
        RECT 4.000 2184.860 2496.000 2200.500 ;
        RECT 4.300 2183.700 2496.000 2184.860 ;
        RECT 4.000 2181.500 2496.000 2183.700 ;
        RECT 4.300 2180.340 2496.000 2181.500 ;
        RECT 4.000 2178.140 2496.000 2180.340 ;
        RECT 4.000 2176.980 2495.700 2178.140 ;
        RECT 4.000 2168.060 2496.000 2176.980 ;
        RECT 4.000 2166.900 2495.700 2168.060 ;
        RECT 4.000 2164.700 2496.000 2166.900 ;
        RECT 4.300 2163.540 2496.000 2164.700 ;
        RECT 4.000 2157.980 2496.000 2163.540 ;
        RECT 4.300 2156.820 2495.700 2157.980 ;
        RECT 4.000 2141.180 2496.000 2156.820 ;
        RECT 4.300 2140.020 2496.000 2141.180 ;
        RECT 4.000 2117.660 2496.000 2140.020 ;
        RECT 4.300 2116.500 2495.700 2117.660 ;
        RECT 4.000 2114.300 2496.000 2116.500 ;
        RECT 4.300 2113.140 2496.000 2114.300 ;
        RECT 4.000 2110.940 2496.000 2113.140 ;
        RECT 4.300 2109.780 2496.000 2110.940 ;
        RECT 4.000 2107.580 2496.000 2109.780 ;
        RECT 4.300 2106.420 2496.000 2107.580 ;
        RECT 4.000 2104.220 2496.000 2106.420 ;
        RECT 4.300 2103.060 2495.700 2104.220 ;
        RECT 4.000 2100.860 2496.000 2103.060 ;
        RECT 4.300 2099.700 2496.000 2100.860 ;
        RECT 4.000 2097.500 2496.000 2099.700 ;
        RECT 4.300 2096.340 2496.000 2097.500 ;
        RECT 4.000 2094.140 2496.000 2096.340 ;
        RECT 4.300 2092.980 2496.000 2094.140 ;
        RECT 4.000 2073.980 2496.000 2092.980 ;
        RECT 4.000 2072.820 2495.700 2073.980 ;
        RECT 4.000 2070.620 2496.000 2072.820 ;
        RECT 4.300 2069.460 2496.000 2070.620 ;
        RECT 4.000 2057.180 2496.000 2069.460 ;
        RECT 4.000 2056.020 2495.700 2057.180 ;
        RECT 4.000 2053.820 2496.000 2056.020 ;
        RECT 4.000 2052.660 2495.700 2053.820 ;
        RECT 4.000 2043.740 2496.000 2052.660 ;
        RECT 4.000 2042.580 2495.700 2043.740 ;
        RECT 4.000 2037.020 2496.000 2042.580 ;
        RECT 4.000 2035.860 2495.700 2037.020 ;
        RECT 4.000 2030.300 2496.000 2035.860 ;
        RECT 4.000 2029.140 2495.700 2030.300 ;
        RECT 4.000 2023.580 2496.000 2029.140 ;
        RECT 4.300 2022.420 2495.700 2023.580 ;
        RECT 4.000 2020.220 2496.000 2022.420 ;
        RECT 4.300 2019.060 2495.700 2020.220 ;
        RECT 4.000 2016.860 2496.000 2019.060 ;
        RECT 4.300 2015.700 2495.700 2016.860 ;
        RECT 4.000 2013.500 2496.000 2015.700 ;
        RECT 4.300 2012.340 2496.000 2013.500 ;
        RECT 4.000 1979.900 2496.000 2012.340 ;
        RECT 4.300 1978.740 2496.000 1979.900 ;
        RECT 4.000 1976.540 2496.000 1978.740 ;
        RECT 4.300 1975.380 2496.000 1976.540 ;
        RECT 4.000 1963.100 2496.000 1975.380 ;
        RECT 4.300 1961.940 2495.700 1963.100 ;
        RECT 4.000 1959.740 2496.000 1961.940 ;
        RECT 4.300 1958.580 2495.700 1959.740 ;
        RECT 4.000 1956.380 2496.000 1958.580 ;
        RECT 4.000 1955.220 2495.700 1956.380 ;
        RECT 4.000 1953.020 2496.000 1955.220 ;
        RECT 4.300 1951.860 2496.000 1953.020 ;
        RECT 4.000 1946.300 2496.000 1951.860 ;
        RECT 4.000 1945.140 2495.700 1946.300 ;
        RECT 4.000 1932.860 2496.000 1945.140 ;
        RECT 4.000 1931.700 2495.700 1932.860 ;
        RECT 4.000 1929.500 2496.000 1931.700 ;
        RECT 4.000 1928.340 2495.700 1929.500 ;
        RECT 4.000 1926.140 2496.000 1928.340 ;
        RECT 4.300 1924.980 2496.000 1926.140 ;
        RECT 4.000 1922.780 2496.000 1924.980 ;
        RECT 4.000 1921.620 2495.700 1922.780 ;
        RECT 4.000 1916.060 2496.000 1921.620 ;
        RECT 4.000 1914.900 2495.700 1916.060 ;
        RECT 4.000 1912.700 2496.000 1914.900 ;
        RECT 4.300 1911.540 2495.700 1912.700 ;
        RECT 4.000 1895.900 2496.000 1911.540 ;
        RECT 4.300 1894.740 2496.000 1895.900 ;
        RECT 4.000 1882.460 2496.000 1894.740 ;
        RECT 4.000 1881.300 2495.700 1882.460 ;
        RECT 4.000 1852.220 2496.000 1881.300 ;
        RECT 4.000 1851.060 2495.700 1852.220 ;
        RECT 4.000 1848.860 2496.000 1851.060 ;
        RECT 4.000 1847.700 2495.700 1848.860 ;
        RECT 4.000 1845.500 2496.000 1847.700 ;
        RECT 4.300 1844.340 2496.000 1845.500 ;
        RECT 4.000 1842.140 2496.000 1844.340 ;
        RECT 4.300 1840.980 2496.000 1842.140 ;
        RECT 4.000 1838.780 2496.000 1840.980 ;
        RECT 4.000 1837.620 2495.700 1838.780 ;
        RECT 4.000 1835.420 2496.000 1837.620 ;
        RECT 4.300 1834.260 2496.000 1835.420 ;
        RECT 4.000 1818.620 2496.000 1834.260 ;
        RECT 4.300 1817.460 2495.700 1818.620 ;
        RECT 4.000 1815.260 2496.000 1817.460 ;
        RECT 4.300 1814.100 2496.000 1815.260 ;
        RECT 4.000 1811.900 2496.000 1814.100 ;
        RECT 4.300 1810.740 2496.000 1811.900 ;
        RECT 4.000 1808.540 2496.000 1810.740 ;
        RECT 4.300 1807.380 2496.000 1808.540 ;
        RECT 4.000 1805.180 2496.000 1807.380 ;
        RECT 4.300 1804.020 2496.000 1805.180 ;
        RECT 4.000 1801.820 2496.000 1804.020 ;
        RECT 4.300 1800.660 2496.000 1801.820 ;
        RECT 4.000 1798.460 2496.000 1800.660 ;
        RECT 4.300 1797.300 2496.000 1798.460 ;
        RECT 4.000 1795.100 2496.000 1797.300 ;
        RECT 4.300 1793.940 2495.700 1795.100 ;
        RECT 4.000 1791.740 2496.000 1793.940 ;
        RECT 4.300 1790.580 2496.000 1791.740 ;
        RECT 4.000 1788.380 2496.000 1790.580 ;
        RECT 4.300 1787.220 2496.000 1788.380 ;
        RECT 4.000 1785.020 2496.000 1787.220 ;
        RECT 4.300 1783.860 2496.000 1785.020 ;
        RECT 4.000 1781.660 2496.000 1783.860 ;
        RECT 4.300 1780.500 2496.000 1781.660 ;
        RECT 4.000 1778.300 2496.000 1780.500 ;
        RECT 4.000 1777.140 2495.700 1778.300 ;
        RECT 4.000 1774.940 2496.000 1777.140 ;
        RECT 4.300 1773.780 2496.000 1774.940 ;
        RECT 4.000 1771.580 2496.000 1773.780 ;
        RECT 4.300 1770.420 2495.700 1771.580 ;
        RECT 4.000 1764.860 2496.000 1770.420 ;
        RECT 4.300 1763.700 2496.000 1764.860 ;
        RECT 4.000 1761.500 2496.000 1763.700 ;
        RECT 4.000 1760.340 2495.700 1761.500 ;
        RECT 4.000 1758.140 2496.000 1760.340 ;
        RECT 4.000 1756.980 2495.700 1758.140 ;
        RECT 4.000 1754.780 2496.000 1756.980 ;
        RECT 4.000 1753.620 2495.700 1754.780 ;
        RECT 4.000 1717.820 2496.000 1753.620 ;
        RECT 4.300 1716.660 2496.000 1717.820 ;
        RECT 4.000 1704.380 2496.000 1716.660 ;
        RECT 4.000 1703.220 2495.700 1704.380 ;
        RECT 4.000 1701.020 2496.000 1703.220 ;
        RECT 4.300 1699.860 2495.700 1701.020 ;
        RECT 4.000 1697.660 2496.000 1699.860 ;
        RECT 4.000 1696.500 2495.700 1697.660 ;
        RECT 4.000 1694.300 2496.000 1696.500 ;
        RECT 4.000 1693.140 2495.700 1694.300 ;
        RECT 4.000 1690.940 2496.000 1693.140 ;
        RECT 4.300 1689.780 2495.700 1690.940 ;
        RECT 4.000 1687.580 2496.000 1689.780 ;
        RECT 4.300 1686.420 2496.000 1687.580 ;
        RECT 4.000 1684.220 2496.000 1686.420 ;
        RECT 4.300 1683.060 2496.000 1684.220 ;
        RECT 4.000 1633.820 2496.000 1683.060 ;
        RECT 4.000 1632.660 2495.700 1633.820 ;
        RECT 4.000 1630.460 2496.000 1632.660 ;
        RECT 4.300 1629.300 2495.700 1630.460 ;
        RECT 4.000 1627.100 2496.000 1629.300 ;
        RECT 4.000 1625.940 2495.700 1627.100 ;
        RECT 4.000 1620.380 2496.000 1625.940 ;
        RECT 4.000 1619.220 2495.700 1620.380 ;
        RECT 4.000 1600.220 2496.000 1619.220 ;
        RECT 4.300 1599.060 2496.000 1600.220 ;
        RECT 4.000 1586.780 2496.000 1599.060 ;
        RECT 4.300 1585.620 2496.000 1586.780 ;
        RECT 4.000 1580.060 2496.000 1585.620 ;
        RECT 4.300 1578.900 2496.000 1580.060 ;
        RECT 4.000 1576.700 2496.000 1578.900 ;
        RECT 4.000 1575.540 2495.700 1576.700 ;
        RECT 4.000 1553.180 2496.000 1575.540 ;
        RECT 4.000 1552.020 2495.700 1553.180 ;
        RECT 4.000 1539.740 2496.000 1552.020 ;
        RECT 4.000 1538.580 2495.700 1539.740 ;
        RECT 4.000 1536.380 2496.000 1538.580 ;
        RECT 4.000 1535.220 2495.700 1536.380 ;
        RECT 4.000 15.540 2496.000 1535.220 ;
      LAYER Metal4 ;
        RECT 1009.260 1507.610 1020.340 2521.590 ;
        RECT 1022.540 1507.610 1097.140 2521.590 ;
        RECT 1099.340 1507.610 1173.940 2521.590 ;
        RECT 1176.140 1507.610 1250.740 2521.590 ;
        RECT 1252.940 1507.610 1327.540 2521.590 ;
        RECT 1329.740 1507.610 1404.340 2521.590 ;
        RECT 1406.540 1507.610 1481.140 2521.590 ;
        RECT 1483.340 1507.610 1492.820 2521.590 ;
  END
END gpu_core
END LIBRARY

