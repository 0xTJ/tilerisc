VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180_ram_128x8_wrapper
  CLASS BLOCK ;
  FOREIGN gf180_ram_128x8_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 444.860 BY 279.880 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.720 275.880 265.280 279.880 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.220 275.880 273.780 279.880 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.720 275.880 282.280 279.880 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.720 275.880 155.280 279.880 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.720 275.880 160.280 279.880 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.720 275.880 164.280 279.880 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.720 275.880 167.280 279.880 ;
    END
  END A[6]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.220 275.880 184.780 279.880 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.220 275.880 296.780 279.880 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 275.880 427.280 279.880 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.720 275.880 375.280 279.880 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 368.720 275.880 369.280 279.880 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.720 275.880 317.280 279.880 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.720 275.880 129.280 279.880 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.220 275.880 77.780 279.880 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.720 275.880 71.280 279.880 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.720 275.880 19.280 279.880 ;
    END
  END D[7]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.840 275.880 233.400 279.880 ;
    END
  END GWEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 419.220 275.880 419.780 279.880 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.220 275.880 378.780 279.880 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.220 275.880 365.780 279.880 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.720 275.880 325.280 279.880 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.220 275.880 121.780 279.880 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.220 275.880 80.780 279.880 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.220 275.880 67.780 279.880 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.720 275.880 27.280 279.880 ;
    END
  END Q[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 5.220 15.680 8.220 262.640 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 428.630 15.680 431.630 262.640 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 9.220 15.680 12.220 262.640 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 432.630 15.680 435.630 262.640 ;
    END
  END VSS
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.220 275.880 423.780 279.880 ;
    END
  END WEN[0]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.720 275.880 373.280 279.880 ;
    END
  END WEN[1]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 275.880 371.280 279.880 ;
    END
  END WEN[2]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.720 275.880 319.280 279.880 ;
    END
  END WEN[3]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.220 275.880 125.780 279.880 ;
    END
  END WEN[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.970 275.880 75.530 279.880 ;
    END
  END WEN[5]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.720 275.880 73.280 279.880 ;
    END
  END WEN[6]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.220 275.880 22.780 279.880 ;
    END
  END WEN[7]
  OBS
      LAYER Metal1 ;
        RECT 5.000 5.000 436.860 273.880 ;
      LAYER Metal2 ;
        RECT 5.000 275.580 18.420 276.360 ;
        RECT 19.580 275.580 21.920 276.360 ;
        RECT 23.080 275.580 26.420 276.360 ;
        RECT 27.580 275.580 66.920 276.360 ;
        RECT 68.080 275.580 70.420 276.360 ;
        RECT 71.580 275.580 72.420 276.360 ;
        RECT 73.580 275.580 74.670 276.360 ;
        RECT 75.830 275.580 76.920 276.360 ;
        RECT 78.080 275.580 79.920 276.360 ;
        RECT 81.080 275.580 120.920 276.360 ;
        RECT 122.080 275.580 124.920 276.360 ;
        RECT 126.080 275.580 128.420 276.360 ;
        RECT 129.580 275.580 154.420 276.360 ;
        RECT 155.580 275.580 159.420 276.360 ;
        RECT 160.580 275.580 163.420 276.360 ;
        RECT 164.580 275.580 166.420 276.360 ;
        RECT 167.580 275.580 183.920 276.360 ;
        RECT 185.080 275.580 232.540 276.360 ;
        RECT 233.700 275.580 264.420 276.360 ;
        RECT 265.580 275.580 272.920 276.360 ;
        RECT 274.080 275.580 281.420 276.360 ;
        RECT 282.580 275.580 295.920 276.360 ;
        RECT 297.080 275.580 316.420 276.360 ;
        RECT 317.580 275.580 318.420 276.360 ;
        RECT 319.580 275.580 324.420 276.360 ;
        RECT 325.580 275.580 364.920 276.360 ;
        RECT 366.080 275.580 368.420 276.360 ;
        RECT 369.580 275.580 370.420 276.360 ;
        RECT 371.580 275.580 372.420 276.360 ;
        RECT 373.580 275.580 374.420 276.360 ;
        RECT 375.580 275.580 377.920 276.360 ;
        RECT 379.080 275.580 418.920 276.360 ;
        RECT 420.080 275.580 422.920 276.360 ;
        RECT 424.080 275.580 426.420 276.360 ;
        RECT 427.580 275.580 436.860 276.360 ;
        RECT 5.000 5.000 436.860 275.580 ;
      LAYER Metal3 ;
        RECT 5.000 5.000 436.860 273.880 ;
  END
END gf180_ram_128x8_wrapper
END LIBRARY

