magic
tech gf180mcuD
magscale 1 10
timestamp 1700157466
<< metal2 >>
rect 3744 69576 3856 70376
rect 4444 69608 4556 70376
rect 5344 69608 5456 70376
rect 4444 69576 4564 69608
rect 5344 69576 5460 69608
rect 13444 69576 13556 70376
rect 14144 69608 14256 70376
rect 14140 69576 14256 69608
rect 14544 69576 14656 70376
rect 14994 69576 15106 70376
rect 15444 69576 15556 70376
rect 16044 69576 16156 70376
rect 24244 69576 24356 70376
rect 25044 69576 25156 70376
rect 25744 69576 25856 70376
rect 30944 69608 31056 70376
rect 30940 69576 31056 69608
rect 31944 69576 32056 70376
rect 32744 69576 32856 70376
rect 33344 69608 33456 70376
rect 33344 69576 33460 69608
rect 36844 69576 36956 70376
rect 46568 69576 46680 70376
rect 52944 69608 53056 70376
rect 52944 69576 53060 69608
rect 54644 69576 54756 70376
rect 56344 69576 56456 70376
rect 57444 69576 57556 70376
rect 59244 69576 59356 70376
rect 63344 69576 63456 70376
rect 63744 69576 63856 70376
rect 64944 69576 65056 70376
rect 73044 69576 73156 70376
rect 73744 69576 73856 70376
rect 74144 69576 74256 70376
rect 74544 69576 74656 70376
rect 74944 69576 75056 70376
rect 75644 69576 75756 70376
rect 83844 69576 83956 70376
rect 84644 69576 84756 70376
rect 85344 69576 85456 70376
rect 3780 69048 3836 69576
rect 4508 69048 4564 69576
rect 5404 69048 5460 69576
rect 13468 69048 13524 69576
rect 14140 69048 14196 69576
rect 14588 69048 14644 69576
rect 15036 69048 15092 69576
rect 15484 69048 15540 69576
rect 16044 69048 16100 69576
rect 24276 69048 24332 69576
rect 25060 69048 25116 69576
rect 25788 69048 25844 69576
rect 30940 69048 30996 69576
rect 31948 69300 32004 69576
rect 31948 69244 32116 69300
rect 32060 69048 32116 69244
rect 32788 69048 32844 69576
rect 33404 69048 33460 69576
rect 36876 69048 36932 69576
rect 46620 69048 46676 69576
rect 53004 69048 53060 69576
rect 54684 69048 54740 69576
rect 56364 69048 56420 69576
rect 57484 69048 57540 69576
rect 59276 69048 59332 69576
rect 63364 69048 63420 69576
rect 63756 69048 63812 69576
rect 64988 69048 65044 69576
rect 73052 69048 73108 69576
rect 73780 69048 73836 69576
rect 74172 69048 74228 69576
rect 74564 69048 74620 69576
rect 74956 69048 75012 69576
rect 75684 69048 75740 69576
rect 83860 69048 83916 69576
rect 84700 69048 84756 69576
rect 85372 69048 85428 69576
<< metal3 >>
rect 1906 66571 2382 66640
rect 1906 66515 1930 66571
rect 1986 66515 2054 66571
rect 2110 66515 2178 66571
rect 2234 66515 2302 66571
rect 2358 66515 2382 66571
rect 1906 66447 2382 66515
rect 1906 66391 1930 66447
rect 1986 66391 2054 66447
rect 2110 66391 2178 66447
rect 2234 66391 2302 66447
rect 2358 66391 2382 66447
rect 1906 66322 2382 66391
rect 86526 66608 86630 66640
rect 86526 66552 86550 66608
rect 86606 66552 86630 66608
rect 86526 66484 86630 66552
rect 86526 66428 86550 66484
rect 86606 66428 86630 66484
rect 86526 66360 86630 66428
rect 86526 66304 86550 66360
rect 86606 66304 86630 66360
rect 86526 66236 86630 66304
rect 86526 66180 86550 66236
rect 86606 66180 86630 66236
rect 86526 66148 86630 66180
rect 86650 66608 87126 66640
rect 86650 66552 86674 66608
rect 86730 66552 86798 66608
rect 86854 66552 86922 66608
rect 86978 66552 87046 66608
rect 87102 66552 87126 66608
rect 86650 66484 87126 66552
rect 86650 66428 86674 66484
rect 86730 66428 86798 66484
rect 86854 66428 86922 66484
rect 86978 66428 87046 66484
rect 87102 66428 87126 66484
rect 86650 66360 87126 66428
rect 86650 66304 86674 66360
rect 86730 66304 86798 66360
rect 86854 66304 86922 66360
rect 86978 66304 87046 66360
rect 87102 66304 87126 66360
rect 86650 66236 87126 66304
rect 86650 66180 86674 66236
rect 86730 66180 86798 66236
rect 86854 66180 86922 66236
rect 86978 66180 87046 66236
rect 87102 66180 87126 66236
rect 86650 66148 87126 66180
rect 86526 66112 86630 66144
rect 86526 66056 86550 66112
rect 86606 66056 86630 66112
rect 86526 65988 86630 66056
rect 86526 65932 86550 65988
rect 86606 65932 86630 65988
rect 86526 65864 86630 65932
rect 86526 65808 86550 65864
rect 86606 65808 86630 65864
rect 1906 65732 2382 65756
rect 1906 65676 1930 65732
rect 1986 65676 2054 65732
rect 2110 65676 2178 65732
rect 2234 65676 2302 65732
rect 2358 65676 2382 65732
rect 1906 65608 2382 65676
rect 86526 65740 86630 65808
rect 86526 65684 86550 65740
rect 86606 65684 86630 65740
rect 86526 65652 86630 65684
rect 86650 66112 87126 66144
rect 86650 66056 86674 66112
rect 86730 66056 86798 66112
rect 86854 66056 86922 66112
rect 86978 66056 87046 66112
rect 87102 66056 87126 66112
rect 86650 65988 87126 66056
rect 86650 65932 86674 65988
rect 86730 65932 86798 65988
rect 86854 65932 86922 65988
rect 86978 65932 87046 65988
rect 87102 65932 87126 65988
rect 86650 65864 87126 65932
rect 86650 65808 86674 65864
rect 86730 65808 86798 65864
rect 86854 65808 86922 65864
rect 86978 65808 87046 65864
rect 87102 65808 87126 65864
rect 86650 65740 87126 65808
rect 86650 65684 86674 65740
rect 86730 65684 86798 65740
rect 86854 65684 86922 65740
rect 86978 65684 87046 65740
rect 87102 65684 87126 65740
rect 86650 65652 87126 65684
rect 1906 65552 1930 65608
rect 1986 65552 2054 65608
rect 2110 65552 2178 65608
rect 2234 65552 2302 65608
rect 2358 65552 2382 65608
rect 1906 65484 2382 65552
rect 1906 65428 1930 65484
rect 1986 65428 2054 65484
rect 2110 65428 2178 65484
rect 2234 65428 2302 65484
rect 2358 65428 2382 65484
rect 1906 65404 2382 65428
rect 86526 65616 86630 65648
rect 86526 65560 86550 65616
rect 86606 65560 86630 65616
rect 86526 65492 86630 65560
rect 86526 65436 86550 65492
rect 86606 65436 86630 65492
rect 86526 65404 86630 65436
rect 86650 65616 87126 65648
rect 86650 65560 86674 65616
rect 86730 65560 86798 65616
rect 86854 65560 86922 65616
rect 86978 65560 87046 65616
rect 87102 65560 87126 65616
rect 86650 65492 87126 65560
rect 86650 65436 86674 65492
rect 86730 65436 86798 65492
rect 86854 65436 86922 65492
rect 86978 65436 87046 65492
rect 87102 65436 87126 65492
rect 86650 65404 87126 65436
rect 1906 63346 2382 63410
rect 1906 63290 1930 63346
rect 1986 63290 2054 63346
rect 2110 63290 2178 63346
rect 2234 63290 2302 63346
rect 2358 63290 2382 63346
rect 1906 63222 2382 63290
rect 1906 63166 1930 63222
rect 1986 63166 2054 63222
rect 2110 63166 2178 63222
rect 2234 63166 2302 63222
rect 2358 63166 2382 63222
rect 1906 63098 2382 63166
rect 1906 63042 1930 63098
rect 1986 63042 2054 63098
rect 2110 63042 2178 63098
rect 2234 63042 2302 63098
rect 2358 63042 2382 63098
rect 1906 62978 2382 63042
rect 86526 63391 86630 63410
rect 86526 63335 86550 63391
rect 86606 63335 86630 63391
rect 86526 63267 86630 63335
rect 86526 63211 86550 63267
rect 86606 63211 86630 63267
rect 86526 63143 86630 63211
rect 86526 63087 86550 63143
rect 86606 63087 86630 63143
rect 86526 63019 86630 63087
rect 86526 62963 86550 63019
rect 86606 62963 86630 63019
rect 86526 62944 86630 62963
rect 86650 63391 87126 63410
rect 86650 63335 86674 63391
rect 86730 63335 86798 63391
rect 86854 63335 86922 63391
rect 86978 63335 87046 63391
rect 87102 63335 87126 63391
rect 86650 63267 87126 63335
rect 86650 63211 86674 63267
rect 86730 63211 86798 63267
rect 86854 63211 86922 63267
rect 86978 63211 87046 63267
rect 87102 63211 87126 63267
rect 86650 63143 87126 63211
rect 86650 63087 86674 63143
rect 86730 63087 86798 63143
rect 86854 63087 86922 63143
rect 86978 63087 87046 63143
rect 87102 63087 87126 63143
rect 86650 63019 87126 63087
rect 86650 62963 86674 63019
rect 86730 62963 86798 63019
rect 86854 62963 86922 63019
rect 86978 62963 87046 63019
rect 87102 62963 87126 63019
rect 86650 62944 87126 62963
rect 86526 62895 86630 62914
rect 86526 62839 86550 62895
rect 86606 62839 86630 62895
rect 86526 62771 86630 62839
rect 86526 62715 86550 62771
rect 86606 62715 86630 62771
rect 86526 62647 86630 62715
rect 86526 62591 86550 62647
rect 86606 62591 86630 62647
rect 86526 62523 86630 62591
rect 86526 62467 86550 62523
rect 86606 62467 86630 62523
rect 86526 62448 86630 62467
rect 86650 62895 87126 62914
rect 86650 62839 86674 62895
rect 86730 62839 86798 62895
rect 86854 62839 86922 62895
rect 86978 62839 87046 62895
rect 87102 62839 87126 62895
rect 86650 62771 87126 62839
rect 86650 62715 86674 62771
rect 86730 62715 86798 62771
rect 86854 62715 86922 62771
rect 86978 62715 87046 62771
rect 87102 62715 87126 62771
rect 86650 62647 87126 62715
rect 86650 62591 86674 62647
rect 86730 62591 86798 62647
rect 86854 62591 86922 62647
rect 86978 62591 87046 62647
rect 87102 62591 87126 62647
rect 86650 62523 87126 62591
rect 86650 62467 86674 62523
rect 86730 62467 86798 62523
rect 86854 62467 86922 62523
rect 86978 62467 87046 62523
rect 87102 62467 87126 62523
rect 86650 62448 87126 62467
rect 86526 62399 86630 62418
rect 86526 62343 86550 62399
rect 86606 62343 86630 62399
rect 86526 62275 86630 62343
rect 86526 62219 86550 62275
rect 86606 62219 86630 62275
rect 86526 62151 86630 62219
rect 1906 62101 2382 62132
rect 1906 62045 1930 62101
rect 1986 62045 2054 62101
rect 2110 62045 2178 62101
rect 2234 62045 2302 62101
rect 2358 62045 2382 62101
rect 1906 61977 2382 62045
rect 1906 61921 1930 61977
rect 1986 61921 2054 61977
rect 2110 61921 2178 61977
rect 2234 61921 2302 61977
rect 2358 61921 2382 61977
rect 86526 62095 86550 62151
rect 86606 62095 86630 62151
rect 86526 62027 86630 62095
rect 86526 61971 86550 62027
rect 86606 61971 86630 62027
rect 86526 61952 86630 61971
rect 86650 62399 87126 62418
rect 86650 62343 86674 62399
rect 86730 62343 86798 62399
rect 86854 62343 86922 62399
rect 86978 62343 87046 62399
rect 87102 62343 87126 62399
rect 86650 62275 87126 62343
rect 86650 62219 86674 62275
rect 86730 62219 86798 62275
rect 86854 62219 86922 62275
rect 86978 62219 87046 62275
rect 87102 62219 87126 62275
rect 86650 62151 87126 62219
rect 86650 62095 86674 62151
rect 86730 62095 86798 62151
rect 86854 62095 86922 62151
rect 86978 62095 87046 62151
rect 87102 62095 87126 62151
rect 86650 62027 87126 62095
rect 86650 61971 86674 62027
rect 86730 61971 86798 62027
rect 86854 61971 86922 62027
rect 86978 61971 87046 62027
rect 87102 61971 87126 62027
rect 86650 61952 87126 61971
rect 1906 61853 2382 61921
rect 1906 61797 1930 61853
rect 1986 61797 2054 61853
rect 2110 61797 2178 61853
rect 2234 61797 2302 61853
rect 2358 61797 2382 61853
rect 1906 61729 2382 61797
rect 1906 61673 1930 61729
rect 1986 61673 2054 61729
rect 2110 61673 2178 61729
rect 2234 61673 2302 61729
rect 2358 61673 2382 61729
rect 1906 61642 2382 61673
rect 86526 61903 86630 61922
rect 86526 61847 86550 61903
rect 86606 61847 86630 61903
rect 86526 61779 86630 61847
rect 86526 61723 86550 61779
rect 86606 61723 86630 61779
rect 86526 61655 86630 61723
rect 86526 61599 86550 61655
rect 86606 61599 86630 61655
rect 86526 61580 86630 61599
rect 86650 61903 87126 61922
rect 86650 61847 86674 61903
rect 86730 61847 86798 61903
rect 86854 61847 86922 61903
rect 86978 61847 87046 61903
rect 87102 61847 87126 61903
rect 86650 61779 87126 61847
rect 86650 61723 86674 61779
rect 86730 61723 86798 61779
rect 86854 61723 86922 61779
rect 86978 61723 87046 61779
rect 87102 61723 87126 61779
rect 86650 61655 87126 61723
rect 86650 61599 86674 61655
rect 86730 61599 86798 61655
rect 86854 61599 86922 61655
rect 86978 61599 87046 61655
rect 87102 61599 87126 61655
rect 86650 61580 87126 61599
rect 85726 60991 85830 61024
rect 85726 60935 85750 60991
rect 85806 60935 85830 60991
rect 85726 60867 85830 60935
rect 85726 60811 85750 60867
rect 85806 60811 85830 60867
rect 85726 60743 85830 60811
rect 85726 60687 85750 60743
rect 85806 60687 85830 60743
rect 85726 60619 85830 60687
rect 85726 60563 85750 60619
rect 85806 60563 85830 60619
rect 85726 60530 85830 60563
rect 85850 60991 86326 61024
rect 85850 60935 85874 60991
rect 85930 60935 85998 60991
rect 86054 60935 86122 60991
rect 86178 60935 86246 60991
rect 86302 60935 86326 60991
rect 85850 60867 86326 60935
rect 85850 60811 85874 60867
rect 85930 60811 85998 60867
rect 86054 60811 86122 60867
rect 86178 60811 86246 60867
rect 86302 60811 86326 60867
rect 85850 60743 86326 60811
rect 85850 60687 85874 60743
rect 85930 60687 85998 60743
rect 86054 60687 86122 60743
rect 86178 60687 86246 60743
rect 86302 60687 86326 60743
rect 85850 60619 86326 60687
rect 85850 60563 85874 60619
rect 85930 60563 85998 60619
rect 86054 60563 86122 60619
rect 86178 60563 86246 60619
rect 86302 60563 86326 60619
rect 85850 60530 86326 60563
rect 85726 60495 85830 60528
rect 85726 60439 85750 60495
rect 85806 60439 85830 60495
rect 85726 60371 85830 60439
rect 85726 60315 85750 60371
rect 85806 60315 85830 60371
rect 85726 60247 85830 60315
rect 85726 60191 85750 60247
rect 85806 60191 85830 60247
rect 85726 60123 85830 60191
rect 85726 60067 85750 60123
rect 85806 60067 85830 60123
rect 85726 60034 85830 60067
rect 85850 60495 86326 60528
rect 85850 60439 85874 60495
rect 85930 60439 85998 60495
rect 86054 60439 86122 60495
rect 86178 60439 86246 60495
rect 86302 60439 86326 60495
rect 85850 60371 86326 60439
rect 85850 60315 85874 60371
rect 85930 60315 85998 60371
rect 86054 60315 86122 60371
rect 86178 60315 86246 60371
rect 86302 60315 86326 60371
rect 85850 60247 86326 60315
rect 85850 60191 85874 60247
rect 85930 60191 85998 60247
rect 86054 60191 86122 60247
rect 86178 60191 86246 60247
rect 86302 60191 86326 60247
rect 85850 60123 86326 60191
rect 85850 60067 85874 60123
rect 85930 60067 85998 60123
rect 86054 60067 86122 60123
rect 86178 60067 86246 60123
rect 86302 60067 86326 60123
rect 85850 60034 86326 60067
rect 85726 59999 85830 60032
rect 85726 59943 85750 59999
rect 85806 59943 85830 59999
rect 85726 59875 85830 59943
rect 85726 59819 85750 59875
rect 85806 59819 85830 59875
rect 85726 59751 85830 59819
rect 85726 59695 85750 59751
rect 85806 59695 85830 59751
rect 85726 59662 85830 59695
rect 85850 59999 86326 60032
rect 85850 59943 85874 59999
rect 85930 59943 85998 59999
rect 86054 59943 86122 59999
rect 86178 59943 86246 59999
rect 86302 59943 86326 59999
rect 85850 59875 86326 59943
rect 85850 59819 85874 59875
rect 85930 59819 85998 59875
rect 86054 59819 86122 59875
rect 86178 59819 86246 59875
rect 86302 59819 86326 59875
rect 85850 59751 86326 59819
rect 85850 59695 85874 59751
rect 85930 59695 85998 59751
rect 86054 59695 86122 59751
rect 86178 59695 86246 59751
rect 86302 59695 86326 59751
rect 85850 59662 86326 59695
rect 1044 57089 1148 57140
rect 1044 57033 1068 57089
rect 1124 57033 1148 57089
rect 1044 56965 1148 57033
rect 1044 56909 1068 56965
rect 1124 56909 1148 56965
rect 1044 56841 1148 56909
rect 1044 56785 1068 56841
rect 1124 56785 1148 56841
rect 1044 56717 1148 56785
rect 1044 56661 1068 56717
rect 1124 56661 1148 56717
rect 1044 56593 1148 56661
rect 1044 56537 1068 56593
rect 1124 56537 1148 56593
rect 1044 56469 1148 56537
rect 1044 56413 1068 56469
rect 1124 56413 1148 56469
rect 1044 56345 1148 56413
rect 1044 56289 1068 56345
rect 1124 56289 1148 56345
rect 1044 56221 1148 56289
rect 1044 56165 1068 56221
rect 1124 56165 1148 56221
rect 1044 56097 1148 56165
rect 1044 56041 1068 56097
rect 1124 56041 1148 56097
rect 1044 55973 1148 56041
rect 1044 55917 1068 55973
rect 1124 55917 1148 55973
rect 1044 55849 1148 55917
rect 1044 55793 1068 55849
rect 1124 55793 1148 55849
rect 1044 55725 1148 55793
rect 1044 55669 1068 55725
rect 1124 55669 1148 55725
rect 1044 55601 1148 55669
rect 1044 55545 1068 55601
rect 1124 55545 1148 55601
rect 1044 55477 1148 55545
rect 1044 55421 1068 55477
rect 1124 55421 1148 55477
rect 1044 55353 1148 55421
rect 1044 55297 1068 55353
rect 1124 55297 1148 55353
rect 1044 55229 1148 55297
rect 1044 55173 1068 55229
rect 1124 55173 1148 55229
rect 1044 55105 1148 55173
rect 1044 55049 1068 55105
rect 1124 55049 1148 55105
rect 1044 54998 1148 55049
rect 1168 57089 1644 57140
rect 1168 57033 1192 57089
rect 1248 57033 1316 57089
rect 1372 57033 1440 57089
rect 1496 57033 1564 57089
rect 1620 57033 1644 57089
rect 1168 56965 1644 57033
rect 1168 56909 1192 56965
rect 1248 56909 1316 56965
rect 1372 56909 1440 56965
rect 1496 56909 1564 56965
rect 1620 56909 1644 56965
rect 1168 56841 1644 56909
rect 1168 56785 1192 56841
rect 1248 56785 1316 56841
rect 1372 56785 1440 56841
rect 1496 56785 1564 56841
rect 1620 56785 1644 56841
rect 1168 56717 1644 56785
rect 1168 56661 1192 56717
rect 1248 56661 1316 56717
rect 1372 56661 1440 56717
rect 1496 56661 1564 56717
rect 1620 56661 1644 56717
rect 1168 56593 1644 56661
rect 1168 56537 1192 56593
rect 1248 56537 1316 56593
rect 1372 56537 1440 56593
rect 1496 56537 1564 56593
rect 1620 56537 1644 56593
rect 1168 56469 1644 56537
rect 1168 56413 1192 56469
rect 1248 56413 1316 56469
rect 1372 56413 1440 56469
rect 1496 56413 1564 56469
rect 1620 56413 1644 56469
rect 1168 56345 1644 56413
rect 1168 56289 1192 56345
rect 1248 56289 1316 56345
rect 1372 56289 1440 56345
rect 1496 56289 1564 56345
rect 1620 56289 1644 56345
rect 1168 56221 1644 56289
rect 1168 56165 1192 56221
rect 1248 56165 1316 56221
rect 1372 56165 1440 56221
rect 1496 56165 1564 56221
rect 1620 56165 1644 56221
rect 1168 56097 1644 56165
rect 1168 56041 1192 56097
rect 1248 56041 1316 56097
rect 1372 56041 1440 56097
rect 1496 56041 1564 56097
rect 1620 56041 1644 56097
rect 1168 55973 1644 56041
rect 1168 55917 1192 55973
rect 1248 55917 1316 55973
rect 1372 55917 1440 55973
rect 1496 55917 1564 55973
rect 1620 55917 1644 55973
rect 1168 55849 1644 55917
rect 1168 55793 1192 55849
rect 1248 55793 1316 55849
rect 1372 55793 1440 55849
rect 1496 55793 1564 55849
rect 1620 55793 1644 55849
rect 1168 55725 1644 55793
rect 1168 55669 1192 55725
rect 1248 55669 1316 55725
rect 1372 55669 1440 55725
rect 1496 55669 1564 55725
rect 1620 55669 1644 55725
rect 1168 55601 1644 55669
rect 1168 55545 1192 55601
rect 1248 55545 1316 55601
rect 1372 55545 1440 55601
rect 1496 55545 1564 55601
rect 1620 55545 1644 55601
rect 1168 55477 1644 55545
rect 1168 55421 1192 55477
rect 1248 55421 1316 55477
rect 1372 55421 1440 55477
rect 1496 55421 1564 55477
rect 1620 55421 1644 55477
rect 1168 55353 1644 55421
rect 1168 55297 1192 55353
rect 1248 55297 1316 55353
rect 1372 55297 1440 55353
rect 1496 55297 1564 55353
rect 1620 55297 1644 55353
rect 1168 55229 1644 55297
rect 1168 55173 1192 55229
rect 1248 55173 1316 55229
rect 1372 55173 1440 55229
rect 1496 55173 1564 55229
rect 1620 55173 1644 55229
rect 1168 55105 1644 55173
rect 1168 55049 1192 55105
rect 1248 55049 1316 55105
rect 1372 55049 1440 55105
rect 1496 55049 1564 55105
rect 1620 55049 1644 55105
rect 1168 54998 1644 55049
rect 85726 57089 85830 57140
rect 85726 57033 85750 57089
rect 85806 57033 85830 57089
rect 85726 56965 85830 57033
rect 85726 56909 85750 56965
rect 85806 56909 85830 56965
rect 85726 56841 85830 56909
rect 85726 56785 85750 56841
rect 85806 56785 85830 56841
rect 85726 56717 85830 56785
rect 85726 56661 85750 56717
rect 85806 56661 85830 56717
rect 85726 56593 85830 56661
rect 85726 56537 85750 56593
rect 85806 56537 85830 56593
rect 85726 56469 85830 56537
rect 85726 56413 85750 56469
rect 85806 56413 85830 56469
rect 85726 56345 85830 56413
rect 85726 56289 85750 56345
rect 85806 56289 85830 56345
rect 85726 56221 85830 56289
rect 85726 56165 85750 56221
rect 85806 56165 85830 56221
rect 85726 56097 85830 56165
rect 85726 56041 85750 56097
rect 85806 56041 85830 56097
rect 85726 55973 85830 56041
rect 85726 55917 85750 55973
rect 85806 55917 85830 55973
rect 85726 55849 85830 55917
rect 85726 55793 85750 55849
rect 85806 55793 85830 55849
rect 85726 55725 85830 55793
rect 85726 55669 85750 55725
rect 85806 55669 85830 55725
rect 85726 55601 85830 55669
rect 85726 55545 85750 55601
rect 85806 55545 85830 55601
rect 85726 55477 85830 55545
rect 85726 55421 85750 55477
rect 85806 55421 85830 55477
rect 85726 55353 85830 55421
rect 85726 55297 85750 55353
rect 85806 55297 85830 55353
rect 85726 55229 85830 55297
rect 85726 55173 85750 55229
rect 85806 55173 85830 55229
rect 85726 55105 85830 55173
rect 85726 55049 85750 55105
rect 85806 55049 85830 55105
rect 85726 54998 85830 55049
rect 85850 57089 86326 57140
rect 85850 57033 85874 57089
rect 85930 57033 85998 57089
rect 86054 57033 86122 57089
rect 86178 57033 86246 57089
rect 86302 57033 86326 57089
rect 85850 56965 86326 57033
rect 85850 56909 85874 56965
rect 85930 56909 85998 56965
rect 86054 56909 86122 56965
rect 86178 56909 86246 56965
rect 86302 56909 86326 56965
rect 85850 56841 86326 56909
rect 85850 56785 85874 56841
rect 85930 56785 85998 56841
rect 86054 56785 86122 56841
rect 86178 56785 86246 56841
rect 86302 56785 86326 56841
rect 85850 56717 86326 56785
rect 85850 56661 85874 56717
rect 85930 56661 85998 56717
rect 86054 56661 86122 56717
rect 86178 56661 86246 56717
rect 86302 56661 86326 56717
rect 85850 56593 86326 56661
rect 85850 56537 85874 56593
rect 85930 56537 85998 56593
rect 86054 56537 86122 56593
rect 86178 56537 86246 56593
rect 86302 56537 86326 56593
rect 85850 56469 86326 56537
rect 85850 56413 85874 56469
rect 85930 56413 85998 56469
rect 86054 56413 86122 56469
rect 86178 56413 86246 56469
rect 86302 56413 86326 56469
rect 85850 56345 86326 56413
rect 85850 56289 85874 56345
rect 85930 56289 85998 56345
rect 86054 56289 86122 56345
rect 86178 56289 86246 56345
rect 86302 56289 86326 56345
rect 85850 56221 86326 56289
rect 85850 56165 85874 56221
rect 85930 56165 85998 56221
rect 86054 56165 86122 56221
rect 86178 56165 86246 56221
rect 86302 56165 86326 56221
rect 85850 56097 86326 56165
rect 85850 56041 85874 56097
rect 85930 56041 85998 56097
rect 86054 56041 86122 56097
rect 86178 56041 86246 56097
rect 86302 56041 86326 56097
rect 85850 55973 86326 56041
rect 85850 55917 85874 55973
rect 85930 55917 85998 55973
rect 86054 55917 86122 55973
rect 86178 55917 86246 55973
rect 86302 55917 86326 55973
rect 85850 55849 86326 55917
rect 85850 55793 85874 55849
rect 85930 55793 85998 55849
rect 86054 55793 86122 55849
rect 86178 55793 86246 55849
rect 86302 55793 86326 55849
rect 85850 55725 86326 55793
rect 85850 55669 85874 55725
rect 85930 55669 85998 55725
rect 86054 55669 86122 55725
rect 86178 55669 86246 55725
rect 86302 55669 86326 55725
rect 85850 55601 86326 55669
rect 85850 55545 85874 55601
rect 85930 55545 85998 55601
rect 86054 55545 86122 55601
rect 86178 55545 86246 55601
rect 86302 55545 86326 55601
rect 85850 55477 86326 55545
rect 85850 55421 85874 55477
rect 85930 55421 85998 55477
rect 86054 55421 86122 55477
rect 86178 55421 86246 55477
rect 86302 55421 86326 55477
rect 85850 55353 86326 55421
rect 85850 55297 85874 55353
rect 85930 55297 85998 55353
rect 86054 55297 86122 55353
rect 86178 55297 86246 55353
rect 86302 55297 86326 55353
rect 85850 55229 86326 55297
rect 85850 55173 85874 55229
rect 85930 55173 85998 55229
rect 86054 55173 86122 55229
rect 86178 55173 86246 55229
rect 86302 55173 86326 55229
rect 85850 55105 86326 55173
rect 85850 55049 85874 55105
rect 85930 55049 85998 55105
rect 86054 55049 86122 55105
rect 86178 55049 86246 55105
rect 86302 55049 86326 55105
rect 85850 54998 86326 55049
rect 1844 54787 1948 54848
rect 1844 54731 1868 54787
rect 1924 54731 1948 54787
rect 1844 54663 1948 54731
rect 1844 54607 1868 54663
rect 1924 54607 1948 54663
rect 1844 54539 1948 54607
rect 1844 54483 1868 54539
rect 1924 54483 1948 54539
rect 1844 54415 1948 54483
rect 1844 54359 1868 54415
rect 1924 54359 1948 54415
rect 1844 54291 1948 54359
rect 1844 54235 1868 54291
rect 1924 54235 1948 54291
rect 1844 54167 1948 54235
rect 1844 54111 1868 54167
rect 1924 54111 1948 54167
rect 1844 54043 1948 54111
rect 1844 53987 1868 54043
rect 1924 53987 1948 54043
rect 1844 53919 1948 53987
rect 1844 53863 1868 53919
rect 1924 53863 1948 53919
rect 1844 53795 1948 53863
rect 1844 53739 1868 53795
rect 1924 53739 1948 53795
rect 1844 53671 1948 53739
rect 1844 53615 1868 53671
rect 1924 53615 1948 53671
rect 1844 53547 1948 53615
rect 1844 53491 1868 53547
rect 1924 53491 1948 53547
rect 1844 53423 1948 53491
rect 1844 53367 1868 53423
rect 1924 53367 1948 53423
rect 1844 53299 1948 53367
rect 1844 53243 1868 53299
rect 1924 53243 1948 53299
rect 1844 53175 1948 53243
rect 1844 53119 1868 53175
rect 1924 53119 1948 53175
rect 1844 53051 1948 53119
rect 1844 52995 1868 53051
rect 1924 52995 1948 53051
rect 1844 52927 1948 52995
rect 1844 52871 1868 52927
rect 1924 52871 1948 52927
rect 1844 52803 1948 52871
rect 1844 52747 1868 52803
rect 1924 52747 1948 52803
rect 1844 52679 1948 52747
rect 1844 52623 1868 52679
rect 1924 52623 1948 52679
rect 1844 52555 1948 52623
rect 1844 52499 1868 52555
rect 1924 52499 1948 52555
rect 1844 52431 1948 52499
rect 1844 52375 1868 52431
rect 1924 52375 1948 52431
rect 1844 52307 1948 52375
rect 1844 52251 1868 52307
rect 1924 52251 1948 52307
rect 1844 52183 1948 52251
rect 1844 52127 1868 52183
rect 1924 52127 1948 52183
rect 1844 52059 1948 52127
rect 1844 52003 1868 52059
rect 1924 52003 1948 52059
rect 1844 51935 1948 52003
rect 1844 51879 1868 51935
rect 1924 51879 1948 51935
rect 1844 51811 1948 51879
rect 1844 51755 1868 51811
rect 1924 51755 1948 51811
rect 1844 51687 1948 51755
rect 1844 51631 1868 51687
rect 1924 51631 1948 51687
rect 1844 51563 1948 51631
rect 1844 51507 1868 51563
rect 1924 51507 1948 51563
rect 1844 51446 1948 51507
rect 1968 54787 2444 54848
rect 1968 54731 1992 54787
rect 2048 54731 2116 54787
rect 2172 54731 2240 54787
rect 2296 54731 2364 54787
rect 2420 54731 2444 54787
rect 1968 54663 2444 54731
rect 1968 54607 1992 54663
rect 2048 54607 2116 54663
rect 2172 54607 2240 54663
rect 2296 54607 2364 54663
rect 2420 54607 2444 54663
rect 1968 54539 2444 54607
rect 1968 54483 1992 54539
rect 2048 54483 2116 54539
rect 2172 54483 2240 54539
rect 2296 54483 2364 54539
rect 2420 54483 2444 54539
rect 1968 54415 2444 54483
rect 1968 54359 1992 54415
rect 2048 54359 2116 54415
rect 2172 54359 2240 54415
rect 2296 54359 2364 54415
rect 2420 54359 2444 54415
rect 1968 54291 2444 54359
rect 1968 54235 1992 54291
rect 2048 54235 2116 54291
rect 2172 54235 2240 54291
rect 2296 54235 2364 54291
rect 2420 54235 2444 54291
rect 1968 54167 2444 54235
rect 1968 54111 1992 54167
rect 2048 54111 2116 54167
rect 2172 54111 2240 54167
rect 2296 54111 2364 54167
rect 2420 54111 2444 54167
rect 1968 54043 2444 54111
rect 1968 53987 1992 54043
rect 2048 53987 2116 54043
rect 2172 53987 2240 54043
rect 2296 53987 2364 54043
rect 2420 53987 2444 54043
rect 1968 53919 2444 53987
rect 1968 53863 1992 53919
rect 2048 53863 2116 53919
rect 2172 53863 2240 53919
rect 2296 53863 2364 53919
rect 2420 53863 2444 53919
rect 1968 53795 2444 53863
rect 1968 53739 1992 53795
rect 2048 53739 2116 53795
rect 2172 53739 2240 53795
rect 2296 53739 2364 53795
rect 2420 53739 2444 53795
rect 1968 53671 2444 53739
rect 1968 53615 1992 53671
rect 2048 53615 2116 53671
rect 2172 53615 2240 53671
rect 2296 53615 2364 53671
rect 2420 53615 2444 53671
rect 1968 53547 2444 53615
rect 1968 53491 1992 53547
rect 2048 53491 2116 53547
rect 2172 53491 2240 53547
rect 2296 53491 2364 53547
rect 2420 53491 2444 53547
rect 1968 53423 2444 53491
rect 1968 53367 1992 53423
rect 2048 53367 2116 53423
rect 2172 53367 2240 53423
rect 2296 53367 2364 53423
rect 2420 53367 2444 53423
rect 1968 53299 2444 53367
rect 1968 53243 1992 53299
rect 2048 53243 2116 53299
rect 2172 53243 2240 53299
rect 2296 53243 2364 53299
rect 2420 53243 2444 53299
rect 1968 53175 2444 53243
rect 1968 53119 1992 53175
rect 2048 53119 2116 53175
rect 2172 53119 2240 53175
rect 2296 53119 2364 53175
rect 2420 53119 2444 53175
rect 1968 53051 2444 53119
rect 1968 52995 1992 53051
rect 2048 52995 2116 53051
rect 2172 52995 2240 53051
rect 2296 52995 2364 53051
rect 2420 52995 2444 53051
rect 1968 52927 2444 52995
rect 1968 52871 1992 52927
rect 2048 52871 2116 52927
rect 2172 52871 2240 52927
rect 2296 52871 2364 52927
rect 2420 52871 2444 52927
rect 1968 52803 2444 52871
rect 1968 52747 1992 52803
rect 2048 52747 2116 52803
rect 2172 52747 2240 52803
rect 2296 52747 2364 52803
rect 2420 52747 2444 52803
rect 1968 52679 2444 52747
rect 1968 52623 1992 52679
rect 2048 52623 2116 52679
rect 2172 52623 2240 52679
rect 2296 52623 2364 52679
rect 2420 52623 2444 52679
rect 1968 52555 2444 52623
rect 1968 52499 1992 52555
rect 2048 52499 2116 52555
rect 2172 52499 2240 52555
rect 2296 52499 2364 52555
rect 2420 52499 2444 52555
rect 1968 52431 2444 52499
rect 1968 52375 1992 52431
rect 2048 52375 2116 52431
rect 2172 52375 2240 52431
rect 2296 52375 2364 52431
rect 2420 52375 2444 52431
rect 1968 52307 2444 52375
rect 1968 52251 1992 52307
rect 2048 52251 2116 52307
rect 2172 52251 2240 52307
rect 2296 52251 2364 52307
rect 2420 52251 2444 52307
rect 1968 52183 2444 52251
rect 1968 52127 1992 52183
rect 2048 52127 2116 52183
rect 2172 52127 2240 52183
rect 2296 52127 2364 52183
rect 2420 52127 2444 52183
rect 1968 52059 2444 52127
rect 1968 52003 1992 52059
rect 2048 52003 2116 52059
rect 2172 52003 2240 52059
rect 2296 52003 2364 52059
rect 2420 52003 2444 52059
rect 1968 51935 2444 52003
rect 1968 51879 1992 51935
rect 2048 51879 2116 51935
rect 2172 51879 2240 51935
rect 2296 51879 2364 51935
rect 2420 51879 2444 51935
rect 1968 51811 2444 51879
rect 1968 51755 1992 51811
rect 2048 51755 2116 51811
rect 2172 51755 2240 51811
rect 2296 51755 2364 51811
rect 2420 51755 2444 51811
rect 1968 51687 2444 51755
rect 1968 51631 1992 51687
rect 2048 51631 2116 51687
rect 2172 51631 2240 51687
rect 2296 51631 2364 51687
rect 2420 51631 2444 51687
rect 1968 51563 2444 51631
rect 1968 51507 1992 51563
rect 2048 51507 2116 51563
rect 2172 51507 2240 51563
rect 2296 51507 2364 51563
rect 2420 51507 2444 51563
rect 1968 51446 2444 51507
rect 86526 54787 86630 54848
rect 86526 54731 86550 54787
rect 86606 54731 86630 54787
rect 86526 54663 86630 54731
rect 86526 54607 86550 54663
rect 86606 54607 86630 54663
rect 86526 54539 86630 54607
rect 86526 54483 86550 54539
rect 86606 54483 86630 54539
rect 86526 54415 86630 54483
rect 86526 54359 86550 54415
rect 86606 54359 86630 54415
rect 86526 54291 86630 54359
rect 86526 54235 86550 54291
rect 86606 54235 86630 54291
rect 86526 54167 86630 54235
rect 86526 54111 86550 54167
rect 86606 54111 86630 54167
rect 86526 54043 86630 54111
rect 86526 53987 86550 54043
rect 86606 53987 86630 54043
rect 86526 53919 86630 53987
rect 86526 53863 86550 53919
rect 86606 53863 86630 53919
rect 86526 53795 86630 53863
rect 86526 53739 86550 53795
rect 86606 53739 86630 53795
rect 86526 53671 86630 53739
rect 86526 53615 86550 53671
rect 86606 53615 86630 53671
rect 86526 53547 86630 53615
rect 86526 53491 86550 53547
rect 86606 53491 86630 53547
rect 86526 53423 86630 53491
rect 86526 53367 86550 53423
rect 86606 53367 86630 53423
rect 86526 53299 86630 53367
rect 86526 53243 86550 53299
rect 86606 53243 86630 53299
rect 86526 53175 86630 53243
rect 86526 53119 86550 53175
rect 86606 53119 86630 53175
rect 86526 53051 86630 53119
rect 86526 52995 86550 53051
rect 86606 52995 86630 53051
rect 86526 52927 86630 52995
rect 86526 52871 86550 52927
rect 86606 52871 86630 52927
rect 86526 52803 86630 52871
rect 86526 52747 86550 52803
rect 86606 52747 86630 52803
rect 86526 52679 86630 52747
rect 86526 52623 86550 52679
rect 86606 52623 86630 52679
rect 86526 52555 86630 52623
rect 86526 52499 86550 52555
rect 86606 52499 86630 52555
rect 86526 52431 86630 52499
rect 86526 52375 86550 52431
rect 86606 52375 86630 52431
rect 86526 52307 86630 52375
rect 86526 52251 86550 52307
rect 86606 52251 86630 52307
rect 86526 52183 86630 52251
rect 86526 52127 86550 52183
rect 86606 52127 86630 52183
rect 86526 52059 86630 52127
rect 86526 52003 86550 52059
rect 86606 52003 86630 52059
rect 86526 51935 86630 52003
rect 86526 51879 86550 51935
rect 86606 51879 86630 51935
rect 86526 51811 86630 51879
rect 86526 51755 86550 51811
rect 86606 51755 86630 51811
rect 86526 51687 86630 51755
rect 86526 51631 86550 51687
rect 86606 51631 86630 51687
rect 86526 51563 86630 51631
rect 86526 51507 86550 51563
rect 86606 51507 86630 51563
rect 86526 51446 86630 51507
rect 86650 54787 87126 54848
rect 86650 54731 86674 54787
rect 86730 54731 86798 54787
rect 86854 54731 86922 54787
rect 86978 54731 87046 54787
rect 87102 54731 87126 54787
rect 86650 54663 87126 54731
rect 86650 54607 86674 54663
rect 86730 54607 86798 54663
rect 86854 54607 86922 54663
rect 86978 54607 87046 54663
rect 87102 54607 87126 54663
rect 86650 54539 87126 54607
rect 86650 54483 86674 54539
rect 86730 54483 86798 54539
rect 86854 54483 86922 54539
rect 86978 54483 87046 54539
rect 87102 54483 87126 54539
rect 86650 54415 87126 54483
rect 86650 54359 86674 54415
rect 86730 54359 86798 54415
rect 86854 54359 86922 54415
rect 86978 54359 87046 54415
rect 87102 54359 87126 54415
rect 86650 54291 87126 54359
rect 86650 54235 86674 54291
rect 86730 54235 86798 54291
rect 86854 54235 86922 54291
rect 86978 54235 87046 54291
rect 87102 54235 87126 54291
rect 86650 54167 87126 54235
rect 86650 54111 86674 54167
rect 86730 54111 86798 54167
rect 86854 54111 86922 54167
rect 86978 54111 87046 54167
rect 87102 54111 87126 54167
rect 86650 54043 87126 54111
rect 86650 53987 86674 54043
rect 86730 53987 86798 54043
rect 86854 53987 86922 54043
rect 86978 53987 87046 54043
rect 87102 53987 87126 54043
rect 86650 53919 87126 53987
rect 86650 53863 86674 53919
rect 86730 53863 86798 53919
rect 86854 53863 86922 53919
rect 86978 53863 87046 53919
rect 87102 53863 87126 53919
rect 86650 53795 87126 53863
rect 86650 53739 86674 53795
rect 86730 53739 86798 53795
rect 86854 53739 86922 53795
rect 86978 53739 87046 53795
rect 87102 53739 87126 53795
rect 86650 53671 87126 53739
rect 86650 53615 86674 53671
rect 86730 53615 86798 53671
rect 86854 53615 86922 53671
rect 86978 53615 87046 53671
rect 87102 53615 87126 53671
rect 86650 53547 87126 53615
rect 86650 53491 86674 53547
rect 86730 53491 86798 53547
rect 86854 53491 86922 53547
rect 86978 53491 87046 53547
rect 87102 53491 87126 53547
rect 86650 53423 87126 53491
rect 86650 53367 86674 53423
rect 86730 53367 86798 53423
rect 86854 53367 86922 53423
rect 86978 53367 87046 53423
rect 87102 53367 87126 53423
rect 86650 53299 87126 53367
rect 86650 53243 86674 53299
rect 86730 53243 86798 53299
rect 86854 53243 86922 53299
rect 86978 53243 87046 53299
rect 87102 53243 87126 53299
rect 86650 53175 87126 53243
rect 86650 53119 86674 53175
rect 86730 53119 86798 53175
rect 86854 53119 86922 53175
rect 86978 53119 87046 53175
rect 87102 53119 87126 53175
rect 86650 53051 87126 53119
rect 86650 52995 86674 53051
rect 86730 52995 86798 53051
rect 86854 52995 86922 53051
rect 86978 52995 87046 53051
rect 87102 52995 87126 53051
rect 86650 52927 87126 52995
rect 86650 52871 86674 52927
rect 86730 52871 86798 52927
rect 86854 52871 86922 52927
rect 86978 52871 87046 52927
rect 87102 52871 87126 52927
rect 86650 52803 87126 52871
rect 86650 52747 86674 52803
rect 86730 52747 86798 52803
rect 86854 52747 86922 52803
rect 86978 52747 87046 52803
rect 87102 52747 87126 52803
rect 86650 52679 87126 52747
rect 86650 52623 86674 52679
rect 86730 52623 86798 52679
rect 86854 52623 86922 52679
rect 86978 52623 87046 52679
rect 87102 52623 87126 52679
rect 86650 52555 87126 52623
rect 86650 52499 86674 52555
rect 86730 52499 86798 52555
rect 86854 52499 86922 52555
rect 86978 52499 87046 52555
rect 87102 52499 87126 52555
rect 86650 52431 87126 52499
rect 86650 52375 86674 52431
rect 86730 52375 86798 52431
rect 86854 52375 86922 52431
rect 86978 52375 87046 52431
rect 87102 52375 87126 52431
rect 86650 52307 87126 52375
rect 86650 52251 86674 52307
rect 86730 52251 86798 52307
rect 86854 52251 86922 52307
rect 86978 52251 87046 52307
rect 87102 52251 87126 52307
rect 86650 52183 87126 52251
rect 86650 52127 86674 52183
rect 86730 52127 86798 52183
rect 86854 52127 86922 52183
rect 86978 52127 87046 52183
rect 87102 52127 87126 52183
rect 86650 52059 87126 52127
rect 86650 52003 86674 52059
rect 86730 52003 86798 52059
rect 86854 52003 86922 52059
rect 86978 52003 87046 52059
rect 87102 52003 87126 52059
rect 86650 51935 87126 52003
rect 86650 51879 86674 51935
rect 86730 51879 86798 51935
rect 86854 51879 86922 51935
rect 86978 51879 87046 51935
rect 87102 51879 87126 51935
rect 86650 51811 87126 51879
rect 86650 51755 86674 51811
rect 86730 51755 86798 51811
rect 86854 51755 86922 51811
rect 86978 51755 87046 51811
rect 87102 51755 87126 51811
rect 86650 51687 87126 51755
rect 86650 51631 86674 51687
rect 86730 51631 86798 51687
rect 86854 51631 86922 51687
rect 86978 51631 87046 51687
rect 87102 51631 87126 51687
rect 86650 51563 87126 51631
rect 86650 51507 86674 51563
rect 86730 51507 86798 51563
rect 86854 51507 86922 51563
rect 86978 51507 87046 51563
rect 87102 51507 87126 51563
rect 86650 51446 87126 51507
rect 86526 47856 86630 47894
rect 86526 47800 86550 47856
rect 86606 47800 86630 47856
rect 86526 47732 86630 47800
rect 86526 47676 86550 47732
rect 86606 47676 86630 47732
rect 86526 47608 86630 47676
rect 86526 47552 86550 47608
rect 86606 47552 86630 47608
rect 86526 47484 86630 47552
rect 86526 47428 86550 47484
rect 86606 47428 86630 47484
rect 86526 47360 86630 47428
rect 86526 47304 86550 47360
rect 86606 47304 86630 47360
rect 86526 47236 86630 47304
rect 86526 47180 86550 47236
rect 86606 47180 86630 47236
rect 86526 47112 86630 47180
rect 86526 47056 86550 47112
rect 86606 47056 86630 47112
rect 86526 46988 86630 47056
rect 86526 46932 86550 46988
rect 86606 46932 86630 46988
rect 86526 46894 86630 46932
rect 86650 47856 87126 47894
rect 86650 47800 86674 47856
rect 86730 47800 86798 47856
rect 86854 47800 86922 47856
rect 86978 47800 87046 47856
rect 87102 47800 87126 47856
rect 86650 47732 87126 47800
rect 86650 47676 86674 47732
rect 86730 47676 86798 47732
rect 86854 47676 86922 47732
rect 86978 47676 87046 47732
rect 87102 47676 87126 47732
rect 86650 47608 87126 47676
rect 86650 47552 86674 47608
rect 86730 47552 86798 47608
rect 86854 47552 86922 47608
rect 86978 47552 87046 47608
rect 87102 47552 87126 47608
rect 86650 47484 87126 47552
rect 86650 47428 86674 47484
rect 86730 47428 86798 47484
rect 86854 47428 86922 47484
rect 86978 47428 87046 47484
rect 87102 47428 87126 47484
rect 86650 47360 87126 47428
rect 86650 47304 86674 47360
rect 86730 47304 86798 47360
rect 86854 47304 86922 47360
rect 86978 47304 87046 47360
rect 87102 47304 87126 47360
rect 86650 47236 87126 47304
rect 86650 47180 86674 47236
rect 86730 47180 86798 47236
rect 86854 47180 86922 47236
rect 86978 47180 87046 47236
rect 87102 47180 87126 47236
rect 86650 47112 87126 47180
rect 86650 47056 86674 47112
rect 86730 47056 86798 47112
rect 86854 47056 86922 47112
rect 86978 47056 87046 47112
rect 87102 47056 87126 47112
rect 86650 46988 87126 47056
rect 86650 46932 86674 46988
rect 86730 46932 86798 46988
rect 86854 46932 86922 46988
rect 86978 46932 87046 46988
rect 87102 46932 87126 46988
rect 86650 46894 87126 46932
rect 1044 46200 1148 46238
rect 1044 46144 1068 46200
rect 1124 46144 1148 46200
rect 1044 46076 1148 46144
rect 1044 46020 1068 46076
rect 1124 46020 1148 46076
rect 1044 45952 1148 46020
rect 1044 45896 1068 45952
rect 1124 45896 1148 45952
rect 1044 45828 1148 45896
rect 1044 45772 1068 45828
rect 1124 45772 1148 45828
rect 1044 45704 1148 45772
rect 1044 45648 1068 45704
rect 1124 45648 1148 45704
rect 1044 45580 1148 45648
rect 1044 45524 1068 45580
rect 1124 45524 1148 45580
rect 1044 45456 1148 45524
rect 1044 45400 1068 45456
rect 1124 45400 1148 45456
rect 1044 45332 1148 45400
rect 1044 45276 1068 45332
rect 1124 45276 1148 45332
rect 1044 45238 1148 45276
rect 1168 46200 1644 46238
rect 1168 46144 1192 46200
rect 1248 46144 1316 46200
rect 1372 46144 1440 46200
rect 1496 46144 1564 46200
rect 1620 46144 1644 46200
rect 1168 46076 1644 46144
rect 1168 46020 1192 46076
rect 1248 46020 1316 46076
rect 1372 46020 1440 46076
rect 1496 46020 1564 46076
rect 1620 46020 1644 46076
rect 1168 45952 1644 46020
rect 1168 45896 1192 45952
rect 1248 45896 1316 45952
rect 1372 45896 1440 45952
rect 1496 45896 1564 45952
rect 1620 45896 1644 45952
rect 1168 45828 1644 45896
rect 1168 45772 1192 45828
rect 1248 45772 1316 45828
rect 1372 45772 1440 45828
rect 1496 45772 1564 45828
rect 1620 45772 1644 45828
rect 1168 45704 1644 45772
rect 1168 45648 1192 45704
rect 1248 45648 1316 45704
rect 1372 45648 1440 45704
rect 1496 45648 1564 45704
rect 1620 45648 1644 45704
rect 1168 45580 1644 45648
rect 1168 45524 1192 45580
rect 1248 45524 1316 45580
rect 1372 45524 1440 45580
rect 1496 45524 1564 45580
rect 1620 45524 1644 45580
rect 1168 45456 1644 45524
rect 1168 45400 1192 45456
rect 1248 45400 1316 45456
rect 1372 45400 1440 45456
rect 1496 45400 1564 45456
rect 1620 45400 1644 45456
rect 1168 45332 1644 45400
rect 1168 45276 1192 45332
rect 1248 45276 1316 45332
rect 1372 45276 1440 45332
rect 1496 45276 1564 45332
rect 1620 45276 1644 45332
rect 1168 45238 1644 45276
rect 85726 46200 85830 46238
rect 85726 46144 85750 46200
rect 85806 46144 85830 46200
rect 85726 46076 85830 46144
rect 85726 46020 85750 46076
rect 85806 46020 85830 46076
rect 85726 45952 85830 46020
rect 85726 45896 85750 45952
rect 85806 45896 85830 45952
rect 85726 45828 85830 45896
rect 85726 45772 85750 45828
rect 85806 45772 85830 45828
rect 85726 45704 85830 45772
rect 85726 45648 85750 45704
rect 85806 45648 85830 45704
rect 85726 45580 85830 45648
rect 85726 45524 85750 45580
rect 85806 45524 85830 45580
rect 85726 45456 85830 45524
rect 85726 45400 85750 45456
rect 85806 45400 85830 45456
rect 85726 45332 85830 45400
rect 85726 45276 85750 45332
rect 85806 45276 85830 45332
rect 85726 45238 85830 45276
rect 85850 46200 86326 46238
rect 85850 46144 85874 46200
rect 85930 46144 85998 46200
rect 86054 46144 86122 46200
rect 86178 46144 86246 46200
rect 86302 46144 86326 46200
rect 85850 46076 86326 46144
rect 85850 46020 85874 46076
rect 85930 46020 85998 46076
rect 86054 46020 86122 46076
rect 86178 46020 86246 46076
rect 86302 46020 86326 46076
rect 85850 45952 86326 46020
rect 85850 45896 85874 45952
rect 85930 45896 85998 45952
rect 86054 45896 86122 45952
rect 86178 45896 86246 45952
rect 86302 45896 86326 45952
rect 85850 45828 86326 45896
rect 85850 45772 85874 45828
rect 85930 45772 85998 45828
rect 86054 45772 86122 45828
rect 86178 45772 86246 45828
rect 86302 45772 86326 45828
rect 85850 45704 86326 45772
rect 85850 45648 85874 45704
rect 85930 45648 85998 45704
rect 86054 45648 86122 45704
rect 86178 45648 86246 45704
rect 86302 45648 86326 45704
rect 85850 45580 86326 45648
rect 85850 45524 85874 45580
rect 85930 45524 85998 45580
rect 86054 45524 86122 45580
rect 86178 45524 86246 45580
rect 86302 45524 86326 45580
rect 85850 45456 86326 45524
rect 85850 45400 85874 45456
rect 85930 45400 85998 45456
rect 86054 45400 86122 45456
rect 86178 45400 86246 45456
rect 86302 45400 86326 45456
rect 85850 45332 86326 45400
rect 85850 45276 85874 45332
rect 85930 45276 85998 45332
rect 86054 45276 86122 45332
rect 86178 45276 86246 45332
rect 86302 45276 86326 45332
rect 85850 45238 86326 45276
rect 1906 34614 2382 34640
rect 1906 34558 1930 34614
rect 1986 34558 2054 34614
rect 2110 34558 2178 34614
rect 2234 34558 2302 34614
rect 2358 34558 2382 34614
rect 1906 34490 2382 34558
rect 1906 34434 1930 34490
rect 1986 34434 2054 34490
rect 2110 34434 2178 34490
rect 2234 34434 2302 34490
rect 2358 34434 2382 34490
rect 1906 34366 2382 34434
rect 1906 34310 1930 34366
rect 1986 34310 2054 34366
rect 2110 34310 2178 34366
rect 2234 34310 2302 34366
rect 2358 34310 2382 34366
rect 1906 34242 2382 34310
rect 1906 34186 1930 34242
rect 1986 34186 2054 34242
rect 2110 34186 2178 34242
rect 2234 34186 2302 34242
rect 2358 34186 2382 34242
rect 1906 34160 2382 34186
rect 86588 34459 87064 34516
rect 86588 34403 86612 34459
rect 86668 34403 86736 34459
rect 86792 34403 86860 34459
rect 86916 34403 86984 34459
rect 87040 34403 87064 34459
rect 86588 34335 87064 34403
rect 86588 34279 86612 34335
rect 86668 34279 86736 34335
rect 86792 34279 86860 34335
rect 86916 34279 86984 34335
rect 87040 34279 87064 34335
rect 86588 34211 87064 34279
rect 86588 34155 86612 34211
rect 86668 34155 86736 34211
rect 86792 34155 86860 34211
rect 86916 34155 86984 34211
rect 87040 34155 87064 34211
rect 86588 34087 87064 34155
rect 86588 34031 86612 34087
rect 86668 34031 86736 34087
rect 86792 34031 86860 34087
rect 86916 34031 86984 34087
rect 87040 34031 87064 34087
rect 86588 33974 87064 34031
rect 1106 33264 1582 33276
rect 1106 33208 1130 33264
rect 1186 33208 1254 33264
rect 1310 33208 1378 33264
rect 1434 33208 1502 33264
rect 1558 33208 1582 33264
rect 1106 33140 1582 33208
rect 1106 33084 1130 33140
rect 1186 33084 1254 33140
rect 1310 33084 1378 33140
rect 1434 33084 1502 33140
rect 1558 33084 1582 33140
rect 1106 33016 1582 33084
rect 1106 32960 1130 33016
rect 1186 32960 1254 33016
rect 1310 32960 1378 33016
rect 1434 32960 1502 33016
rect 1558 32960 1582 33016
rect 1106 32892 1582 32960
rect 1106 32836 1130 32892
rect 1186 32836 1254 32892
rect 1310 32836 1378 32892
rect 1434 32836 1502 32892
rect 1558 32836 1582 32892
rect 1106 32824 1582 32836
rect 85788 33264 86264 33276
rect 85788 33208 85812 33264
rect 85868 33208 85936 33264
rect 85992 33208 86060 33264
rect 86116 33208 86184 33264
rect 86240 33208 86264 33264
rect 85788 33140 86264 33208
rect 85788 33084 85812 33140
rect 85868 33084 85936 33140
rect 85992 33084 86060 33140
rect 86116 33084 86184 33140
rect 86240 33084 86264 33140
rect 85788 33016 86264 33084
rect 85788 32960 85812 33016
rect 85868 32960 85936 33016
rect 85992 32960 86060 33016
rect 86116 32960 86184 33016
rect 86240 32960 86264 33016
rect 85788 32892 86264 32960
rect 85788 32836 85812 32892
rect 85868 32836 85936 32892
rect 85992 32836 86060 32892
rect 86116 32836 86184 32892
rect 86240 32836 86264 32892
rect 85788 32824 86264 32836
rect 86588 32364 87064 32376
rect 86588 32308 86612 32364
rect 86668 32308 86736 32364
rect 86792 32308 86860 32364
rect 86916 32308 86984 32364
rect 87040 32308 87064 32364
rect 1906 32240 2382 32300
rect 1906 32184 1930 32240
rect 1986 32184 2054 32240
rect 2110 32184 2178 32240
rect 2234 32184 2302 32240
rect 2358 32184 2382 32240
rect 1906 32116 2382 32184
rect 1906 32060 1930 32116
rect 1986 32060 2054 32116
rect 2110 32060 2178 32116
rect 2234 32060 2302 32116
rect 2358 32060 2382 32116
rect 1906 32000 2382 32060
rect 86588 32240 87064 32308
rect 86588 32184 86612 32240
rect 86668 32184 86736 32240
rect 86792 32184 86860 32240
rect 86916 32184 86984 32240
rect 87040 32184 87064 32240
rect 86588 32116 87064 32184
rect 86588 32060 86612 32116
rect 86668 32060 86736 32116
rect 86792 32060 86860 32116
rect 86916 32060 86984 32116
rect 87040 32060 87064 32116
rect 86588 31992 87064 32060
rect 86588 31936 86612 31992
rect 86668 31936 86736 31992
rect 86792 31936 86860 31992
rect 86916 31936 86984 31992
rect 87040 31936 87064 31992
rect 86588 31924 87064 31936
rect 1106 31464 1582 31476
rect 1106 31408 1130 31464
rect 1186 31408 1254 31464
rect 1310 31408 1378 31464
rect 1434 31408 1502 31464
rect 1558 31408 1582 31464
rect 1106 31340 1582 31408
rect 1106 31284 1130 31340
rect 1186 31284 1254 31340
rect 1310 31284 1378 31340
rect 1434 31284 1502 31340
rect 1558 31284 1582 31340
rect 1106 31216 1582 31284
rect 1106 31160 1130 31216
rect 1186 31160 1254 31216
rect 1310 31160 1378 31216
rect 1434 31160 1502 31216
rect 1558 31160 1582 31216
rect 1106 31092 1582 31160
rect 1106 31036 1130 31092
rect 1186 31036 1254 31092
rect 1310 31036 1378 31092
rect 1434 31036 1502 31092
rect 1558 31036 1582 31092
rect 1106 31024 1582 31036
rect 85788 31464 86264 31476
rect 85788 31408 85812 31464
rect 85868 31408 85936 31464
rect 85992 31408 86060 31464
rect 86116 31408 86184 31464
rect 86240 31408 86264 31464
rect 85788 31340 86264 31408
rect 85788 31284 85812 31340
rect 85868 31284 85936 31340
rect 85992 31284 86060 31340
rect 86116 31284 86184 31340
rect 86240 31284 86264 31340
rect 85788 31216 86264 31284
rect 85788 31160 85812 31216
rect 85868 31160 85936 31216
rect 85992 31160 86060 31216
rect 86116 31160 86184 31216
rect 86240 31160 86264 31216
rect 85788 31092 86264 31160
rect 85788 31036 85812 31092
rect 85868 31036 85936 31092
rect 85992 31036 86060 31092
rect 86116 31036 86184 31092
rect 86240 31036 86264 31092
rect 85788 31024 86264 31036
rect 86588 30564 87064 30576
rect 86588 30508 86612 30564
rect 86668 30508 86736 30564
rect 86792 30508 86860 30564
rect 86916 30508 86984 30564
rect 87040 30508 87064 30564
rect 1906 30440 2382 30500
rect 1906 30384 1930 30440
rect 1986 30384 2054 30440
rect 2110 30384 2178 30440
rect 2234 30384 2302 30440
rect 2358 30384 2382 30440
rect 1906 30316 2382 30384
rect 1906 30260 1930 30316
rect 1986 30260 2054 30316
rect 2110 30260 2178 30316
rect 2234 30260 2302 30316
rect 2358 30260 2382 30316
rect 1906 30200 2382 30260
rect 86588 30440 87064 30508
rect 86588 30384 86612 30440
rect 86668 30384 86736 30440
rect 86792 30384 86860 30440
rect 86916 30384 86984 30440
rect 87040 30384 87064 30440
rect 86588 30316 87064 30384
rect 86588 30260 86612 30316
rect 86668 30260 86736 30316
rect 86792 30260 86860 30316
rect 86916 30260 86984 30316
rect 87040 30260 87064 30316
rect 86588 30192 87064 30260
rect 86588 30136 86612 30192
rect 86668 30136 86736 30192
rect 86792 30136 86860 30192
rect 86916 30136 86984 30192
rect 87040 30136 87064 30192
rect 86588 30124 87064 30136
rect 1106 29664 1582 29676
rect 1106 29608 1130 29664
rect 1186 29608 1254 29664
rect 1310 29608 1378 29664
rect 1434 29608 1502 29664
rect 1558 29608 1582 29664
rect 1106 29540 1582 29608
rect 1106 29484 1130 29540
rect 1186 29484 1254 29540
rect 1310 29484 1378 29540
rect 1434 29484 1502 29540
rect 1558 29484 1582 29540
rect 1106 29416 1582 29484
rect 1106 29360 1130 29416
rect 1186 29360 1254 29416
rect 1310 29360 1378 29416
rect 1434 29360 1502 29416
rect 1558 29360 1582 29416
rect 1106 29292 1582 29360
rect 1106 29236 1130 29292
rect 1186 29236 1254 29292
rect 1310 29236 1378 29292
rect 1434 29236 1502 29292
rect 1558 29236 1582 29292
rect 1106 29224 1582 29236
rect 85788 29664 86264 29676
rect 85788 29608 85812 29664
rect 85868 29608 85936 29664
rect 85992 29608 86060 29664
rect 86116 29608 86184 29664
rect 86240 29608 86264 29664
rect 85788 29540 86264 29608
rect 85788 29484 85812 29540
rect 85868 29484 85936 29540
rect 85992 29484 86060 29540
rect 86116 29484 86184 29540
rect 86240 29484 86264 29540
rect 85788 29416 86264 29484
rect 85788 29360 85812 29416
rect 85868 29360 85936 29416
rect 85992 29360 86060 29416
rect 86116 29360 86184 29416
rect 86240 29360 86264 29416
rect 85788 29292 86264 29360
rect 85788 29236 85812 29292
rect 85868 29236 85936 29292
rect 85992 29236 86060 29292
rect 86116 29236 86184 29292
rect 86240 29236 86264 29292
rect 85788 29224 86264 29236
rect 86588 28764 87064 28776
rect 86588 28708 86612 28764
rect 86668 28708 86736 28764
rect 86792 28708 86860 28764
rect 86916 28708 86984 28764
rect 87040 28708 87064 28764
rect 1906 28640 2382 28700
rect 1906 28584 1930 28640
rect 1986 28584 2054 28640
rect 2110 28584 2178 28640
rect 2234 28584 2302 28640
rect 2358 28584 2382 28640
rect 1906 28516 2382 28584
rect 1906 28460 1930 28516
rect 1986 28460 2054 28516
rect 2110 28460 2178 28516
rect 2234 28460 2302 28516
rect 2358 28460 2382 28516
rect 1906 28400 2382 28460
rect 86588 28640 87064 28708
rect 86588 28584 86612 28640
rect 86668 28584 86736 28640
rect 86792 28584 86860 28640
rect 86916 28584 86984 28640
rect 87040 28584 87064 28640
rect 86588 28516 87064 28584
rect 86588 28460 86612 28516
rect 86668 28460 86736 28516
rect 86792 28460 86860 28516
rect 86916 28460 86984 28516
rect 87040 28460 87064 28516
rect 86588 28392 87064 28460
rect 86588 28336 86612 28392
rect 86668 28336 86736 28392
rect 86792 28336 86860 28392
rect 86916 28336 86984 28392
rect 87040 28336 87064 28392
rect 86588 28324 87064 28336
rect 1106 27864 1582 27876
rect 1106 27808 1130 27864
rect 1186 27808 1254 27864
rect 1310 27808 1378 27864
rect 1434 27808 1502 27864
rect 1558 27808 1582 27864
rect 1106 27740 1582 27808
rect 1106 27684 1130 27740
rect 1186 27684 1254 27740
rect 1310 27684 1378 27740
rect 1434 27684 1502 27740
rect 1558 27684 1582 27740
rect 1106 27616 1582 27684
rect 1106 27560 1130 27616
rect 1186 27560 1254 27616
rect 1310 27560 1378 27616
rect 1434 27560 1502 27616
rect 1558 27560 1582 27616
rect 1106 27492 1582 27560
rect 1106 27436 1130 27492
rect 1186 27436 1254 27492
rect 1310 27436 1378 27492
rect 1434 27436 1502 27492
rect 1558 27436 1582 27492
rect 1106 27424 1582 27436
rect 85788 27864 86264 27876
rect 85788 27808 85812 27864
rect 85868 27808 85936 27864
rect 85992 27808 86060 27864
rect 86116 27808 86184 27864
rect 86240 27808 86264 27864
rect 85788 27740 86264 27808
rect 85788 27684 85812 27740
rect 85868 27684 85936 27740
rect 85992 27684 86060 27740
rect 86116 27684 86184 27740
rect 86240 27684 86264 27740
rect 85788 27616 86264 27684
rect 85788 27560 85812 27616
rect 85868 27560 85936 27616
rect 85992 27560 86060 27616
rect 86116 27560 86184 27616
rect 86240 27560 86264 27616
rect 85788 27492 86264 27560
rect 85788 27436 85812 27492
rect 85868 27436 85936 27492
rect 85992 27436 86060 27492
rect 86116 27436 86184 27492
rect 86240 27436 86264 27492
rect 85788 27424 86264 27436
rect 86588 26964 87064 26976
rect 86588 26908 86612 26964
rect 86668 26908 86736 26964
rect 86792 26908 86860 26964
rect 86916 26908 86984 26964
rect 87040 26908 87064 26964
rect 1906 26840 2382 26900
rect 1906 26784 1930 26840
rect 1986 26784 2054 26840
rect 2110 26784 2178 26840
rect 2234 26784 2302 26840
rect 2358 26784 2382 26840
rect 1906 26716 2382 26784
rect 1906 26660 1930 26716
rect 1986 26660 2054 26716
rect 2110 26660 2178 26716
rect 2234 26660 2302 26716
rect 2358 26660 2382 26716
rect 1906 26600 2382 26660
rect 86588 26840 87064 26908
rect 86588 26784 86612 26840
rect 86668 26784 86736 26840
rect 86792 26784 86860 26840
rect 86916 26784 86984 26840
rect 87040 26784 87064 26840
rect 86588 26716 87064 26784
rect 86588 26660 86612 26716
rect 86668 26660 86736 26716
rect 86792 26660 86860 26716
rect 86916 26660 86984 26716
rect 87040 26660 87064 26716
rect 86588 26592 87064 26660
rect 86588 26536 86612 26592
rect 86668 26536 86736 26592
rect 86792 26536 86860 26592
rect 86916 26536 86984 26592
rect 87040 26536 87064 26592
rect 86588 26524 87064 26536
rect 1106 26064 1582 26076
rect 1106 26008 1130 26064
rect 1186 26008 1254 26064
rect 1310 26008 1378 26064
rect 1434 26008 1502 26064
rect 1558 26008 1582 26064
rect 1106 25940 1582 26008
rect 1106 25884 1130 25940
rect 1186 25884 1254 25940
rect 1310 25884 1378 25940
rect 1434 25884 1502 25940
rect 1558 25884 1582 25940
rect 1106 25816 1582 25884
rect 1106 25760 1130 25816
rect 1186 25760 1254 25816
rect 1310 25760 1378 25816
rect 1434 25760 1502 25816
rect 1558 25760 1582 25816
rect 1106 25692 1582 25760
rect 1106 25636 1130 25692
rect 1186 25636 1254 25692
rect 1310 25636 1378 25692
rect 1434 25636 1502 25692
rect 1558 25636 1582 25692
rect 1106 25624 1582 25636
rect 85788 26064 86264 26076
rect 85788 26008 85812 26064
rect 85868 26008 85936 26064
rect 85992 26008 86060 26064
rect 86116 26008 86184 26064
rect 86240 26008 86264 26064
rect 85788 25940 86264 26008
rect 85788 25884 85812 25940
rect 85868 25884 85936 25940
rect 85992 25884 86060 25940
rect 86116 25884 86184 25940
rect 86240 25884 86264 25940
rect 85788 25816 86264 25884
rect 85788 25760 85812 25816
rect 85868 25760 85936 25816
rect 85992 25760 86060 25816
rect 86116 25760 86184 25816
rect 86240 25760 86264 25816
rect 85788 25692 86264 25760
rect 85788 25636 85812 25692
rect 85868 25636 85936 25692
rect 85992 25636 86060 25692
rect 86116 25636 86184 25692
rect 86240 25636 86264 25692
rect 85788 25624 86264 25636
rect 86588 25164 87064 25176
rect 86588 25108 86612 25164
rect 86668 25108 86736 25164
rect 86792 25108 86860 25164
rect 86916 25108 86984 25164
rect 87040 25108 87064 25164
rect 1906 25040 2382 25100
rect 1906 24984 1930 25040
rect 1986 24984 2054 25040
rect 2110 24984 2178 25040
rect 2234 24984 2302 25040
rect 2358 24984 2382 25040
rect 1906 24916 2382 24984
rect 1906 24860 1930 24916
rect 1986 24860 2054 24916
rect 2110 24860 2178 24916
rect 2234 24860 2302 24916
rect 2358 24860 2382 24916
rect 1906 24800 2382 24860
rect 86588 25040 87064 25108
rect 86588 24984 86612 25040
rect 86668 24984 86736 25040
rect 86792 24984 86860 25040
rect 86916 24984 86984 25040
rect 87040 24984 87064 25040
rect 86588 24916 87064 24984
rect 86588 24860 86612 24916
rect 86668 24860 86736 24916
rect 86792 24860 86860 24916
rect 86916 24860 86984 24916
rect 87040 24860 87064 24916
rect 86588 24792 87064 24860
rect 86588 24736 86612 24792
rect 86668 24736 86736 24792
rect 86792 24736 86860 24792
rect 86916 24736 86984 24792
rect 87040 24736 87064 24792
rect 86588 24724 87064 24736
rect 1106 24264 1582 24276
rect 1106 24208 1130 24264
rect 1186 24208 1254 24264
rect 1310 24208 1378 24264
rect 1434 24208 1502 24264
rect 1558 24208 1582 24264
rect 1106 24140 1582 24208
rect 1106 24084 1130 24140
rect 1186 24084 1254 24140
rect 1310 24084 1378 24140
rect 1434 24084 1502 24140
rect 1558 24084 1582 24140
rect 1106 24016 1582 24084
rect 1106 23960 1130 24016
rect 1186 23960 1254 24016
rect 1310 23960 1378 24016
rect 1434 23960 1502 24016
rect 1558 23960 1582 24016
rect 1106 23892 1582 23960
rect 1106 23836 1130 23892
rect 1186 23836 1254 23892
rect 1310 23836 1378 23892
rect 1434 23836 1502 23892
rect 1558 23836 1582 23892
rect 1106 23824 1582 23836
rect 85788 24264 86264 24276
rect 85788 24208 85812 24264
rect 85868 24208 85936 24264
rect 85992 24208 86060 24264
rect 86116 24208 86184 24264
rect 86240 24208 86264 24264
rect 85788 24140 86264 24208
rect 85788 24084 85812 24140
rect 85868 24084 85936 24140
rect 85992 24084 86060 24140
rect 86116 24084 86184 24140
rect 86240 24084 86264 24140
rect 85788 24016 86264 24084
rect 85788 23960 85812 24016
rect 85868 23960 85936 24016
rect 85992 23960 86060 24016
rect 86116 23960 86184 24016
rect 86240 23960 86264 24016
rect 85788 23892 86264 23960
rect 85788 23836 85812 23892
rect 85868 23836 85936 23892
rect 85992 23836 86060 23892
rect 86116 23836 86184 23892
rect 86240 23836 86264 23892
rect 85788 23824 86264 23836
rect 86588 23364 87064 23376
rect 86588 23308 86612 23364
rect 86668 23308 86736 23364
rect 86792 23308 86860 23364
rect 86916 23308 86984 23364
rect 87040 23308 87064 23364
rect 1906 23240 2382 23300
rect 1906 23184 1930 23240
rect 1986 23184 2054 23240
rect 2110 23184 2178 23240
rect 2234 23184 2302 23240
rect 2358 23184 2382 23240
rect 1906 23116 2382 23184
rect 1906 23060 1930 23116
rect 1986 23060 2054 23116
rect 2110 23060 2178 23116
rect 2234 23060 2302 23116
rect 2358 23060 2382 23116
rect 1906 23000 2382 23060
rect 86588 23240 87064 23308
rect 86588 23184 86612 23240
rect 86668 23184 86736 23240
rect 86792 23184 86860 23240
rect 86916 23184 86984 23240
rect 87040 23184 87064 23240
rect 86588 23116 87064 23184
rect 86588 23060 86612 23116
rect 86668 23060 86736 23116
rect 86792 23060 86860 23116
rect 86916 23060 86984 23116
rect 87040 23060 87064 23116
rect 86588 22992 87064 23060
rect 86588 22936 86612 22992
rect 86668 22936 86736 22992
rect 86792 22936 86860 22992
rect 86916 22936 86984 22992
rect 87040 22936 87064 22992
rect 86588 22924 87064 22936
rect 1106 22464 1582 22476
rect 1106 22408 1130 22464
rect 1186 22408 1254 22464
rect 1310 22408 1378 22464
rect 1434 22408 1502 22464
rect 1558 22408 1582 22464
rect 1106 22340 1582 22408
rect 1106 22284 1130 22340
rect 1186 22284 1254 22340
rect 1310 22284 1378 22340
rect 1434 22284 1502 22340
rect 1558 22284 1582 22340
rect 1106 22216 1582 22284
rect 1106 22160 1130 22216
rect 1186 22160 1254 22216
rect 1310 22160 1378 22216
rect 1434 22160 1502 22216
rect 1558 22160 1582 22216
rect 1106 22092 1582 22160
rect 1106 22036 1130 22092
rect 1186 22036 1254 22092
rect 1310 22036 1378 22092
rect 1434 22036 1502 22092
rect 1558 22036 1582 22092
rect 1106 22024 1582 22036
rect 85788 22464 86264 22476
rect 85788 22408 85812 22464
rect 85868 22408 85936 22464
rect 85992 22408 86060 22464
rect 86116 22408 86184 22464
rect 86240 22408 86264 22464
rect 85788 22340 86264 22408
rect 85788 22284 85812 22340
rect 85868 22284 85936 22340
rect 85992 22284 86060 22340
rect 86116 22284 86184 22340
rect 86240 22284 86264 22340
rect 85788 22216 86264 22284
rect 85788 22160 85812 22216
rect 85868 22160 85936 22216
rect 85992 22160 86060 22216
rect 86116 22160 86184 22216
rect 86240 22160 86264 22216
rect 85788 22092 86264 22160
rect 85788 22036 85812 22092
rect 85868 22036 85936 22092
rect 85992 22036 86060 22092
rect 86116 22036 86184 22092
rect 86240 22036 86264 22092
rect 85788 22024 86264 22036
rect 86588 21564 87064 21576
rect 86588 21508 86612 21564
rect 86668 21508 86736 21564
rect 86792 21508 86860 21564
rect 86916 21508 86984 21564
rect 87040 21508 87064 21564
rect 1906 21440 2382 21500
rect 1906 21384 1930 21440
rect 1986 21384 2054 21440
rect 2110 21384 2178 21440
rect 2234 21384 2302 21440
rect 2358 21384 2382 21440
rect 1906 21316 2382 21384
rect 1906 21260 1930 21316
rect 1986 21260 2054 21316
rect 2110 21260 2178 21316
rect 2234 21260 2302 21316
rect 2358 21260 2382 21316
rect 1906 21200 2382 21260
rect 86588 21440 87064 21508
rect 86588 21384 86612 21440
rect 86668 21384 86736 21440
rect 86792 21384 86860 21440
rect 86916 21384 86984 21440
rect 87040 21384 87064 21440
rect 86588 21316 87064 21384
rect 86588 21260 86612 21316
rect 86668 21260 86736 21316
rect 86792 21260 86860 21316
rect 86916 21260 86984 21316
rect 87040 21260 87064 21316
rect 86588 21192 87064 21260
rect 86588 21136 86612 21192
rect 86668 21136 86736 21192
rect 86792 21136 86860 21192
rect 86916 21136 86984 21192
rect 87040 21136 87064 21192
rect 86588 21124 87064 21136
rect 1106 20664 1582 20676
rect 1106 20608 1130 20664
rect 1186 20608 1254 20664
rect 1310 20608 1378 20664
rect 1434 20608 1502 20664
rect 1558 20608 1582 20664
rect 1106 20540 1582 20608
rect 1106 20484 1130 20540
rect 1186 20484 1254 20540
rect 1310 20484 1378 20540
rect 1434 20484 1502 20540
rect 1558 20484 1582 20540
rect 1106 20416 1582 20484
rect 1106 20360 1130 20416
rect 1186 20360 1254 20416
rect 1310 20360 1378 20416
rect 1434 20360 1502 20416
rect 1558 20360 1582 20416
rect 1106 20292 1582 20360
rect 1106 20236 1130 20292
rect 1186 20236 1254 20292
rect 1310 20236 1378 20292
rect 1434 20236 1502 20292
rect 1558 20236 1582 20292
rect 1106 20224 1582 20236
rect 85788 20664 86264 20676
rect 85788 20608 85812 20664
rect 85868 20608 85936 20664
rect 85992 20608 86060 20664
rect 86116 20608 86184 20664
rect 86240 20608 86264 20664
rect 85788 20540 86264 20608
rect 85788 20484 85812 20540
rect 85868 20484 85936 20540
rect 85992 20484 86060 20540
rect 86116 20484 86184 20540
rect 86240 20484 86264 20540
rect 85788 20416 86264 20484
rect 85788 20360 85812 20416
rect 85868 20360 85936 20416
rect 85992 20360 86060 20416
rect 86116 20360 86184 20416
rect 86240 20360 86264 20416
rect 85788 20292 86264 20360
rect 85788 20236 85812 20292
rect 85868 20236 85936 20292
rect 85992 20236 86060 20292
rect 86116 20236 86184 20292
rect 86240 20236 86264 20292
rect 85788 20224 86264 20236
rect 86588 19764 87064 19776
rect 86588 19708 86612 19764
rect 86668 19708 86736 19764
rect 86792 19708 86860 19764
rect 86916 19708 86984 19764
rect 87040 19708 87064 19764
rect 1906 19640 2382 19700
rect 1906 19584 1930 19640
rect 1986 19584 2054 19640
rect 2110 19584 2178 19640
rect 2234 19584 2302 19640
rect 2358 19584 2382 19640
rect 1906 19516 2382 19584
rect 1906 19460 1930 19516
rect 1986 19460 2054 19516
rect 2110 19460 2178 19516
rect 2234 19460 2302 19516
rect 2358 19460 2382 19516
rect 1906 19400 2382 19460
rect 86588 19640 87064 19708
rect 86588 19584 86612 19640
rect 86668 19584 86736 19640
rect 86792 19584 86860 19640
rect 86916 19584 86984 19640
rect 87040 19584 87064 19640
rect 86588 19516 87064 19584
rect 86588 19460 86612 19516
rect 86668 19460 86736 19516
rect 86792 19460 86860 19516
rect 86916 19460 86984 19516
rect 87040 19460 87064 19516
rect 86588 19392 87064 19460
rect 86588 19336 86612 19392
rect 86668 19336 86736 19392
rect 86792 19336 86860 19392
rect 86916 19336 86984 19392
rect 87040 19336 87064 19392
rect 86588 19324 87064 19336
rect 1106 18864 1582 18876
rect 1106 18808 1130 18864
rect 1186 18808 1254 18864
rect 1310 18808 1378 18864
rect 1434 18808 1502 18864
rect 1558 18808 1582 18864
rect 1106 18740 1582 18808
rect 1106 18684 1130 18740
rect 1186 18684 1254 18740
rect 1310 18684 1378 18740
rect 1434 18684 1502 18740
rect 1558 18684 1582 18740
rect 1106 18616 1582 18684
rect 1106 18560 1130 18616
rect 1186 18560 1254 18616
rect 1310 18560 1378 18616
rect 1434 18560 1502 18616
rect 1558 18560 1582 18616
rect 1106 18492 1582 18560
rect 1106 18436 1130 18492
rect 1186 18436 1254 18492
rect 1310 18436 1378 18492
rect 1434 18436 1502 18492
rect 1558 18436 1582 18492
rect 1106 18424 1582 18436
rect 85788 18864 86264 18876
rect 85788 18808 85812 18864
rect 85868 18808 85936 18864
rect 85992 18808 86060 18864
rect 86116 18808 86184 18864
rect 86240 18808 86264 18864
rect 85788 18740 86264 18808
rect 85788 18684 85812 18740
rect 85868 18684 85936 18740
rect 85992 18684 86060 18740
rect 86116 18684 86184 18740
rect 86240 18684 86264 18740
rect 85788 18616 86264 18684
rect 85788 18560 85812 18616
rect 85868 18560 85936 18616
rect 85992 18560 86060 18616
rect 86116 18560 86184 18616
rect 86240 18560 86264 18616
rect 85788 18492 86264 18560
rect 85788 18436 85812 18492
rect 85868 18436 85936 18492
rect 85992 18436 86060 18492
rect 86116 18436 86184 18492
rect 86240 18436 86264 18492
rect 85788 18424 86264 18436
rect 86588 17964 87064 17976
rect 86588 17908 86612 17964
rect 86668 17908 86736 17964
rect 86792 17908 86860 17964
rect 86916 17908 86984 17964
rect 87040 17908 87064 17964
rect 1906 17840 2382 17900
rect 1906 17784 1930 17840
rect 1986 17784 2054 17840
rect 2110 17784 2178 17840
rect 2234 17784 2302 17840
rect 2358 17784 2382 17840
rect 1906 17716 2382 17784
rect 1906 17660 1930 17716
rect 1986 17660 2054 17716
rect 2110 17660 2178 17716
rect 2234 17660 2302 17716
rect 2358 17660 2382 17716
rect 1906 17600 2382 17660
rect 86588 17840 87064 17908
rect 86588 17784 86612 17840
rect 86668 17784 86736 17840
rect 86792 17784 86860 17840
rect 86916 17784 86984 17840
rect 87040 17784 87064 17840
rect 86588 17716 87064 17784
rect 86588 17660 86612 17716
rect 86668 17660 86736 17716
rect 86792 17660 86860 17716
rect 86916 17660 86984 17716
rect 87040 17660 87064 17716
rect 86588 17592 87064 17660
rect 86588 17536 86612 17592
rect 86668 17536 86736 17592
rect 86792 17536 86860 17592
rect 86916 17536 86984 17592
rect 87040 17536 87064 17592
rect 86588 17524 87064 17536
rect 1106 17064 1582 17076
rect 1106 17008 1130 17064
rect 1186 17008 1254 17064
rect 1310 17008 1378 17064
rect 1434 17008 1502 17064
rect 1558 17008 1582 17064
rect 1106 16940 1582 17008
rect 1106 16884 1130 16940
rect 1186 16884 1254 16940
rect 1310 16884 1378 16940
rect 1434 16884 1502 16940
rect 1558 16884 1582 16940
rect 1106 16816 1582 16884
rect 1106 16760 1130 16816
rect 1186 16760 1254 16816
rect 1310 16760 1378 16816
rect 1434 16760 1502 16816
rect 1558 16760 1582 16816
rect 1106 16692 1582 16760
rect 1106 16636 1130 16692
rect 1186 16636 1254 16692
rect 1310 16636 1378 16692
rect 1434 16636 1502 16692
rect 1558 16636 1582 16692
rect 1106 16624 1582 16636
rect 85788 17064 86264 17076
rect 85788 17008 85812 17064
rect 85868 17008 85936 17064
rect 85992 17008 86060 17064
rect 86116 17008 86184 17064
rect 86240 17008 86264 17064
rect 85788 16940 86264 17008
rect 85788 16884 85812 16940
rect 85868 16884 85936 16940
rect 85992 16884 86060 16940
rect 86116 16884 86184 16940
rect 86240 16884 86264 16940
rect 85788 16816 86264 16884
rect 85788 16760 85812 16816
rect 85868 16760 85936 16816
rect 85992 16760 86060 16816
rect 86116 16760 86184 16816
rect 86240 16760 86264 16816
rect 85788 16692 86264 16760
rect 85788 16636 85812 16692
rect 85868 16636 85936 16692
rect 85992 16636 86060 16692
rect 86116 16636 86184 16692
rect 86240 16636 86264 16692
rect 85788 16624 86264 16636
rect 86588 16164 87064 16176
rect 86588 16108 86612 16164
rect 86668 16108 86736 16164
rect 86792 16108 86860 16164
rect 86916 16108 86984 16164
rect 87040 16108 87064 16164
rect 1906 16040 2382 16100
rect 1906 15984 1930 16040
rect 1986 15984 2054 16040
rect 2110 15984 2178 16040
rect 2234 15984 2302 16040
rect 2358 15984 2382 16040
rect 1906 15916 2382 15984
rect 1906 15860 1930 15916
rect 1986 15860 2054 15916
rect 2110 15860 2178 15916
rect 2234 15860 2302 15916
rect 2358 15860 2382 15916
rect 1906 15800 2382 15860
rect 86588 16040 87064 16108
rect 86588 15984 86612 16040
rect 86668 15984 86736 16040
rect 86792 15984 86860 16040
rect 86916 15984 86984 16040
rect 87040 15984 87064 16040
rect 86588 15916 87064 15984
rect 86588 15860 86612 15916
rect 86668 15860 86736 15916
rect 86792 15860 86860 15916
rect 86916 15860 86984 15916
rect 87040 15860 87064 15916
rect 86588 15792 87064 15860
rect 86588 15736 86612 15792
rect 86668 15736 86736 15792
rect 86792 15736 86860 15792
rect 86916 15736 86984 15792
rect 87040 15736 87064 15792
rect 86588 15724 87064 15736
rect 1106 15264 1582 15276
rect 1106 15208 1130 15264
rect 1186 15208 1254 15264
rect 1310 15208 1378 15264
rect 1434 15208 1502 15264
rect 1558 15208 1582 15264
rect 1106 15140 1582 15208
rect 1106 15084 1130 15140
rect 1186 15084 1254 15140
rect 1310 15084 1378 15140
rect 1434 15084 1502 15140
rect 1558 15084 1582 15140
rect 1106 15016 1582 15084
rect 1106 14960 1130 15016
rect 1186 14960 1254 15016
rect 1310 14960 1378 15016
rect 1434 14960 1502 15016
rect 1558 14960 1582 15016
rect 1106 14892 1582 14960
rect 1106 14836 1130 14892
rect 1186 14836 1254 14892
rect 1310 14836 1378 14892
rect 1434 14836 1502 14892
rect 1558 14836 1582 14892
rect 1106 14824 1582 14836
rect 85788 15264 86264 15276
rect 85788 15208 85812 15264
rect 85868 15208 85936 15264
rect 85992 15208 86060 15264
rect 86116 15208 86184 15264
rect 86240 15208 86264 15264
rect 85788 15140 86264 15208
rect 85788 15084 85812 15140
rect 85868 15084 85936 15140
rect 85992 15084 86060 15140
rect 86116 15084 86184 15140
rect 86240 15084 86264 15140
rect 85788 15016 86264 15084
rect 85788 14960 85812 15016
rect 85868 14960 85936 15016
rect 85992 14960 86060 15016
rect 86116 14960 86184 15016
rect 86240 14960 86264 15016
rect 85788 14892 86264 14960
rect 85788 14836 85812 14892
rect 85868 14836 85936 14892
rect 85992 14836 86060 14892
rect 86116 14836 86184 14892
rect 86240 14836 86264 14892
rect 85788 14824 86264 14836
rect 86588 14364 87064 14376
rect 86588 14308 86612 14364
rect 86668 14308 86736 14364
rect 86792 14308 86860 14364
rect 86916 14308 86984 14364
rect 87040 14308 87064 14364
rect 1906 14240 2382 14300
rect 1906 14184 1930 14240
rect 1986 14184 2054 14240
rect 2110 14184 2178 14240
rect 2234 14184 2302 14240
rect 2358 14184 2382 14240
rect 1906 14116 2382 14184
rect 1906 14060 1930 14116
rect 1986 14060 2054 14116
rect 2110 14060 2178 14116
rect 2234 14060 2302 14116
rect 2358 14060 2382 14116
rect 1906 14000 2382 14060
rect 86588 14240 87064 14308
rect 86588 14184 86612 14240
rect 86668 14184 86736 14240
rect 86792 14184 86860 14240
rect 86916 14184 86984 14240
rect 87040 14184 87064 14240
rect 86588 14116 87064 14184
rect 86588 14060 86612 14116
rect 86668 14060 86736 14116
rect 86792 14060 86860 14116
rect 86916 14060 86984 14116
rect 87040 14060 87064 14116
rect 86588 13992 87064 14060
rect 86588 13936 86612 13992
rect 86668 13936 86736 13992
rect 86792 13936 86860 13992
rect 86916 13936 86984 13992
rect 87040 13936 87064 13992
rect 86588 13924 87064 13936
rect 1106 13464 1582 13476
rect 1106 13408 1130 13464
rect 1186 13408 1254 13464
rect 1310 13408 1378 13464
rect 1434 13408 1502 13464
rect 1558 13408 1582 13464
rect 1106 13340 1582 13408
rect 1106 13284 1130 13340
rect 1186 13284 1254 13340
rect 1310 13284 1378 13340
rect 1434 13284 1502 13340
rect 1558 13284 1582 13340
rect 1106 13216 1582 13284
rect 1106 13160 1130 13216
rect 1186 13160 1254 13216
rect 1310 13160 1378 13216
rect 1434 13160 1502 13216
rect 1558 13160 1582 13216
rect 1106 13092 1582 13160
rect 1106 13036 1130 13092
rect 1186 13036 1254 13092
rect 1310 13036 1378 13092
rect 1434 13036 1502 13092
rect 1558 13036 1582 13092
rect 1106 13024 1582 13036
rect 85788 13464 86264 13476
rect 85788 13408 85812 13464
rect 85868 13408 85936 13464
rect 85992 13408 86060 13464
rect 86116 13408 86184 13464
rect 86240 13408 86264 13464
rect 85788 13340 86264 13408
rect 85788 13284 85812 13340
rect 85868 13284 85936 13340
rect 85992 13284 86060 13340
rect 86116 13284 86184 13340
rect 86240 13284 86264 13340
rect 85788 13216 86264 13284
rect 85788 13160 85812 13216
rect 85868 13160 85936 13216
rect 85992 13160 86060 13216
rect 86116 13160 86184 13216
rect 86240 13160 86264 13216
rect 85788 13092 86264 13160
rect 85788 13036 85812 13092
rect 85868 13036 85936 13092
rect 85992 13036 86060 13092
rect 86116 13036 86184 13092
rect 86240 13036 86264 13092
rect 85788 13024 86264 13036
rect 86588 12564 87064 12576
rect 86588 12508 86612 12564
rect 86668 12508 86736 12564
rect 86792 12508 86860 12564
rect 86916 12508 86984 12564
rect 87040 12508 87064 12564
rect 1906 12440 2382 12500
rect 1906 12384 1930 12440
rect 1986 12384 2054 12440
rect 2110 12384 2178 12440
rect 2234 12384 2302 12440
rect 2358 12384 2382 12440
rect 1906 12316 2382 12384
rect 1906 12260 1930 12316
rect 1986 12260 2054 12316
rect 2110 12260 2178 12316
rect 2234 12260 2302 12316
rect 2358 12260 2382 12316
rect 1906 12200 2382 12260
rect 86588 12440 87064 12508
rect 86588 12384 86612 12440
rect 86668 12384 86736 12440
rect 86792 12384 86860 12440
rect 86916 12384 86984 12440
rect 87040 12384 87064 12440
rect 86588 12316 87064 12384
rect 86588 12260 86612 12316
rect 86668 12260 86736 12316
rect 86792 12260 86860 12316
rect 86916 12260 86984 12316
rect 87040 12260 87064 12316
rect 86588 12192 87064 12260
rect 86588 12136 86612 12192
rect 86668 12136 86736 12192
rect 86792 12136 86860 12192
rect 86916 12136 86984 12192
rect 87040 12136 87064 12192
rect 86588 12124 87064 12136
rect 1106 11664 1582 11676
rect 1106 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1582 11664
rect 1106 11540 1582 11608
rect 1106 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1582 11540
rect 1106 11416 1582 11484
rect 1106 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1582 11416
rect 1106 11292 1582 11360
rect 1106 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1582 11292
rect 1106 11224 1582 11236
rect 85788 11664 86264 11676
rect 85788 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86264 11664
rect 85788 11540 86264 11608
rect 85788 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86264 11540
rect 85788 11416 86264 11484
rect 85788 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86264 11416
rect 85788 11292 86264 11360
rect 85788 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86264 11292
rect 85788 11224 86264 11236
rect 86588 10764 87064 10776
rect 86588 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87064 10764
rect 1906 10640 2382 10700
rect 1906 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2382 10640
rect 1906 10516 2382 10584
rect 1906 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2382 10516
rect 1906 10400 2382 10460
rect 86588 10640 87064 10708
rect 86588 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87064 10640
rect 86588 10516 87064 10584
rect 86588 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87064 10516
rect 86588 10392 87064 10460
rect 86588 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87064 10392
rect 86588 10324 87064 10336
rect 1106 9864 1582 9876
rect 1106 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1582 9864
rect 1106 9740 1582 9808
rect 1106 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1582 9740
rect 1106 9616 1582 9684
rect 1106 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1582 9616
rect 1106 9492 1582 9560
rect 1106 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1582 9492
rect 1106 9424 1582 9436
rect 85788 9864 86264 9876
rect 85788 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86264 9864
rect 85788 9740 86264 9808
rect 85788 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86264 9740
rect 85788 9616 86264 9684
rect 85788 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86264 9616
rect 85788 9492 86264 9560
rect 85788 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86264 9492
rect 85788 9424 86264 9436
rect 86588 8964 87064 8976
rect 86588 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87064 8964
rect 1906 8840 2382 8900
rect 1906 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2382 8840
rect 1906 8716 2382 8784
rect 1906 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2382 8716
rect 1906 8600 2382 8660
rect 86588 8840 87064 8908
rect 86588 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87064 8840
rect 86588 8716 87064 8784
rect 86588 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87064 8716
rect 86588 8592 87064 8660
rect 86588 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87064 8592
rect 86588 8524 87064 8536
rect 1106 8064 1582 8076
rect 1106 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1582 8064
rect 1106 7940 1582 8008
rect 1106 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1582 7940
rect 1106 7816 1582 7884
rect 1106 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1582 7816
rect 1106 7692 1582 7760
rect 1106 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1582 7692
rect 1106 7624 1582 7636
rect 85788 8064 86264 8076
rect 85788 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86264 8064
rect 85788 7940 86264 8008
rect 85788 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86264 7940
rect 85788 7816 86264 7884
rect 85788 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86264 7816
rect 85788 7692 86264 7760
rect 85788 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86264 7692
rect 85788 7624 86264 7636
rect 86588 7164 87064 7176
rect 86588 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87064 7164
rect 1906 7040 2382 7100
rect 1906 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2382 7040
rect 1906 6916 2382 6984
rect 1906 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2382 6916
rect 1906 6800 2382 6860
rect 86588 7040 87064 7108
rect 86588 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87064 7040
rect 86588 6916 87064 6984
rect 86588 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87064 6916
rect 86588 6792 87064 6860
rect 86588 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87064 6792
rect 86588 6724 87064 6736
rect 1106 6264 1582 6276
rect 1106 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1582 6264
rect 1106 6140 1582 6208
rect 1106 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1582 6140
rect 1106 6016 1582 6084
rect 1106 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1582 6016
rect 1106 5892 1582 5960
rect 1106 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1582 5892
rect 1106 5824 1582 5836
rect 85788 6264 86264 6276
rect 85788 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86264 6264
rect 85788 6140 86264 6208
rect 85788 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86264 6140
rect 85788 6016 86264 6084
rect 85788 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86264 6016
rect 85788 5892 86264 5960
rect 85788 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86264 5892
rect 85788 5824 86264 5836
rect 86588 5364 87064 5376
rect 86588 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87064 5364
rect 1906 5240 2382 5300
rect 1906 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2382 5240
rect 1906 5116 2382 5184
rect 1906 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2382 5116
rect 1906 5000 2382 5060
rect 86588 5240 87064 5308
rect 86588 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87064 5240
rect 86588 5116 87064 5184
rect 86588 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87064 5116
rect 86588 4992 87064 5060
rect 86588 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87064 4992
rect 86588 4924 87064 4936
rect 1106 4464 1582 4476
rect 1106 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1582 4464
rect 1106 4340 1582 4408
rect 1106 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1582 4340
rect 1106 4216 1582 4284
rect 1106 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1582 4216
rect 1106 4092 1582 4160
rect 1106 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1582 4092
rect 1106 4024 1582 4036
rect 85788 4464 86264 4476
rect 85788 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86264 4464
rect 85788 4340 86264 4408
rect 85788 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86264 4340
rect 85788 4216 86264 4284
rect 85788 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86264 4216
rect 85788 4092 86264 4160
rect 85788 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86264 4092
rect 85788 4024 86264 4036
rect 86588 3632 87064 3700
rect 86588 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87064 3632
rect 86588 3508 87064 3576
rect 1906 3440 2382 3500
rect 1906 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2382 3440
rect 1906 3316 2382 3384
rect 1906 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2382 3316
rect 1906 3200 2382 3260
rect 86588 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87064 3508
rect 86588 3384 87064 3452
rect 86588 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87064 3384
rect 86588 3260 87064 3328
rect 86588 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87064 3260
rect 86588 3136 87064 3204
<< via3 >>
rect 1930 66515 1986 66571
rect 2054 66515 2110 66571
rect 2178 66515 2234 66571
rect 2302 66515 2358 66571
rect 1930 66391 1986 66447
rect 2054 66391 2110 66447
rect 2178 66391 2234 66447
rect 2302 66391 2358 66447
rect 86550 66552 86606 66608
rect 86550 66428 86606 66484
rect 86550 66304 86606 66360
rect 86550 66180 86606 66236
rect 86674 66552 86730 66608
rect 86798 66552 86854 66608
rect 86922 66552 86978 66608
rect 87046 66552 87102 66608
rect 86674 66428 86730 66484
rect 86798 66428 86854 66484
rect 86922 66428 86978 66484
rect 87046 66428 87102 66484
rect 86674 66304 86730 66360
rect 86798 66304 86854 66360
rect 86922 66304 86978 66360
rect 87046 66304 87102 66360
rect 86674 66180 86730 66236
rect 86798 66180 86854 66236
rect 86922 66180 86978 66236
rect 87046 66180 87102 66236
rect 86550 66056 86606 66112
rect 86550 65932 86606 65988
rect 86550 65808 86606 65864
rect 1930 65676 1986 65732
rect 2054 65676 2110 65732
rect 2178 65676 2234 65732
rect 2302 65676 2358 65732
rect 86550 65684 86606 65740
rect 86674 66056 86730 66112
rect 86798 66056 86854 66112
rect 86922 66056 86978 66112
rect 87046 66056 87102 66112
rect 86674 65932 86730 65988
rect 86798 65932 86854 65988
rect 86922 65932 86978 65988
rect 87046 65932 87102 65988
rect 86674 65808 86730 65864
rect 86798 65808 86854 65864
rect 86922 65808 86978 65864
rect 87046 65808 87102 65864
rect 86674 65684 86730 65740
rect 86798 65684 86854 65740
rect 86922 65684 86978 65740
rect 87046 65684 87102 65740
rect 1930 65552 1986 65608
rect 2054 65552 2110 65608
rect 2178 65552 2234 65608
rect 2302 65552 2358 65608
rect 1930 65428 1986 65484
rect 2054 65428 2110 65484
rect 2178 65428 2234 65484
rect 2302 65428 2358 65484
rect 86550 65560 86606 65616
rect 86550 65436 86606 65492
rect 86674 65560 86730 65616
rect 86798 65560 86854 65616
rect 86922 65560 86978 65616
rect 87046 65560 87102 65616
rect 86674 65436 86730 65492
rect 86798 65436 86854 65492
rect 86922 65436 86978 65492
rect 87046 65436 87102 65492
rect 1930 63290 1986 63346
rect 2054 63290 2110 63346
rect 2178 63290 2234 63346
rect 2302 63290 2358 63346
rect 1930 63166 1986 63222
rect 2054 63166 2110 63222
rect 2178 63166 2234 63222
rect 2302 63166 2358 63222
rect 1930 63042 1986 63098
rect 2054 63042 2110 63098
rect 2178 63042 2234 63098
rect 2302 63042 2358 63098
rect 86550 63335 86606 63391
rect 86550 63211 86606 63267
rect 86550 63087 86606 63143
rect 86550 62963 86606 63019
rect 86674 63335 86730 63391
rect 86798 63335 86854 63391
rect 86922 63335 86978 63391
rect 87046 63335 87102 63391
rect 86674 63211 86730 63267
rect 86798 63211 86854 63267
rect 86922 63211 86978 63267
rect 87046 63211 87102 63267
rect 86674 63087 86730 63143
rect 86798 63087 86854 63143
rect 86922 63087 86978 63143
rect 87046 63087 87102 63143
rect 86674 62963 86730 63019
rect 86798 62963 86854 63019
rect 86922 62963 86978 63019
rect 87046 62963 87102 63019
rect 86550 62839 86606 62895
rect 86550 62715 86606 62771
rect 86550 62591 86606 62647
rect 86550 62467 86606 62523
rect 86674 62839 86730 62895
rect 86798 62839 86854 62895
rect 86922 62839 86978 62895
rect 87046 62839 87102 62895
rect 86674 62715 86730 62771
rect 86798 62715 86854 62771
rect 86922 62715 86978 62771
rect 87046 62715 87102 62771
rect 86674 62591 86730 62647
rect 86798 62591 86854 62647
rect 86922 62591 86978 62647
rect 87046 62591 87102 62647
rect 86674 62467 86730 62523
rect 86798 62467 86854 62523
rect 86922 62467 86978 62523
rect 87046 62467 87102 62523
rect 86550 62343 86606 62399
rect 86550 62219 86606 62275
rect 1930 62045 1986 62101
rect 2054 62045 2110 62101
rect 2178 62045 2234 62101
rect 2302 62045 2358 62101
rect 1930 61921 1986 61977
rect 2054 61921 2110 61977
rect 2178 61921 2234 61977
rect 2302 61921 2358 61977
rect 86550 62095 86606 62151
rect 86550 61971 86606 62027
rect 86674 62343 86730 62399
rect 86798 62343 86854 62399
rect 86922 62343 86978 62399
rect 87046 62343 87102 62399
rect 86674 62219 86730 62275
rect 86798 62219 86854 62275
rect 86922 62219 86978 62275
rect 87046 62219 87102 62275
rect 86674 62095 86730 62151
rect 86798 62095 86854 62151
rect 86922 62095 86978 62151
rect 87046 62095 87102 62151
rect 86674 61971 86730 62027
rect 86798 61971 86854 62027
rect 86922 61971 86978 62027
rect 87046 61971 87102 62027
rect 1930 61797 1986 61853
rect 2054 61797 2110 61853
rect 2178 61797 2234 61853
rect 2302 61797 2358 61853
rect 1930 61673 1986 61729
rect 2054 61673 2110 61729
rect 2178 61673 2234 61729
rect 2302 61673 2358 61729
rect 86550 61847 86606 61903
rect 86550 61723 86606 61779
rect 86550 61599 86606 61655
rect 86674 61847 86730 61903
rect 86798 61847 86854 61903
rect 86922 61847 86978 61903
rect 87046 61847 87102 61903
rect 86674 61723 86730 61779
rect 86798 61723 86854 61779
rect 86922 61723 86978 61779
rect 87046 61723 87102 61779
rect 86674 61599 86730 61655
rect 86798 61599 86854 61655
rect 86922 61599 86978 61655
rect 87046 61599 87102 61655
rect 85750 60935 85806 60991
rect 85750 60811 85806 60867
rect 85750 60687 85806 60743
rect 85750 60563 85806 60619
rect 85874 60935 85930 60991
rect 85998 60935 86054 60991
rect 86122 60935 86178 60991
rect 86246 60935 86302 60991
rect 85874 60811 85930 60867
rect 85998 60811 86054 60867
rect 86122 60811 86178 60867
rect 86246 60811 86302 60867
rect 85874 60687 85930 60743
rect 85998 60687 86054 60743
rect 86122 60687 86178 60743
rect 86246 60687 86302 60743
rect 85874 60563 85930 60619
rect 85998 60563 86054 60619
rect 86122 60563 86178 60619
rect 86246 60563 86302 60619
rect 85750 60439 85806 60495
rect 85750 60315 85806 60371
rect 85750 60191 85806 60247
rect 85750 60067 85806 60123
rect 85874 60439 85930 60495
rect 85998 60439 86054 60495
rect 86122 60439 86178 60495
rect 86246 60439 86302 60495
rect 85874 60315 85930 60371
rect 85998 60315 86054 60371
rect 86122 60315 86178 60371
rect 86246 60315 86302 60371
rect 85874 60191 85930 60247
rect 85998 60191 86054 60247
rect 86122 60191 86178 60247
rect 86246 60191 86302 60247
rect 85874 60067 85930 60123
rect 85998 60067 86054 60123
rect 86122 60067 86178 60123
rect 86246 60067 86302 60123
rect 85750 59943 85806 59999
rect 85750 59819 85806 59875
rect 85750 59695 85806 59751
rect 85874 59943 85930 59999
rect 85998 59943 86054 59999
rect 86122 59943 86178 59999
rect 86246 59943 86302 59999
rect 85874 59819 85930 59875
rect 85998 59819 86054 59875
rect 86122 59819 86178 59875
rect 86246 59819 86302 59875
rect 85874 59695 85930 59751
rect 85998 59695 86054 59751
rect 86122 59695 86178 59751
rect 86246 59695 86302 59751
rect 1068 57033 1124 57089
rect 1068 56909 1124 56965
rect 1068 56785 1124 56841
rect 1068 56661 1124 56717
rect 1068 56537 1124 56593
rect 1068 56413 1124 56469
rect 1068 56289 1124 56345
rect 1068 56165 1124 56221
rect 1068 56041 1124 56097
rect 1068 55917 1124 55973
rect 1068 55793 1124 55849
rect 1068 55669 1124 55725
rect 1068 55545 1124 55601
rect 1068 55421 1124 55477
rect 1068 55297 1124 55353
rect 1068 55173 1124 55229
rect 1068 55049 1124 55105
rect 1192 57033 1248 57089
rect 1316 57033 1372 57089
rect 1440 57033 1496 57089
rect 1564 57033 1620 57089
rect 1192 56909 1248 56965
rect 1316 56909 1372 56965
rect 1440 56909 1496 56965
rect 1564 56909 1620 56965
rect 1192 56785 1248 56841
rect 1316 56785 1372 56841
rect 1440 56785 1496 56841
rect 1564 56785 1620 56841
rect 1192 56661 1248 56717
rect 1316 56661 1372 56717
rect 1440 56661 1496 56717
rect 1564 56661 1620 56717
rect 1192 56537 1248 56593
rect 1316 56537 1372 56593
rect 1440 56537 1496 56593
rect 1564 56537 1620 56593
rect 1192 56413 1248 56469
rect 1316 56413 1372 56469
rect 1440 56413 1496 56469
rect 1564 56413 1620 56469
rect 1192 56289 1248 56345
rect 1316 56289 1372 56345
rect 1440 56289 1496 56345
rect 1564 56289 1620 56345
rect 1192 56165 1248 56221
rect 1316 56165 1372 56221
rect 1440 56165 1496 56221
rect 1564 56165 1620 56221
rect 1192 56041 1248 56097
rect 1316 56041 1372 56097
rect 1440 56041 1496 56097
rect 1564 56041 1620 56097
rect 1192 55917 1248 55973
rect 1316 55917 1372 55973
rect 1440 55917 1496 55973
rect 1564 55917 1620 55973
rect 1192 55793 1248 55849
rect 1316 55793 1372 55849
rect 1440 55793 1496 55849
rect 1564 55793 1620 55849
rect 1192 55669 1248 55725
rect 1316 55669 1372 55725
rect 1440 55669 1496 55725
rect 1564 55669 1620 55725
rect 1192 55545 1248 55601
rect 1316 55545 1372 55601
rect 1440 55545 1496 55601
rect 1564 55545 1620 55601
rect 1192 55421 1248 55477
rect 1316 55421 1372 55477
rect 1440 55421 1496 55477
rect 1564 55421 1620 55477
rect 1192 55297 1248 55353
rect 1316 55297 1372 55353
rect 1440 55297 1496 55353
rect 1564 55297 1620 55353
rect 1192 55173 1248 55229
rect 1316 55173 1372 55229
rect 1440 55173 1496 55229
rect 1564 55173 1620 55229
rect 1192 55049 1248 55105
rect 1316 55049 1372 55105
rect 1440 55049 1496 55105
rect 1564 55049 1620 55105
rect 85750 57033 85806 57089
rect 85750 56909 85806 56965
rect 85750 56785 85806 56841
rect 85750 56661 85806 56717
rect 85750 56537 85806 56593
rect 85750 56413 85806 56469
rect 85750 56289 85806 56345
rect 85750 56165 85806 56221
rect 85750 56041 85806 56097
rect 85750 55917 85806 55973
rect 85750 55793 85806 55849
rect 85750 55669 85806 55725
rect 85750 55545 85806 55601
rect 85750 55421 85806 55477
rect 85750 55297 85806 55353
rect 85750 55173 85806 55229
rect 85750 55049 85806 55105
rect 85874 57033 85930 57089
rect 85998 57033 86054 57089
rect 86122 57033 86178 57089
rect 86246 57033 86302 57089
rect 85874 56909 85930 56965
rect 85998 56909 86054 56965
rect 86122 56909 86178 56965
rect 86246 56909 86302 56965
rect 85874 56785 85930 56841
rect 85998 56785 86054 56841
rect 86122 56785 86178 56841
rect 86246 56785 86302 56841
rect 85874 56661 85930 56717
rect 85998 56661 86054 56717
rect 86122 56661 86178 56717
rect 86246 56661 86302 56717
rect 85874 56537 85930 56593
rect 85998 56537 86054 56593
rect 86122 56537 86178 56593
rect 86246 56537 86302 56593
rect 85874 56413 85930 56469
rect 85998 56413 86054 56469
rect 86122 56413 86178 56469
rect 86246 56413 86302 56469
rect 85874 56289 85930 56345
rect 85998 56289 86054 56345
rect 86122 56289 86178 56345
rect 86246 56289 86302 56345
rect 85874 56165 85930 56221
rect 85998 56165 86054 56221
rect 86122 56165 86178 56221
rect 86246 56165 86302 56221
rect 85874 56041 85930 56097
rect 85998 56041 86054 56097
rect 86122 56041 86178 56097
rect 86246 56041 86302 56097
rect 85874 55917 85930 55973
rect 85998 55917 86054 55973
rect 86122 55917 86178 55973
rect 86246 55917 86302 55973
rect 85874 55793 85930 55849
rect 85998 55793 86054 55849
rect 86122 55793 86178 55849
rect 86246 55793 86302 55849
rect 85874 55669 85930 55725
rect 85998 55669 86054 55725
rect 86122 55669 86178 55725
rect 86246 55669 86302 55725
rect 85874 55545 85930 55601
rect 85998 55545 86054 55601
rect 86122 55545 86178 55601
rect 86246 55545 86302 55601
rect 85874 55421 85930 55477
rect 85998 55421 86054 55477
rect 86122 55421 86178 55477
rect 86246 55421 86302 55477
rect 85874 55297 85930 55353
rect 85998 55297 86054 55353
rect 86122 55297 86178 55353
rect 86246 55297 86302 55353
rect 85874 55173 85930 55229
rect 85998 55173 86054 55229
rect 86122 55173 86178 55229
rect 86246 55173 86302 55229
rect 85874 55049 85930 55105
rect 85998 55049 86054 55105
rect 86122 55049 86178 55105
rect 86246 55049 86302 55105
rect 1868 54731 1924 54787
rect 1868 54607 1924 54663
rect 1868 54483 1924 54539
rect 1868 54359 1924 54415
rect 1868 54235 1924 54291
rect 1868 54111 1924 54167
rect 1868 53987 1924 54043
rect 1868 53863 1924 53919
rect 1868 53739 1924 53795
rect 1868 53615 1924 53671
rect 1868 53491 1924 53547
rect 1868 53367 1924 53423
rect 1868 53243 1924 53299
rect 1868 53119 1924 53175
rect 1868 52995 1924 53051
rect 1868 52871 1924 52927
rect 1868 52747 1924 52803
rect 1868 52623 1924 52679
rect 1868 52499 1924 52555
rect 1868 52375 1924 52431
rect 1868 52251 1924 52307
rect 1868 52127 1924 52183
rect 1868 52003 1924 52059
rect 1868 51879 1924 51935
rect 1868 51755 1924 51811
rect 1868 51631 1924 51687
rect 1868 51507 1924 51563
rect 1992 54731 2048 54787
rect 2116 54731 2172 54787
rect 2240 54731 2296 54787
rect 2364 54731 2420 54787
rect 1992 54607 2048 54663
rect 2116 54607 2172 54663
rect 2240 54607 2296 54663
rect 2364 54607 2420 54663
rect 1992 54483 2048 54539
rect 2116 54483 2172 54539
rect 2240 54483 2296 54539
rect 2364 54483 2420 54539
rect 1992 54359 2048 54415
rect 2116 54359 2172 54415
rect 2240 54359 2296 54415
rect 2364 54359 2420 54415
rect 1992 54235 2048 54291
rect 2116 54235 2172 54291
rect 2240 54235 2296 54291
rect 2364 54235 2420 54291
rect 1992 54111 2048 54167
rect 2116 54111 2172 54167
rect 2240 54111 2296 54167
rect 2364 54111 2420 54167
rect 1992 53987 2048 54043
rect 2116 53987 2172 54043
rect 2240 53987 2296 54043
rect 2364 53987 2420 54043
rect 1992 53863 2048 53919
rect 2116 53863 2172 53919
rect 2240 53863 2296 53919
rect 2364 53863 2420 53919
rect 1992 53739 2048 53795
rect 2116 53739 2172 53795
rect 2240 53739 2296 53795
rect 2364 53739 2420 53795
rect 1992 53615 2048 53671
rect 2116 53615 2172 53671
rect 2240 53615 2296 53671
rect 2364 53615 2420 53671
rect 1992 53491 2048 53547
rect 2116 53491 2172 53547
rect 2240 53491 2296 53547
rect 2364 53491 2420 53547
rect 1992 53367 2048 53423
rect 2116 53367 2172 53423
rect 2240 53367 2296 53423
rect 2364 53367 2420 53423
rect 1992 53243 2048 53299
rect 2116 53243 2172 53299
rect 2240 53243 2296 53299
rect 2364 53243 2420 53299
rect 1992 53119 2048 53175
rect 2116 53119 2172 53175
rect 2240 53119 2296 53175
rect 2364 53119 2420 53175
rect 1992 52995 2048 53051
rect 2116 52995 2172 53051
rect 2240 52995 2296 53051
rect 2364 52995 2420 53051
rect 1992 52871 2048 52927
rect 2116 52871 2172 52927
rect 2240 52871 2296 52927
rect 2364 52871 2420 52927
rect 1992 52747 2048 52803
rect 2116 52747 2172 52803
rect 2240 52747 2296 52803
rect 2364 52747 2420 52803
rect 1992 52623 2048 52679
rect 2116 52623 2172 52679
rect 2240 52623 2296 52679
rect 2364 52623 2420 52679
rect 1992 52499 2048 52555
rect 2116 52499 2172 52555
rect 2240 52499 2296 52555
rect 2364 52499 2420 52555
rect 1992 52375 2048 52431
rect 2116 52375 2172 52431
rect 2240 52375 2296 52431
rect 2364 52375 2420 52431
rect 1992 52251 2048 52307
rect 2116 52251 2172 52307
rect 2240 52251 2296 52307
rect 2364 52251 2420 52307
rect 1992 52127 2048 52183
rect 2116 52127 2172 52183
rect 2240 52127 2296 52183
rect 2364 52127 2420 52183
rect 1992 52003 2048 52059
rect 2116 52003 2172 52059
rect 2240 52003 2296 52059
rect 2364 52003 2420 52059
rect 1992 51879 2048 51935
rect 2116 51879 2172 51935
rect 2240 51879 2296 51935
rect 2364 51879 2420 51935
rect 1992 51755 2048 51811
rect 2116 51755 2172 51811
rect 2240 51755 2296 51811
rect 2364 51755 2420 51811
rect 1992 51631 2048 51687
rect 2116 51631 2172 51687
rect 2240 51631 2296 51687
rect 2364 51631 2420 51687
rect 1992 51507 2048 51563
rect 2116 51507 2172 51563
rect 2240 51507 2296 51563
rect 2364 51507 2420 51563
rect 86550 54731 86606 54787
rect 86550 54607 86606 54663
rect 86550 54483 86606 54539
rect 86550 54359 86606 54415
rect 86550 54235 86606 54291
rect 86550 54111 86606 54167
rect 86550 53987 86606 54043
rect 86550 53863 86606 53919
rect 86550 53739 86606 53795
rect 86550 53615 86606 53671
rect 86550 53491 86606 53547
rect 86550 53367 86606 53423
rect 86550 53243 86606 53299
rect 86550 53119 86606 53175
rect 86550 52995 86606 53051
rect 86550 52871 86606 52927
rect 86550 52747 86606 52803
rect 86550 52623 86606 52679
rect 86550 52499 86606 52555
rect 86550 52375 86606 52431
rect 86550 52251 86606 52307
rect 86550 52127 86606 52183
rect 86550 52003 86606 52059
rect 86550 51879 86606 51935
rect 86550 51755 86606 51811
rect 86550 51631 86606 51687
rect 86550 51507 86606 51563
rect 86674 54731 86730 54787
rect 86798 54731 86854 54787
rect 86922 54731 86978 54787
rect 87046 54731 87102 54787
rect 86674 54607 86730 54663
rect 86798 54607 86854 54663
rect 86922 54607 86978 54663
rect 87046 54607 87102 54663
rect 86674 54483 86730 54539
rect 86798 54483 86854 54539
rect 86922 54483 86978 54539
rect 87046 54483 87102 54539
rect 86674 54359 86730 54415
rect 86798 54359 86854 54415
rect 86922 54359 86978 54415
rect 87046 54359 87102 54415
rect 86674 54235 86730 54291
rect 86798 54235 86854 54291
rect 86922 54235 86978 54291
rect 87046 54235 87102 54291
rect 86674 54111 86730 54167
rect 86798 54111 86854 54167
rect 86922 54111 86978 54167
rect 87046 54111 87102 54167
rect 86674 53987 86730 54043
rect 86798 53987 86854 54043
rect 86922 53987 86978 54043
rect 87046 53987 87102 54043
rect 86674 53863 86730 53919
rect 86798 53863 86854 53919
rect 86922 53863 86978 53919
rect 87046 53863 87102 53919
rect 86674 53739 86730 53795
rect 86798 53739 86854 53795
rect 86922 53739 86978 53795
rect 87046 53739 87102 53795
rect 86674 53615 86730 53671
rect 86798 53615 86854 53671
rect 86922 53615 86978 53671
rect 87046 53615 87102 53671
rect 86674 53491 86730 53547
rect 86798 53491 86854 53547
rect 86922 53491 86978 53547
rect 87046 53491 87102 53547
rect 86674 53367 86730 53423
rect 86798 53367 86854 53423
rect 86922 53367 86978 53423
rect 87046 53367 87102 53423
rect 86674 53243 86730 53299
rect 86798 53243 86854 53299
rect 86922 53243 86978 53299
rect 87046 53243 87102 53299
rect 86674 53119 86730 53175
rect 86798 53119 86854 53175
rect 86922 53119 86978 53175
rect 87046 53119 87102 53175
rect 86674 52995 86730 53051
rect 86798 52995 86854 53051
rect 86922 52995 86978 53051
rect 87046 52995 87102 53051
rect 86674 52871 86730 52927
rect 86798 52871 86854 52927
rect 86922 52871 86978 52927
rect 87046 52871 87102 52927
rect 86674 52747 86730 52803
rect 86798 52747 86854 52803
rect 86922 52747 86978 52803
rect 87046 52747 87102 52803
rect 86674 52623 86730 52679
rect 86798 52623 86854 52679
rect 86922 52623 86978 52679
rect 87046 52623 87102 52679
rect 86674 52499 86730 52555
rect 86798 52499 86854 52555
rect 86922 52499 86978 52555
rect 87046 52499 87102 52555
rect 86674 52375 86730 52431
rect 86798 52375 86854 52431
rect 86922 52375 86978 52431
rect 87046 52375 87102 52431
rect 86674 52251 86730 52307
rect 86798 52251 86854 52307
rect 86922 52251 86978 52307
rect 87046 52251 87102 52307
rect 86674 52127 86730 52183
rect 86798 52127 86854 52183
rect 86922 52127 86978 52183
rect 87046 52127 87102 52183
rect 86674 52003 86730 52059
rect 86798 52003 86854 52059
rect 86922 52003 86978 52059
rect 87046 52003 87102 52059
rect 86674 51879 86730 51935
rect 86798 51879 86854 51935
rect 86922 51879 86978 51935
rect 87046 51879 87102 51935
rect 86674 51755 86730 51811
rect 86798 51755 86854 51811
rect 86922 51755 86978 51811
rect 87046 51755 87102 51811
rect 86674 51631 86730 51687
rect 86798 51631 86854 51687
rect 86922 51631 86978 51687
rect 87046 51631 87102 51687
rect 86674 51507 86730 51563
rect 86798 51507 86854 51563
rect 86922 51507 86978 51563
rect 87046 51507 87102 51563
rect 86550 47800 86606 47856
rect 86550 47676 86606 47732
rect 86550 47552 86606 47608
rect 86550 47428 86606 47484
rect 86550 47304 86606 47360
rect 86550 47180 86606 47236
rect 86550 47056 86606 47112
rect 86550 46932 86606 46988
rect 86674 47800 86730 47856
rect 86798 47800 86854 47856
rect 86922 47800 86978 47856
rect 87046 47800 87102 47856
rect 86674 47676 86730 47732
rect 86798 47676 86854 47732
rect 86922 47676 86978 47732
rect 87046 47676 87102 47732
rect 86674 47552 86730 47608
rect 86798 47552 86854 47608
rect 86922 47552 86978 47608
rect 87046 47552 87102 47608
rect 86674 47428 86730 47484
rect 86798 47428 86854 47484
rect 86922 47428 86978 47484
rect 87046 47428 87102 47484
rect 86674 47304 86730 47360
rect 86798 47304 86854 47360
rect 86922 47304 86978 47360
rect 87046 47304 87102 47360
rect 86674 47180 86730 47236
rect 86798 47180 86854 47236
rect 86922 47180 86978 47236
rect 87046 47180 87102 47236
rect 86674 47056 86730 47112
rect 86798 47056 86854 47112
rect 86922 47056 86978 47112
rect 87046 47056 87102 47112
rect 86674 46932 86730 46988
rect 86798 46932 86854 46988
rect 86922 46932 86978 46988
rect 87046 46932 87102 46988
rect 1068 46144 1124 46200
rect 1068 46020 1124 46076
rect 1068 45896 1124 45952
rect 1068 45772 1124 45828
rect 1068 45648 1124 45704
rect 1068 45524 1124 45580
rect 1068 45400 1124 45456
rect 1068 45276 1124 45332
rect 1192 46144 1248 46200
rect 1316 46144 1372 46200
rect 1440 46144 1496 46200
rect 1564 46144 1620 46200
rect 1192 46020 1248 46076
rect 1316 46020 1372 46076
rect 1440 46020 1496 46076
rect 1564 46020 1620 46076
rect 1192 45896 1248 45952
rect 1316 45896 1372 45952
rect 1440 45896 1496 45952
rect 1564 45896 1620 45952
rect 1192 45772 1248 45828
rect 1316 45772 1372 45828
rect 1440 45772 1496 45828
rect 1564 45772 1620 45828
rect 1192 45648 1248 45704
rect 1316 45648 1372 45704
rect 1440 45648 1496 45704
rect 1564 45648 1620 45704
rect 1192 45524 1248 45580
rect 1316 45524 1372 45580
rect 1440 45524 1496 45580
rect 1564 45524 1620 45580
rect 1192 45400 1248 45456
rect 1316 45400 1372 45456
rect 1440 45400 1496 45456
rect 1564 45400 1620 45456
rect 1192 45276 1248 45332
rect 1316 45276 1372 45332
rect 1440 45276 1496 45332
rect 1564 45276 1620 45332
rect 85750 46144 85806 46200
rect 85750 46020 85806 46076
rect 85750 45896 85806 45952
rect 85750 45772 85806 45828
rect 85750 45648 85806 45704
rect 85750 45524 85806 45580
rect 85750 45400 85806 45456
rect 85750 45276 85806 45332
rect 85874 46144 85930 46200
rect 85998 46144 86054 46200
rect 86122 46144 86178 46200
rect 86246 46144 86302 46200
rect 85874 46020 85930 46076
rect 85998 46020 86054 46076
rect 86122 46020 86178 46076
rect 86246 46020 86302 46076
rect 85874 45896 85930 45952
rect 85998 45896 86054 45952
rect 86122 45896 86178 45952
rect 86246 45896 86302 45952
rect 85874 45772 85930 45828
rect 85998 45772 86054 45828
rect 86122 45772 86178 45828
rect 86246 45772 86302 45828
rect 85874 45648 85930 45704
rect 85998 45648 86054 45704
rect 86122 45648 86178 45704
rect 86246 45648 86302 45704
rect 85874 45524 85930 45580
rect 85998 45524 86054 45580
rect 86122 45524 86178 45580
rect 86246 45524 86302 45580
rect 85874 45400 85930 45456
rect 85998 45400 86054 45456
rect 86122 45400 86178 45456
rect 86246 45400 86302 45456
rect 85874 45276 85930 45332
rect 85998 45276 86054 45332
rect 86122 45276 86178 45332
rect 86246 45276 86302 45332
rect 1930 34558 1986 34614
rect 2054 34558 2110 34614
rect 2178 34558 2234 34614
rect 2302 34558 2358 34614
rect 1930 34434 1986 34490
rect 2054 34434 2110 34490
rect 2178 34434 2234 34490
rect 2302 34434 2358 34490
rect 1930 34310 1986 34366
rect 2054 34310 2110 34366
rect 2178 34310 2234 34366
rect 2302 34310 2358 34366
rect 1930 34186 1986 34242
rect 2054 34186 2110 34242
rect 2178 34186 2234 34242
rect 2302 34186 2358 34242
rect 86612 34403 86668 34459
rect 86736 34403 86792 34459
rect 86860 34403 86916 34459
rect 86984 34403 87040 34459
rect 86612 34279 86668 34335
rect 86736 34279 86792 34335
rect 86860 34279 86916 34335
rect 86984 34279 87040 34335
rect 86612 34155 86668 34211
rect 86736 34155 86792 34211
rect 86860 34155 86916 34211
rect 86984 34155 87040 34211
rect 86612 34031 86668 34087
rect 86736 34031 86792 34087
rect 86860 34031 86916 34087
rect 86984 34031 87040 34087
rect 1130 33208 1186 33264
rect 1254 33208 1310 33264
rect 1378 33208 1434 33264
rect 1502 33208 1558 33264
rect 1130 33084 1186 33140
rect 1254 33084 1310 33140
rect 1378 33084 1434 33140
rect 1502 33084 1558 33140
rect 1130 32960 1186 33016
rect 1254 32960 1310 33016
rect 1378 32960 1434 33016
rect 1502 32960 1558 33016
rect 1130 32836 1186 32892
rect 1254 32836 1310 32892
rect 1378 32836 1434 32892
rect 1502 32836 1558 32892
rect 85812 33208 85868 33264
rect 85936 33208 85992 33264
rect 86060 33208 86116 33264
rect 86184 33208 86240 33264
rect 85812 33084 85868 33140
rect 85936 33084 85992 33140
rect 86060 33084 86116 33140
rect 86184 33084 86240 33140
rect 85812 32960 85868 33016
rect 85936 32960 85992 33016
rect 86060 32960 86116 33016
rect 86184 32960 86240 33016
rect 85812 32836 85868 32892
rect 85936 32836 85992 32892
rect 86060 32836 86116 32892
rect 86184 32836 86240 32892
rect 86612 32308 86668 32364
rect 86736 32308 86792 32364
rect 86860 32308 86916 32364
rect 86984 32308 87040 32364
rect 1930 32184 1986 32240
rect 2054 32184 2110 32240
rect 2178 32184 2234 32240
rect 2302 32184 2358 32240
rect 1930 32060 1986 32116
rect 2054 32060 2110 32116
rect 2178 32060 2234 32116
rect 2302 32060 2358 32116
rect 86612 32184 86668 32240
rect 86736 32184 86792 32240
rect 86860 32184 86916 32240
rect 86984 32184 87040 32240
rect 86612 32060 86668 32116
rect 86736 32060 86792 32116
rect 86860 32060 86916 32116
rect 86984 32060 87040 32116
rect 86612 31936 86668 31992
rect 86736 31936 86792 31992
rect 86860 31936 86916 31992
rect 86984 31936 87040 31992
rect 1130 31408 1186 31464
rect 1254 31408 1310 31464
rect 1378 31408 1434 31464
rect 1502 31408 1558 31464
rect 1130 31284 1186 31340
rect 1254 31284 1310 31340
rect 1378 31284 1434 31340
rect 1502 31284 1558 31340
rect 1130 31160 1186 31216
rect 1254 31160 1310 31216
rect 1378 31160 1434 31216
rect 1502 31160 1558 31216
rect 1130 31036 1186 31092
rect 1254 31036 1310 31092
rect 1378 31036 1434 31092
rect 1502 31036 1558 31092
rect 85812 31408 85868 31464
rect 85936 31408 85992 31464
rect 86060 31408 86116 31464
rect 86184 31408 86240 31464
rect 85812 31284 85868 31340
rect 85936 31284 85992 31340
rect 86060 31284 86116 31340
rect 86184 31284 86240 31340
rect 85812 31160 85868 31216
rect 85936 31160 85992 31216
rect 86060 31160 86116 31216
rect 86184 31160 86240 31216
rect 85812 31036 85868 31092
rect 85936 31036 85992 31092
rect 86060 31036 86116 31092
rect 86184 31036 86240 31092
rect 86612 30508 86668 30564
rect 86736 30508 86792 30564
rect 86860 30508 86916 30564
rect 86984 30508 87040 30564
rect 1930 30384 1986 30440
rect 2054 30384 2110 30440
rect 2178 30384 2234 30440
rect 2302 30384 2358 30440
rect 1930 30260 1986 30316
rect 2054 30260 2110 30316
rect 2178 30260 2234 30316
rect 2302 30260 2358 30316
rect 86612 30384 86668 30440
rect 86736 30384 86792 30440
rect 86860 30384 86916 30440
rect 86984 30384 87040 30440
rect 86612 30260 86668 30316
rect 86736 30260 86792 30316
rect 86860 30260 86916 30316
rect 86984 30260 87040 30316
rect 86612 30136 86668 30192
rect 86736 30136 86792 30192
rect 86860 30136 86916 30192
rect 86984 30136 87040 30192
rect 1130 29608 1186 29664
rect 1254 29608 1310 29664
rect 1378 29608 1434 29664
rect 1502 29608 1558 29664
rect 1130 29484 1186 29540
rect 1254 29484 1310 29540
rect 1378 29484 1434 29540
rect 1502 29484 1558 29540
rect 1130 29360 1186 29416
rect 1254 29360 1310 29416
rect 1378 29360 1434 29416
rect 1502 29360 1558 29416
rect 1130 29236 1186 29292
rect 1254 29236 1310 29292
rect 1378 29236 1434 29292
rect 1502 29236 1558 29292
rect 85812 29608 85868 29664
rect 85936 29608 85992 29664
rect 86060 29608 86116 29664
rect 86184 29608 86240 29664
rect 85812 29484 85868 29540
rect 85936 29484 85992 29540
rect 86060 29484 86116 29540
rect 86184 29484 86240 29540
rect 85812 29360 85868 29416
rect 85936 29360 85992 29416
rect 86060 29360 86116 29416
rect 86184 29360 86240 29416
rect 85812 29236 85868 29292
rect 85936 29236 85992 29292
rect 86060 29236 86116 29292
rect 86184 29236 86240 29292
rect 86612 28708 86668 28764
rect 86736 28708 86792 28764
rect 86860 28708 86916 28764
rect 86984 28708 87040 28764
rect 1930 28584 1986 28640
rect 2054 28584 2110 28640
rect 2178 28584 2234 28640
rect 2302 28584 2358 28640
rect 1930 28460 1986 28516
rect 2054 28460 2110 28516
rect 2178 28460 2234 28516
rect 2302 28460 2358 28516
rect 86612 28584 86668 28640
rect 86736 28584 86792 28640
rect 86860 28584 86916 28640
rect 86984 28584 87040 28640
rect 86612 28460 86668 28516
rect 86736 28460 86792 28516
rect 86860 28460 86916 28516
rect 86984 28460 87040 28516
rect 86612 28336 86668 28392
rect 86736 28336 86792 28392
rect 86860 28336 86916 28392
rect 86984 28336 87040 28392
rect 1130 27808 1186 27864
rect 1254 27808 1310 27864
rect 1378 27808 1434 27864
rect 1502 27808 1558 27864
rect 1130 27684 1186 27740
rect 1254 27684 1310 27740
rect 1378 27684 1434 27740
rect 1502 27684 1558 27740
rect 1130 27560 1186 27616
rect 1254 27560 1310 27616
rect 1378 27560 1434 27616
rect 1502 27560 1558 27616
rect 1130 27436 1186 27492
rect 1254 27436 1310 27492
rect 1378 27436 1434 27492
rect 1502 27436 1558 27492
rect 85812 27808 85868 27864
rect 85936 27808 85992 27864
rect 86060 27808 86116 27864
rect 86184 27808 86240 27864
rect 85812 27684 85868 27740
rect 85936 27684 85992 27740
rect 86060 27684 86116 27740
rect 86184 27684 86240 27740
rect 85812 27560 85868 27616
rect 85936 27560 85992 27616
rect 86060 27560 86116 27616
rect 86184 27560 86240 27616
rect 85812 27436 85868 27492
rect 85936 27436 85992 27492
rect 86060 27436 86116 27492
rect 86184 27436 86240 27492
rect 86612 26908 86668 26964
rect 86736 26908 86792 26964
rect 86860 26908 86916 26964
rect 86984 26908 87040 26964
rect 1930 26784 1986 26840
rect 2054 26784 2110 26840
rect 2178 26784 2234 26840
rect 2302 26784 2358 26840
rect 1930 26660 1986 26716
rect 2054 26660 2110 26716
rect 2178 26660 2234 26716
rect 2302 26660 2358 26716
rect 86612 26784 86668 26840
rect 86736 26784 86792 26840
rect 86860 26784 86916 26840
rect 86984 26784 87040 26840
rect 86612 26660 86668 26716
rect 86736 26660 86792 26716
rect 86860 26660 86916 26716
rect 86984 26660 87040 26716
rect 86612 26536 86668 26592
rect 86736 26536 86792 26592
rect 86860 26536 86916 26592
rect 86984 26536 87040 26592
rect 1130 26008 1186 26064
rect 1254 26008 1310 26064
rect 1378 26008 1434 26064
rect 1502 26008 1558 26064
rect 1130 25884 1186 25940
rect 1254 25884 1310 25940
rect 1378 25884 1434 25940
rect 1502 25884 1558 25940
rect 1130 25760 1186 25816
rect 1254 25760 1310 25816
rect 1378 25760 1434 25816
rect 1502 25760 1558 25816
rect 1130 25636 1186 25692
rect 1254 25636 1310 25692
rect 1378 25636 1434 25692
rect 1502 25636 1558 25692
rect 85812 26008 85868 26064
rect 85936 26008 85992 26064
rect 86060 26008 86116 26064
rect 86184 26008 86240 26064
rect 85812 25884 85868 25940
rect 85936 25884 85992 25940
rect 86060 25884 86116 25940
rect 86184 25884 86240 25940
rect 85812 25760 85868 25816
rect 85936 25760 85992 25816
rect 86060 25760 86116 25816
rect 86184 25760 86240 25816
rect 85812 25636 85868 25692
rect 85936 25636 85992 25692
rect 86060 25636 86116 25692
rect 86184 25636 86240 25692
rect 86612 25108 86668 25164
rect 86736 25108 86792 25164
rect 86860 25108 86916 25164
rect 86984 25108 87040 25164
rect 1930 24984 1986 25040
rect 2054 24984 2110 25040
rect 2178 24984 2234 25040
rect 2302 24984 2358 25040
rect 1930 24860 1986 24916
rect 2054 24860 2110 24916
rect 2178 24860 2234 24916
rect 2302 24860 2358 24916
rect 86612 24984 86668 25040
rect 86736 24984 86792 25040
rect 86860 24984 86916 25040
rect 86984 24984 87040 25040
rect 86612 24860 86668 24916
rect 86736 24860 86792 24916
rect 86860 24860 86916 24916
rect 86984 24860 87040 24916
rect 86612 24736 86668 24792
rect 86736 24736 86792 24792
rect 86860 24736 86916 24792
rect 86984 24736 87040 24792
rect 1130 24208 1186 24264
rect 1254 24208 1310 24264
rect 1378 24208 1434 24264
rect 1502 24208 1558 24264
rect 1130 24084 1186 24140
rect 1254 24084 1310 24140
rect 1378 24084 1434 24140
rect 1502 24084 1558 24140
rect 1130 23960 1186 24016
rect 1254 23960 1310 24016
rect 1378 23960 1434 24016
rect 1502 23960 1558 24016
rect 1130 23836 1186 23892
rect 1254 23836 1310 23892
rect 1378 23836 1434 23892
rect 1502 23836 1558 23892
rect 85812 24208 85868 24264
rect 85936 24208 85992 24264
rect 86060 24208 86116 24264
rect 86184 24208 86240 24264
rect 85812 24084 85868 24140
rect 85936 24084 85992 24140
rect 86060 24084 86116 24140
rect 86184 24084 86240 24140
rect 85812 23960 85868 24016
rect 85936 23960 85992 24016
rect 86060 23960 86116 24016
rect 86184 23960 86240 24016
rect 85812 23836 85868 23892
rect 85936 23836 85992 23892
rect 86060 23836 86116 23892
rect 86184 23836 86240 23892
rect 86612 23308 86668 23364
rect 86736 23308 86792 23364
rect 86860 23308 86916 23364
rect 86984 23308 87040 23364
rect 1930 23184 1986 23240
rect 2054 23184 2110 23240
rect 2178 23184 2234 23240
rect 2302 23184 2358 23240
rect 1930 23060 1986 23116
rect 2054 23060 2110 23116
rect 2178 23060 2234 23116
rect 2302 23060 2358 23116
rect 86612 23184 86668 23240
rect 86736 23184 86792 23240
rect 86860 23184 86916 23240
rect 86984 23184 87040 23240
rect 86612 23060 86668 23116
rect 86736 23060 86792 23116
rect 86860 23060 86916 23116
rect 86984 23060 87040 23116
rect 86612 22936 86668 22992
rect 86736 22936 86792 22992
rect 86860 22936 86916 22992
rect 86984 22936 87040 22992
rect 1130 22408 1186 22464
rect 1254 22408 1310 22464
rect 1378 22408 1434 22464
rect 1502 22408 1558 22464
rect 1130 22284 1186 22340
rect 1254 22284 1310 22340
rect 1378 22284 1434 22340
rect 1502 22284 1558 22340
rect 1130 22160 1186 22216
rect 1254 22160 1310 22216
rect 1378 22160 1434 22216
rect 1502 22160 1558 22216
rect 1130 22036 1186 22092
rect 1254 22036 1310 22092
rect 1378 22036 1434 22092
rect 1502 22036 1558 22092
rect 85812 22408 85868 22464
rect 85936 22408 85992 22464
rect 86060 22408 86116 22464
rect 86184 22408 86240 22464
rect 85812 22284 85868 22340
rect 85936 22284 85992 22340
rect 86060 22284 86116 22340
rect 86184 22284 86240 22340
rect 85812 22160 85868 22216
rect 85936 22160 85992 22216
rect 86060 22160 86116 22216
rect 86184 22160 86240 22216
rect 85812 22036 85868 22092
rect 85936 22036 85992 22092
rect 86060 22036 86116 22092
rect 86184 22036 86240 22092
rect 86612 21508 86668 21564
rect 86736 21508 86792 21564
rect 86860 21508 86916 21564
rect 86984 21508 87040 21564
rect 1930 21384 1986 21440
rect 2054 21384 2110 21440
rect 2178 21384 2234 21440
rect 2302 21384 2358 21440
rect 1930 21260 1986 21316
rect 2054 21260 2110 21316
rect 2178 21260 2234 21316
rect 2302 21260 2358 21316
rect 86612 21384 86668 21440
rect 86736 21384 86792 21440
rect 86860 21384 86916 21440
rect 86984 21384 87040 21440
rect 86612 21260 86668 21316
rect 86736 21260 86792 21316
rect 86860 21260 86916 21316
rect 86984 21260 87040 21316
rect 86612 21136 86668 21192
rect 86736 21136 86792 21192
rect 86860 21136 86916 21192
rect 86984 21136 87040 21192
rect 1130 20608 1186 20664
rect 1254 20608 1310 20664
rect 1378 20608 1434 20664
rect 1502 20608 1558 20664
rect 1130 20484 1186 20540
rect 1254 20484 1310 20540
rect 1378 20484 1434 20540
rect 1502 20484 1558 20540
rect 1130 20360 1186 20416
rect 1254 20360 1310 20416
rect 1378 20360 1434 20416
rect 1502 20360 1558 20416
rect 1130 20236 1186 20292
rect 1254 20236 1310 20292
rect 1378 20236 1434 20292
rect 1502 20236 1558 20292
rect 85812 20608 85868 20664
rect 85936 20608 85992 20664
rect 86060 20608 86116 20664
rect 86184 20608 86240 20664
rect 85812 20484 85868 20540
rect 85936 20484 85992 20540
rect 86060 20484 86116 20540
rect 86184 20484 86240 20540
rect 85812 20360 85868 20416
rect 85936 20360 85992 20416
rect 86060 20360 86116 20416
rect 86184 20360 86240 20416
rect 85812 20236 85868 20292
rect 85936 20236 85992 20292
rect 86060 20236 86116 20292
rect 86184 20236 86240 20292
rect 86612 19708 86668 19764
rect 86736 19708 86792 19764
rect 86860 19708 86916 19764
rect 86984 19708 87040 19764
rect 1930 19584 1986 19640
rect 2054 19584 2110 19640
rect 2178 19584 2234 19640
rect 2302 19584 2358 19640
rect 1930 19460 1986 19516
rect 2054 19460 2110 19516
rect 2178 19460 2234 19516
rect 2302 19460 2358 19516
rect 86612 19584 86668 19640
rect 86736 19584 86792 19640
rect 86860 19584 86916 19640
rect 86984 19584 87040 19640
rect 86612 19460 86668 19516
rect 86736 19460 86792 19516
rect 86860 19460 86916 19516
rect 86984 19460 87040 19516
rect 86612 19336 86668 19392
rect 86736 19336 86792 19392
rect 86860 19336 86916 19392
rect 86984 19336 87040 19392
rect 1130 18808 1186 18864
rect 1254 18808 1310 18864
rect 1378 18808 1434 18864
rect 1502 18808 1558 18864
rect 1130 18684 1186 18740
rect 1254 18684 1310 18740
rect 1378 18684 1434 18740
rect 1502 18684 1558 18740
rect 1130 18560 1186 18616
rect 1254 18560 1310 18616
rect 1378 18560 1434 18616
rect 1502 18560 1558 18616
rect 1130 18436 1186 18492
rect 1254 18436 1310 18492
rect 1378 18436 1434 18492
rect 1502 18436 1558 18492
rect 85812 18808 85868 18864
rect 85936 18808 85992 18864
rect 86060 18808 86116 18864
rect 86184 18808 86240 18864
rect 85812 18684 85868 18740
rect 85936 18684 85992 18740
rect 86060 18684 86116 18740
rect 86184 18684 86240 18740
rect 85812 18560 85868 18616
rect 85936 18560 85992 18616
rect 86060 18560 86116 18616
rect 86184 18560 86240 18616
rect 85812 18436 85868 18492
rect 85936 18436 85992 18492
rect 86060 18436 86116 18492
rect 86184 18436 86240 18492
rect 86612 17908 86668 17964
rect 86736 17908 86792 17964
rect 86860 17908 86916 17964
rect 86984 17908 87040 17964
rect 1930 17784 1986 17840
rect 2054 17784 2110 17840
rect 2178 17784 2234 17840
rect 2302 17784 2358 17840
rect 1930 17660 1986 17716
rect 2054 17660 2110 17716
rect 2178 17660 2234 17716
rect 2302 17660 2358 17716
rect 86612 17784 86668 17840
rect 86736 17784 86792 17840
rect 86860 17784 86916 17840
rect 86984 17784 87040 17840
rect 86612 17660 86668 17716
rect 86736 17660 86792 17716
rect 86860 17660 86916 17716
rect 86984 17660 87040 17716
rect 86612 17536 86668 17592
rect 86736 17536 86792 17592
rect 86860 17536 86916 17592
rect 86984 17536 87040 17592
rect 1130 17008 1186 17064
rect 1254 17008 1310 17064
rect 1378 17008 1434 17064
rect 1502 17008 1558 17064
rect 1130 16884 1186 16940
rect 1254 16884 1310 16940
rect 1378 16884 1434 16940
rect 1502 16884 1558 16940
rect 1130 16760 1186 16816
rect 1254 16760 1310 16816
rect 1378 16760 1434 16816
rect 1502 16760 1558 16816
rect 1130 16636 1186 16692
rect 1254 16636 1310 16692
rect 1378 16636 1434 16692
rect 1502 16636 1558 16692
rect 85812 17008 85868 17064
rect 85936 17008 85992 17064
rect 86060 17008 86116 17064
rect 86184 17008 86240 17064
rect 85812 16884 85868 16940
rect 85936 16884 85992 16940
rect 86060 16884 86116 16940
rect 86184 16884 86240 16940
rect 85812 16760 85868 16816
rect 85936 16760 85992 16816
rect 86060 16760 86116 16816
rect 86184 16760 86240 16816
rect 85812 16636 85868 16692
rect 85936 16636 85992 16692
rect 86060 16636 86116 16692
rect 86184 16636 86240 16692
rect 86612 16108 86668 16164
rect 86736 16108 86792 16164
rect 86860 16108 86916 16164
rect 86984 16108 87040 16164
rect 1930 15984 1986 16040
rect 2054 15984 2110 16040
rect 2178 15984 2234 16040
rect 2302 15984 2358 16040
rect 1930 15860 1986 15916
rect 2054 15860 2110 15916
rect 2178 15860 2234 15916
rect 2302 15860 2358 15916
rect 86612 15984 86668 16040
rect 86736 15984 86792 16040
rect 86860 15984 86916 16040
rect 86984 15984 87040 16040
rect 86612 15860 86668 15916
rect 86736 15860 86792 15916
rect 86860 15860 86916 15916
rect 86984 15860 87040 15916
rect 86612 15736 86668 15792
rect 86736 15736 86792 15792
rect 86860 15736 86916 15792
rect 86984 15736 87040 15792
rect 1130 15208 1186 15264
rect 1254 15208 1310 15264
rect 1378 15208 1434 15264
rect 1502 15208 1558 15264
rect 1130 15084 1186 15140
rect 1254 15084 1310 15140
rect 1378 15084 1434 15140
rect 1502 15084 1558 15140
rect 1130 14960 1186 15016
rect 1254 14960 1310 15016
rect 1378 14960 1434 15016
rect 1502 14960 1558 15016
rect 1130 14836 1186 14892
rect 1254 14836 1310 14892
rect 1378 14836 1434 14892
rect 1502 14836 1558 14892
rect 85812 15208 85868 15264
rect 85936 15208 85992 15264
rect 86060 15208 86116 15264
rect 86184 15208 86240 15264
rect 85812 15084 85868 15140
rect 85936 15084 85992 15140
rect 86060 15084 86116 15140
rect 86184 15084 86240 15140
rect 85812 14960 85868 15016
rect 85936 14960 85992 15016
rect 86060 14960 86116 15016
rect 86184 14960 86240 15016
rect 85812 14836 85868 14892
rect 85936 14836 85992 14892
rect 86060 14836 86116 14892
rect 86184 14836 86240 14892
rect 86612 14308 86668 14364
rect 86736 14308 86792 14364
rect 86860 14308 86916 14364
rect 86984 14308 87040 14364
rect 1930 14184 1986 14240
rect 2054 14184 2110 14240
rect 2178 14184 2234 14240
rect 2302 14184 2358 14240
rect 1930 14060 1986 14116
rect 2054 14060 2110 14116
rect 2178 14060 2234 14116
rect 2302 14060 2358 14116
rect 86612 14184 86668 14240
rect 86736 14184 86792 14240
rect 86860 14184 86916 14240
rect 86984 14184 87040 14240
rect 86612 14060 86668 14116
rect 86736 14060 86792 14116
rect 86860 14060 86916 14116
rect 86984 14060 87040 14116
rect 86612 13936 86668 13992
rect 86736 13936 86792 13992
rect 86860 13936 86916 13992
rect 86984 13936 87040 13992
rect 1130 13408 1186 13464
rect 1254 13408 1310 13464
rect 1378 13408 1434 13464
rect 1502 13408 1558 13464
rect 1130 13284 1186 13340
rect 1254 13284 1310 13340
rect 1378 13284 1434 13340
rect 1502 13284 1558 13340
rect 1130 13160 1186 13216
rect 1254 13160 1310 13216
rect 1378 13160 1434 13216
rect 1502 13160 1558 13216
rect 1130 13036 1186 13092
rect 1254 13036 1310 13092
rect 1378 13036 1434 13092
rect 1502 13036 1558 13092
rect 85812 13408 85868 13464
rect 85936 13408 85992 13464
rect 86060 13408 86116 13464
rect 86184 13408 86240 13464
rect 85812 13284 85868 13340
rect 85936 13284 85992 13340
rect 86060 13284 86116 13340
rect 86184 13284 86240 13340
rect 85812 13160 85868 13216
rect 85936 13160 85992 13216
rect 86060 13160 86116 13216
rect 86184 13160 86240 13216
rect 85812 13036 85868 13092
rect 85936 13036 85992 13092
rect 86060 13036 86116 13092
rect 86184 13036 86240 13092
rect 86612 12508 86668 12564
rect 86736 12508 86792 12564
rect 86860 12508 86916 12564
rect 86984 12508 87040 12564
rect 1930 12384 1986 12440
rect 2054 12384 2110 12440
rect 2178 12384 2234 12440
rect 2302 12384 2358 12440
rect 1930 12260 1986 12316
rect 2054 12260 2110 12316
rect 2178 12260 2234 12316
rect 2302 12260 2358 12316
rect 86612 12384 86668 12440
rect 86736 12384 86792 12440
rect 86860 12384 86916 12440
rect 86984 12384 87040 12440
rect 86612 12260 86668 12316
rect 86736 12260 86792 12316
rect 86860 12260 86916 12316
rect 86984 12260 87040 12316
rect 86612 12136 86668 12192
rect 86736 12136 86792 12192
rect 86860 12136 86916 12192
rect 86984 12136 87040 12192
rect 1130 11608 1186 11664
rect 1254 11608 1310 11664
rect 1378 11608 1434 11664
rect 1502 11608 1558 11664
rect 1130 11484 1186 11540
rect 1254 11484 1310 11540
rect 1378 11484 1434 11540
rect 1502 11484 1558 11540
rect 1130 11360 1186 11416
rect 1254 11360 1310 11416
rect 1378 11360 1434 11416
rect 1502 11360 1558 11416
rect 1130 11236 1186 11292
rect 1254 11236 1310 11292
rect 1378 11236 1434 11292
rect 1502 11236 1558 11292
rect 85812 11608 85868 11664
rect 85936 11608 85992 11664
rect 86060 11608 86116 11664
rect 86184 11608 86240 11664
rect 85812 11484 85868 11540
rect 85936 11484 85992 11540
rect 86060 11484 86116 11540
rect 86184 11484 86240 11540
rect 85812 11360 85868 11416
rect 85936 11360 85992 11416
rect 86060 11360 86116 11416
rect 86184 11360 86240 11416
rect 85812 11236 85868 11292
rect 85936 11236 85992 11292
rect 86060 11236 86116 11292
rect 86184 11236 86240 11292
rect 86612 10708 86668 10764
rect 86736 10708 86792 10764
rect 86860 10708 86916 10764
rect 86984 10708 87040 10764
rect 1930 10584 1986 10640
rect 2054 10584 2110 10640
rect 2178 10584 2234 10640
rect 2302 10584 2358 10640
rect 1930 10460 1986 10516
rect 2054 10460 2110 10516
rect 2178 10460 2234 10516
rect 2302 10460 2358 10516
rect 86612 10584 86668 10640
rect 86736 10584 86792 10640
rect 86860 10584 86916 10640
rect 86984 10584 87040 10640
rect 86612 10460 86668 10516
rect 86736 10460 86792 10516
rect 86860 10460 86916 10516
rect 86984 10460 87040 10516
rect 86612 10336 86668 10392
rect 86736 10336 86792 10392
rect 86860 10336 86916 10392
rect 86984 10336 87040 10392
rect 1130 9808 1186 9864
rect 1254 9808 1310 9864
rect 1378 9808 1434 9864
rect 1502 9808 1558 9864
rect 1130 9684 1186 9740
rect 1254 9684 1310 9740
rect 1378 9684 1434 9740
rect 1502 9684 1558 9740
rect 1130 9560 1186 9616
rect 1254 9560 1310 9616
rect 1378 9560 1434 9616
rect 1502 9560 1558 9616
rect 1130 9436 1186 9492
rect 1254 9436 1310 9492
rect 1378 9436 1434 9492
rect 1502 9436 1558 9492
rect 85812 9808 85868 9864
rect 85936 9808 85992 9864
rect 86060 9808 86116 9864
rect 86184 9808 86240 9864
rect 85812 9684 85868 9740
rect 85936 9684 85992 9740
rect 86060 9684 86116 9740
rect 86184 9684 86240 9740
rect 85812 9560 85868 9616
rect 85936 9560 85992 9616
rect 86060 9560 86116 9616
rect 86184 9560 86240 9616
rect 85812 9436 85868 9492
rect 85936 9436 85992 9492
rect 86060 9436 86116 9492
rect 86184 9436 86240 9492
rect 86612 8908 86668 8964
rect 86736 8908 86792 8964
rect 86860 8908 86916 8964
rect 86984 8908 87040 8964
rect 1930 8784 1986 8840
rect 2054 8784 2110 8840
rect 2178 8784 2234 8840
rect 2302 8784 2358 8840
rect 1930 8660 1986 8716
rect 2054 8660 2110 8716
rect 2178 8660 2234 8716
rect 2302 8660 2358 8716
rect 86612 8784 86668 8840
rect 86736 8784 86792 8840
rect 86860 8784 86916 8840
rect 86984 8784 87040 8840
rect 86612 8660 86668 8716
rect 86736 8660 86792 8716
rect 86860 8660 86916 8716
rect 86984 8660 87040 8716
rect 86612 8536 86668 8592
rect 86736 8536 86792 8592
rect 86860 8536 86916 8592
rect 86984 8536 87040 8592
rect 1130 8008 1186 8064
rect 1254 8008 1310 8064
rect 1378 8008 1434 8064
rect 1502 8008 1558 8064
rect 1130 7884 1186 7940
rect 1254 7884 1310 7940
rect 1378 7884 1434 7940
rect 1502 7884 1558 7940
rect 1130 7760 1186 7816
rect 1254 7760 1310 7816
rect 1378 7760 1434 7816
rect 1502 7760 1558 7816
rect 1130 7636 1186 7692
rect 1254 7636 1310 7692
rect 1378 7636 1434 7692
rect 1502 7636 1558 7692
rect 85812 8008 85868 8064
rect 85936 8008 85992 8064
rect 86060 8008 86116 8064
rect 86184 8008 86240 8064
rect 85812 7884 85868 7940
rect 85936 7884 85992 7940
rect 86060 7884 86116 7940
rect 86184 7884 86240 7940
rect 85812 7760 85868 7816
rect 85936 7760 85992 7816
rect 86060 7760 86116 7816
rect 86184 7760 86240 7816
rect 85812 7636 85868 7692
rect 85936 7636 85992 7692
rect 86060 7636 86116 7692
rect 86184 7636 86240 7692
rect 86612 7108 86668 7164
rect 86736 7108 86792 7164
rect 86860 7108 86916 7164
rect 86984 7108 87040 7164
rect 1930 6984 1986 7040
rect 2054 6984 2110 7040
rect 2178 6984 2234 7040
rect 2302 6984 2358 7040
rect 1930 6860 1986 6916
rect 2054 6860 2110 6916
rect 2178 6860 2234 6916
rect 2302 6860 2358 6916
rect 86612 6984 86668 7040
rect 86736 6984 86792 7040
rect 86860 6984 86916 7040
rect 86984 6984 87040 7040
rect 86612 6860 86668 6916
rect 86736 6860 86792 6916
rect 86860 6860 86916 6916
rect 86984 6860 87040 6916
rect 86612 6736 86668 6792
rect 86736 6736 86792 6792
rect 86860 6736 86916 6792
rect 86984 6736 87040 6792
rect 1130 6208 1186 6264
rect 1254 6208 1310 6264
rect 1378 6208 1434 6264
rect 1502 6208 1558 6264
rect 1130 6084 1186 6140
rect 1254 6084 1310 6140
rect 1378 6084 1434 6140
rect 1502 6084 1558 6140
rect 1130 5960 1186 6016
rect 1254 5960 1310 6016
rect 1378 5960 1434 6016
rect 1502 5960 1558 6016
rect 1130 5836 1186 5892
rect 1254 5836 1310 5892
rect 1378 5836 1434 5892
rect 1502 5836 1558 5892
rect 85812 6208 85868 6264
rect 85936 6208 85992 6264
rect 86060 6208 86116 6264
rect 86184 6208 86240 6264
rect 85812 6084 85868 6140
rect 85936 6084 85992 6140
rect 86060 6084 86116 6140
rect 86184 6084 86240 6140
rect 85812 5960 85868 6016
rect 85936 5960 85992 6016
rect 86060 5960 86116 6016
rect 86184 5960 86240 6016
rect 85812 5836 85868 5892
rect 85936 5836 85992 5892
rect 86060 5836 86116 5892
rect 86184 5836 86240 5892
rect 86612 5308 86668 5364
rect 86736 5308 86792 5364
rect 86860 5308 86916 5364
rect 86984 5308 87040 5364
rect 1930 5184 1986 5240
rect 2054 5184 2110 5240
rect 2178 5184 2234 5240
rect 2302 5184 2358 5240
rect 1930 5060 1986 5116
rect 2054 5060 2110 5116
rect 2178 5060 2234 5116
rect 2302 5060 2358 5116
rect 86612 5184 86668 5240
rect 86736 5184 86792 5240
rect 86860 5184 86916 5240
rect 86984 5184 87040 5240
rect 86612 5060 86668 5116
rect 86736 5060 86792 5116
rect 86860 5060 86916 5116
rect 86984 5060 87040 5116
rect 86612 4936 86668 4992
rect 86736 4936 86792 4992
rect 86860 4936 86916 4992
rect 86984 4936 87040 4992
rect 1130 4408 1186 4464
rect 1254 4408 1310 4464
rect 1378 4408 1434 4464
rect 1502 4408 1558 4464
rect 1130 4284 1186 4340
rect 1254 4284 1310 4340
rect 1378 4284 1434 4340
rect 1502 4284 1558 4340
rect 1130 4160 1186 4216
rect 1254 4160 1310 4216
rect 1378 4160 1434 4216
rect 1502 4160 1558 4216
rect 1130 4036 1186 4092
rect 1254 4036 1310 4092
rect 1378 4036 1434 4092
rect 1502 4036 1558 4092
rect 85812 4408 85868 4464
rect 85936 4408 85992 4464
rect 86060 4408 86116 4464
rect 86184 4408 86240 4464
rect 85812 4284 85868 4340
rect 85936 4284 85992 4340
rect 86060 4284 86116 4340
rect 86184 4284 86240 4340
rect 85812 4160 85868 4216
rect 85936 4160 85992 4216
rect 86060 4160 86116 4216
rect 86184 4160 86240 4216
rect 85812 4036 85868 4092
rect 85936 4036 85992 4092
rect 86060 4036 86116 4092
rect 86184 4036 86240 4092
rect 86612 3576 86668 3632
rect 86736 3576 86792 3632
rect 86860 3576 86916 3632
rect 86984 3576 87040 3632
rect 1930 3384 1986 3440
rect 2054 3384 2110 3440
rect 2178 3384 2234 3440
rect 2302 3384 2358 3440
rect 1930 3260 1986 3316
rect 2054 3260 2110 3316
rect 2178 3260 2234 3316
rect 2302 3260 2358 3316
rect 86612 3452 86668 3508
rect 86736 3452 86792 3508
rect 86860 3452 86916 3508
rect 86984 3452 87040 3508
rect 86612 3328 86668 3384
rect 86736 3328 86792 3384
rect 86860 3328 86916 3384
rect 86984 3328 87040 3384
rect 86612 3204 86668 3260
rect 86736 3204 86792 3260
rect 86860 3204 86916 3260
rect 86984 3204 87040 3260
<< metal4 >>
rect 1044 57089 1644 66640
rect 1044 57033 1068 57089
rect 1124 57033 1192 57089
rect 1248 57033 1316 57089
rect 1372 57033 1440 57089
rect 1496 57033 1564 57089
rect 1620 57033 1644 57089
rect 1044 56965 1644 57033
rect 1044 56909 1068 56965
rect 1124 56909 1192 56965
rect 1248 56909 1316 56965
rect 1372 56909 1440 56965
rect 1496 56909 1564 56965
rect 1620 56909 1644 56965
rect 1044 56841 1644 56909
rect 1044 56785 1068 56841
rect 1124 56785 1192 56841
rect 1248 56785 1316 56841
rect 1372 56785 1440 56841
rect 1496 56785 1564 56841
rect 1620 56785 1644 56841
rect 1044 56717 1644 56785
rect 1044 56661 1068 56717
rect 1124 56661 1192 56717
rect 1248 56661 1316 56717
rect 1372 56661 1440 56717
rect 1496 56661 1564 56717
rect 1620 56661 1644 56717
rect 1044 56593 1644 56661
rect 1044 56537 1068 56593
rect 1124 56537 1192 56593
rect 1248 56537 1316 56593
rect 1372 56537 1440 56593
rect 1496 56537 1564 56593
rect 1620 56537 1644 56593
rect 1044 56469 1644 56537
rect 1044 56413 1068 56469
rect 1124 56413 1192 56469
rect 1248 56413 1316 56469
rect 1372 56413 1440 56469
rect 1496 56413 1564 56469
rect 1620 56413 1644 56469
rect 1044 56345 1644 56413
rect 1044 56289 1068 56345
rect 1124 56289 1192 56345
rect 1248 56289 1316 56345
rect 1372 56289 1440 56345
rect 1496 56289 1564 56345
rect 1620 56289 1644 56345
rect 1044 56221 1644 56289
rect 1044 56165 1068 56221
rect 1124 56165 1192 56221
rect 1248 56165 1316 56221
rect 1372 56165 1440 56221
rect 1496 56165 1564 56221
rect 1620 56165 1644 56221
rect 1044 56097 1644 56165
rect 1044 56041 1068 56097
rect 1124 56041 1192 56097
rect 1248 56041 1316 56097
rect 1372 56041 1440 56097
rect 1496 56041 1564 56097
rect 1620 56041 1644 56097
rect 1044 55973 1644 56041
rect 1044 55917 1068 55973
rect 1124 55917 1192 55973
rect 1248 55917 1316 55973
rect 1372 55917 1440 55973
rect 1496 55917 1564 55973
rect 1620 55917 1644 55973
rect 1044 55849 1644 55917
rect 1044 55793 1068 55849
rect 1124 55793 1192 55849
rect 1248 55793 1316 55849
rect 1372 55793 1440 55849
rect 1496 55793 1564 55849
rect 1620 55793 1644 55849
rect 1044 55725 1644 55793
rect 1044 55669 1068 55725
rect 1124 55669 1192 55725
rect 1248 55669 1316 55725
rect 1372 55669 1440 55725
rect 1496 55669 1564 55725
rect 1620 55669 1644 55725
rect 1044 55601 1644 55669
rect 1044 55545 1068 55601
rect 1124 55545 1192 55601
rect 1248 55545 1316 55601
rect 1372 55545 1440 55601
rect 1496 55545 1564 55601
rect 1620 55545 1644 55601
rect 1044 55477 1644 55545
rect 1044 55421 1068 55477
rect 1124 55421 1192 55477
rect 1248 55421 1316 55477
rect 1372 55421 1440 55477
rect 1496 55421 1564 55477
rect 1620 55421 1644 55477
rect 1044 55353 1644 55421
rect 1044 55297 1068 55353
rect 1124 55297 1192 55353
rect 1248 55297 1316 55353
rect 1372 55297 1440 55353
rect 1496 55297 1564 55353
rect 1620 55297 1644 55353
rect 1044 55229 1644 55297
rect 1044 55173 1068 55229
rect 1124 55173 1192 55229
rect 1248 55173 1316 55229
rect 1372 55173 1440 55229
rect 1496 55173 1564 55229
rect 1620 55173 1644 55229
rect 1044 55105 1644 55173
rect 1044 55049 1068 55105
rect 1124 55049 1192 55105
rect 1248 55049 1316 55105
rect 1372 55049 1440 55105
rect 1496 55049 1564 55105
rect 1620 55049 1644 55105
rect 1044 46200 1644 55049
rect 1044 46144 1068 46200
rect 1124 46144 1192 46200
rect 1248 46144 1316 46200
rect 1372 46144 1440 46200
rect 1496 46144 1564 46200
rect 1620 46144 1644 46200
rect 1044 46076 1644 46144
rect 1044 46020 1068 46076
rect 1124 46020 1192 46076
rect 1248 46020 1316 46076
rect 1372 46020 1440 46076
rect 1496 46020 1564 46076
rect 1620 46020 1644 46076
rect 1044 45952 1644 46020
rect 1044 45896 1068 45952
rect 1124 45896 1192 45952
rect 1248 45896 1316 45952
rect 1372 45896 1440 45952
rect 1496 45896 1564 45952
rect 1620 45896 1644 45952
rect 1044 45828 1644 45896
rect 1044 45772 1068 45828
rect 1124 45772 1192 45828
rect 1248 45772 1316 45828
rect 1372 45772 1440 45828
rect 1496 45772 1564 45828
rect 1620 45772 1644 45828
rect 1044 45704 1644 45772
rect 1044 45648 1068 45704
rect 1124 45648 1192 45704
rect 1248 45648 1316 45704
rect 1372 45648 1440 45704
rect 1496 45648 1564 45704
rect 1620 45648 1644 45704
rect 1044 45580 1644 45648
rect 1044 45524 1068 45580
rect 1124 45524 1192 45580
rect 1248 45524 1316 45580
rect 1372 45524 1440 45580
rect 1496 45524 1564 45580
rect 1620 45524 1644 45580
rect 1044 45456 1644 45524
rect 1044 45400 1068 45456
rect 1124 45400 1192 45456
rect 1248 45400 1316 45456
rect 1372 45400 1440 45456
rect 1496 45400 1564 45456
rect 1620 45400 1644 45456
rect 1044 45332 1644 45400
rect 1044 45276 1068 45332
rect 1124 45276 1192 45332
rect 1248 45276 1316 45332
rect 1372 45276 1440 45332
rect 1496 45276 1564 45332
rect 1620 45276 1644 45332
rect 1044 33264 1644 45276
rect 1044 33208 1130 33264
rect 1186 33208 1254 33264
rect 1310 33208 1378 33264
rect 1434 33208 1502 33264
rect 1558 33208 1644 33264
rect 1044 33140 1644 33208
rect 1044 33084 1130 33140
rect 1186 33084 1254 33140
rect 1310 33084 1378 33140
rect 1434 33084 1502 33140
rect 1558 33084 1644 33140
rect 1044 33016 1644 33084
rect 1044 32960 1130 33016
rect 1186 32960 1254 33016
rect 1310 32960 1378 33016
rect 1434 32960 1502 33016
rect 1558 32960 1644 33016
rect 1044 32892 1644 32960
rect 1044 32836 1130 32892
rect 1186 32836 1254 32892
rect 1310 32836 1378 32892
rect 1434 32836 1502 32892
rect 1558 32836 1644 32892
rect 1044 31464 1644 32836
rect 1044 31408 1130 31464
rect 1186 31408 1254 31464
rect 1310 31408 1378 31464
rect 1434 31408 1502 31464
rect 1558 31408 1644 31464
rect 1044 31340 1644 31408
rect 1044 31284 1130 31340
rect 1186 31284 1254 31340
rect 1310 31284 1378 31340
rect 1434 31284 1502 31340
rect 1558 31284 1644 31340
rect 1044 31216 1644 31284
rect 1044 31160 1130 31216
rect 1186 31160 1254 31216
rect 1310 31160 1378 31216
rect 1434 31160 1502 31216
rect 1558 31160 1644 31216
rect 1044 31092 1644 31160
rect 1044 31036 1130 31092
rect 1186 31036 1254 31092
rect 1310 31036 1378 31092
rect 1434 31036 1502 31092
rect 1558 31036 1644 31092
rect 1044 29664 1644 31036
rect 1044 29608 1130 29664
rect 1186 29608 1254 29664
rect 1310 29608 1378 29664
rect 1434 29608 1502 29664
rect 1558 29608 1644 29664
rect 1044 29540 1644 29608
rect 1044 29484 1130 29540
rect 1186 29484 1254 29540
rect 1310 29484 1378 29540
rect 1434 29484 1502 29540
rect 1558 29484 1644 29540
rect 1044 29416 1644 29484
rect 1044 29360 1130 29416
rect 1186 29360 1254 29416
rect 1310 29360 1378 29416
rect 1434 29360 1502 29416
rect 1558 29360 1644 29416
rect 1044 29292 1644 29360
rect 1044 29236 1130 29292
rect 1186 29236 1254 29292
rect 1310 29236 1378 29292
rect 1434 29236 1502 29292
rect 1558 29236 1644 29292
rect 1044 27864 1644 29236
rect 1044 27808 1130 27864
rect 1186 27808 1254 27864
rect 1310 27808 1378 27864
rect 1434 27808 1502 27864
rect 1558 27808 1644 27864
rect 1044 27740 1644 27808
rect 1044 27684 1130 27740
rect 1186 27684 1254 27740
rect 1310 27684 1378 27740
rect 1434 27684 1502 27740
rect 1558 27684 1644 27740
rect 1044 27616 1644 27684
rect 1044 27560 1130 27616
rect 1186 27560 1254 27616
rect 1310 27560 1378 27616
rect 1434 27560 1502 27616
rect 1558 27560 1644 27616
rect 1044 27492 1644 27560
rect 1044 27436 1130 27492
rect 1186 27436 1254 27492
rect 1310 27436 1378 27492
rect 1434 27436 1502 27492
rect 1558 27436 1644 27492
rect 1044 26064 1644 27436
rect 1044 26008 1130 26064
rect 1186 26008 1254 26064
rect 1310 26008 1378 26064
rect 1434 26008 1502 26064
rect 1558 26008 1644 26064
rect 1044 25940 1644 26008
rect 1044 25884 1130 25940
rect 1186 25884 1254 25940
rect 1310 25884 1378 25940
rect 1434 25884 1502 25940
rect 1558 25884 1644 25940
rect 1044 25816 1644 25884
rect 1044 25760 1130 25816
rect 1186 25760 1254 25816
rect 1310 25760 1378 25816
rect 1434 25760 1502 25816
rect 1558 25760 1644 25816
rect 1044 25692 1644 25760
rect 1044 25636 1130 25692
rect 1186 25636 1254 25692
rect 1310 25636 1378 25692
rect 1434 25636 1502 25692
rect 1558 25636 1644 25692
rect 1044 24264 1644 25636
rect 1044 24208 1130 24264
rect 1186 24208 1254 24264
rect 1310 24208 1378 24264
rect 1434 24208 1502 24264
rect 1558 24208 1644 24264
rect 1044 24140 1644 24208
rect 1044 24084 1130 24140
rect 1186 24084 1254 24140
rect 1310 24084 1378 24140
rect 1434 24084 1502 24140
rect 1558 24084 1644 24140
rect 1044 24016 1644 24084
rect 1044 23960 1130 24016
rect 1186 23960 1254 24016
rect 1310 23960 1378 24016
rect 1434 23960 1502 24016
rect 1558 23960 1644 24016
rect 1044 23892 1644 23960
rect 1044 23836 1130 23892
rect 1186 23836 1254 23892
rect 1310 23836 1378 23892
rect 1434 23836 1502 23892
rect 1558 23836 1644 23892
rect 1044 22464 1644 23836
rect 1044 22408 1130 22464
rect 1186 22408 1254 22464
rect 1310 22408 1378 22464
rect 1434 22408 1502 22464
rect 1558 22408 1644 22464
rect 1044 22340 1644 22408
rect 1044 22284 1130 22340
rect 1186 22284 1254 22340
rect 1310 22284 1378 22340
rect 1434 22284 1502 22340
rect 1558 22284 1644 22340
rect 1044 22216 1644 22284
rect 1044 22160 1130 22216
rect 1186 22160 1254 22216
rect 1310 22160 1378 22216
rect 1434 22160 1502 22216
rect 1558 22160 1644 22216
rect 1044 22092 1644 22160
rect 1044 22036 1130 22092
rect 1186 22036 1254 22092
rect 1310 22036 1378 22092
rect 1434 22036 1502 22092
rect 1558 22036 1644 22092
rect 1044 20664 1644 22036
rect 1044 20608 1130 20664
rect 1186 20608 1254 20664
rect 1310 20608 1378 20664
rect 1434 20608 1502 20664
rect 1558 20608 1644 20664
rect 1044 20540 1644 20608
rect 1044 20484 1130 20540
rect 1186 20484 1254 20540
rect 1310 20484 1378 20540
rect 1434 20484 1502 20540
rect 1558 20484 1644 20540
rect 1044 20416 1644 20484
rect 1044 20360 1130 20416
rect 1186 20360 1254 20416
rect 1310 20360 1378 20416
rect 1434 20360 1502 20416
rect 1558 20360 1644 20416
rect 1044 20292 1644 20360
rect 1044 20236 1130 20292
rect 1186 20236 1254 20292
rect 1310 20236 1378 20292
rect 1434 20236 1502 20292
rect 1558 20236 1644 20292
rect 1044 18864 1644 20236
rect 1044 18808 1130 18864
rect 1186 18808 1254 18864
rect 1310 18808 1378 18864
rect 1434 18808 1502 18864
rect 1558 18808 1644 18864
rect 1044 18740 1644 18808
rect 1044 18684 1130 18740
rect 1186 18684 1254 18740
rect 1310 18684 1378 18740
rect 1434 18684 1502 18740
rect 1558 18684 1644 18740
rect 1044 18616 1644 18684
rect 1044 18560 1130 18616
rect 1186 18560 1254 18616
rect 1310 18560 1378 18616
rect 1434 18560 1502 18616
rect 1558 18560 1644 18616
rect 1044 18492 1644 18560
rect 1044 18436 1130 18492
rect 1186 18436 1254 18492
rect 1310 18436 1378 18492
rect 1434 18436 1502 18492
rect 1558 18436 1644 18492
rect 1044 17064 1644 18436
rect 1044 17008 1130 17064
rect 1186 17008 1254 17064
rect 1310 17008 1378 17064
rect 1434 17008 1502 17064
rect 1558 17008 1644 17064
rect 1044 16940 1644 17008
rect 1044 16884 1130 16940
rect 1186 16884 1254 16940
rect 1310 16884 1378 16940
rect 1434 16884 1502 16940
rect 1558 16884 1644 16940
rect 1044 16816 1644 16884
rect 1044 16760 1130 16816
rect 1186 16760 1254 16816
rect 1310 16760 1378 16816
rect 1434 16760 1502 16816
rect 1558 16760 1644 16816
rect 1044 16692 1644 16760
rect 1044 16636 1130 16692
rect 1186 16636 1254 16692
rect 1310 16636 1378 16692
rect 1434 16636 1502 16692
rect 1558 16636 1644 16692
rect 1044 15264 1644 16636
rect 1044 15208 1130 15264
rect 1186 15208 1254 15264
rect 1310 15208 1378 15264
rect 1434 15208 1502 15264
rect 1558 15208 1644 15264
rect 1044 15140 1644 15208
rect 1044 15084 1130 15140
rect 1186 15084 1254 15140
rect 1310 15084 1378 15140
rect 1434 15084 1502 15140
rect 1558 15084 1644 15140
rect 1044 15016 1644 15084
rect 1044 14960 1130 15016
rect 1186 14960 1254 15016
rect 1310 14960 1378 15016
rect 1434 14960 1502 15016
rect 1558 14960 1644 15016
rect 1044 14892 1644 14960
rect 1044 14836 1130 14892
rect 1186 14836 1254 14892
rect 1310 14836 1378 14892
rect 1434 14836 1502 14892
rect 1558 14836 1644 14892
rect 1044 13464 1644 14836
rect 1044 13408 1130 13464
rect 1186 13408 1254 13464
rect 1310 13408 1378 13464
rect 1434 13408 1502 13464
rect 1558 13408 1644 13464
rect 1044 13340 1644 13408
rect 1044 13284 1130 13340
rect 1186 13284 1254 13340
rect 1310 13284 1378 13340
rect 1434 13284 1502 13340
rect 1558 13284 1644 13340
rect 1044 13216 1644 13284
rect 1044 13160 1130 13216
rect 1186 13160 1254 13216
rect 1310 13160 1378 13216
rect 1434 13160 1502 13216
rect 1558 13160 1644 13216
rect 1044 13092 1644 13160
rect 1044 13036 1130 13092
rect 1186 13036 1254 13092
rect 1310 13036 1378 13092
rect 1434 13036 1502 13092
rect 1558 13036 1644 13092
rect 1044 11664 1644 13036
rect 1044 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1644 11664
rect 1044 11540 1644 11608
rect 1044 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1644 11540
rect 1044 11416 1644 11484
rect 1044 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1644 11416
rect 1044 11292 1644 11360
rect 1044 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1644 11292
rect 1044 9864 1644 11236
rect 1044 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1644 9864
rect 1044 9740 1644 9808
rect 1044 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1644 9740
rect 1044 9616 1644 9684
rect 1044 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1644 9616
rect 1044 9492 1644 9560
rect 1044 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1644 9492
rect 1044 8064 1644 9436
rect 1044 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1644 8064
rect 1044 7940 1644 8008
rect 1044 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1644 7940
rect 1044 7816 1644 7884
rect 1044 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1644 7816
rect 1044 7692 1644 7760
rect 1044 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1644 7692
rect 1044 6264 1644 7636
rect 1044 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1644 6264
rect 1044 6140 1644 6208
rect 1044 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1644 6140
rect 1044 6016 1644 6084
rect 1044 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1644 6016
rect 1044 5892 1644 5960
rect 1044 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1644 5892
rect 1044 4464 1644 5836
rect 1044 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1644 4464
rect 1044 4340 1644 4408
rect 1044 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1644 4340
rect 1044 4216 1644 4284
rect 1044 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1644 4216
rect 1044 4092 1644 4160
rect 1044 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1644 4092
rect 1044 3136 1644 4036
rect 1844 66571 2444 66640
rect 1844 66515 1930 66571
rect 1986 66515 2054 66571
rect 2110 66515 2178 66571
rect 2234 66515 2302 66571
rect 2358 66515 2444 66571
rect 1844 66447 2444 66515
rect 1844 66391 1930 66447
rect 1986 66391 2054 66447
rect 2110 66391 2178 66447
rect 2234 66391 2302 66447
rect 2358 66391 2444 66447
rect 1844 65732 2444 66391
rect 1844 65676 1930 65732
rect 1986 65676 2054 65732
rect 2110 65676 2178 65732
rect 2234 65676 2302 65732
rect 2358 65676 2444 65732
rect 1844 65608 2444 65676
rect 1844 65552 1930 65608
rect 1986 65552 2054 65608
rect 2110 65552 2178 65608
rect 2234 65552 2302 65608
rect 2358 65552 2444 65608
rect 1844 65484 2444 65552
rect 1844 65428 1930 65484
rect 1986 65428 2054 65484
rect 2110 65428 2178 65484
rect 2234 65428 2302 65484
rect 2358 65428 2444 65484
rect 1844 63346 2444 65428
rect 1844 63290 1930 63346
rect 1986 63290 2054 63346
rect 2110 63290 2178 63346
rect 2234 63290 2302 63346
rect 2358 63290 2444 63346
rect 1844 63222 2444 63290
rect 1844 63166 1930 63222
rect 1986 63166 2054 63222
rect 2110 63166 2178 63222
rect 2234 63166 2302 63222
rect 2358 63166 2444 63222
rect 1844 63098 2444 63166
rect 1844 63042 1930 63098
rect 1986 63042 2054 63098
rect 2110 63042 2178 63098
rect 2234 63042 2302 63098
rect 2358 63042 2444 63098
rect 1844 62101 2444 63042
rect 1844 62045 1930 62101
rect 1986 62045 2054 62101
rect 2110 62045 2178 62101
rect 2234 62045 2302 62101
rect 2358 62045 2444 62101
rect 1844 61977 2444 62045
rect 1844 61921 1930 61977
rect 1986 61921 2054 61977
rect 2110 61921 2178 61977
rect 2234 61921 2302 61977
rect 2358 61921 2444 61977
rect 1844 61853 2444 61921
rect 1844 61797 1930 61853
rect 1986 61797 2054 61853
rect 2110 61797 2178 61853
rect 2234 61797 2302 61853
rect 2358 61797 2444 61853
rect 1844 61729 2444 61797
rect 1844 61673 1930 61729
rect 1986 61673 2054 61729
rect 2110 61673 2178 61729
rect 2234 61673 2302 61729
rect 2358 61673 2444 61729
rect 1844 54787 2444 61673
rect 1844 54731 1868 54787
rect 1924 54731 1992 54787
rect 2048 54731 2116 54787
rect 2172 54731 2240 54787
rect 2296 54731 2364 54787
rect 2420 54731 2444 54787
rect 1844 54663 2444 54731
rect 1844 54607 1868 54663
rect 1924 54607 1992 54663
rect 2048 54607 2116 54663
rect 2172 54607 2240 54663
rect 2296 54607 2364 54663
rect 2420 54607 2444 54663
rect 1844 54539 2444 54607
rect 1844 54483 1868 54539
rect 1924 54483 1992 54539
rect 2048 54483 2116 54539
rect 2172 54483 2240 54539
rect 2296 54483 2364 54539
rect 2420 54483 2444 54539
rect 1844 54415 2444 54483
rect 1844 54359 1868 54415
rect 1924 54359 1992 54415
rect 2048 54359 2116 54415
rect 2172 54359 2240 54415
rect 2296 54359 2364 54415
rect 2420 54359 2444 54415
rect 1844 54291 2444 54359
rect 1844 54235 1868 54291
rect 1924 54235 1992 54291
rect 2048 54235 2116 54291
rect 2172 54235 2240 54291
rect 2296 54235 2364 54291
rect 2420 54235 2444 54291
rect 1844 54167 2444 54235
rect 1844 54111 1868 54167
rect 1924 54111 1992 54167
rect 2048 54111 2116 54167
rect 2172 54111 2240 54167
rect 2296 54111 2364 54167
rect 2420 54111 2444 54167
rect 1844 54043 2444 54111
rect 1844 53987 1868 54043
rect 1924 53987 1992 54043
rect 2048 53987 2116 54043
rect 2172 53987 2240 54043
rect 2296 53987 2364 54043
rect 2420 53987 2444 54043
rect 1844 53919 2444 53987
rect 1844 53863 1868 53919
rect 1924 53863 1992 53919
rect 2048 53863 2116 53919
rect 2172 53863 2240 53919
rect 2296 53863 2364 53919
rect 2420 53863 2444 53919
rect 1844 53795 2444 53863
rect 1844 53739 1868 53795
rect 1924 53739 1992 53795
rect 2048 53739 2116 53795
rect 2172 53739 2240 53795
rect 2296 53739 2364 53795
rect 2420 53739 2444 53795
rect 1844 53671 2444 53739
rect 1844 53615 1868 53671
rect 1924 53615 1992 53671
rect 2048 53615 2116 53671
rect 2172 53615 2240 53671
rect 2296 53615 2364 53671
rect 2420 53615 2444 53671
rect 1844 53547 2444 53615
rect 1844 53491 1868 53547
rect 1924 53491 1992 53547
rect 2048 53491 2116 53547
rect 2172 53491 2240 53547
rect 2296 53491 2364 53547
rect 2420 53491 2444 53547
rect 1844 53423 2444 53491
rect 1844 53367 1868 53423
rect 1924 53367 1992 53423
rect 2048 53367 2116 53423
rect 2172 53367 2240 53423
rect 2296 53367 2364 53423
rect 2420 53367 2444 53423
rect 1844 53299 2444 53367
rect 1844 53243 1868 53299
rect 1924 53243 1992 53299
rect 2048 53243 2116 53299
rect 2172 53243 2240 53299
rect 2296 53243 2364 53299
rect 2420 53243 2444 53299
rect 1844 53175 2444 53243
rect 1844 53119 1868 53175
rect 1924 53119 1992 53175
rect 2048 53119 2116 53175
rect 2172 53119 2240 53175
rect 2296 53119 2364 53175
rect 2420 53119 2444 53175
rect 1844 53051 2444 53119
rect 1844 52995 1868 53051
rect 1924 52995 1992 53051
rect 2048 52995 2116 53051
rect 2172 52995 2240 53051
rect 2296 52995 2364 53051
rect 2420 52995 2444 53051
rect 1844 52927 2444 52995
rect 1844 52871 1868 52927
rect 1924 52871 1992 52927
rect 2048 52871 2116 52927
rect 2172 52871 2240 52927
rect 2296 52871 2364 52927
rect 2420 52871 2444 52927
rect 1844 52803 2444 52871
rect 1844 52747 1868 52803
rect 1924 52747 1992 52803
rect 2048 52747 2116 52803
rect 2172 52747 2240 52803
rect 2296 52747 2364 52803
rect 2420 52747 2444 52803
rect 1844 52679 2444 52747
rect 1844 52623 1868 52679
rect 1924 52623 1992 52679
rect 2048 52623 2116 52679
rect 2172 52623 2240 52679
rect 2296 52623 2364 52679
rect 2420 52623 2444 52679
rect 1844 52555 2444 52623
rect 1844 52499 1868 52555
rect 1924 52499 1992 52555
rect 2048 52499 2116 52555
rect 2172 52499 2240 52555
rect 2296 52499 2364 52555
rect 2420 52499 2444 52555
rect 1844 52431 2444 52499
rect 1844 52375 1868 52431
rect 1924 52375 1992 52431
rect 2048 52375 2116 52431
rect 2172 52375 2240 52431
rect 2296 52375 2364 52431
rect 2420 52375 2444 52431
rect 1844 52307 2444 52375
rect 1844 52251 1868 52307
rect 1924 52251 1992 52307
rect 2048 52251 2116 52307
rect 2172 52251 2240 52307
rect 2296 52251 2364 52307
rect 2420 52251 2444 52307
rect 1844 52183 2444 52251
rect 1844 52127 1868 52183
rect 1924 52127 1992 52183
rect 2048 52127 2116 52183
rect 2172 52127 2240 52183
rect 2296 52127 2364 52183
rect 2420 52127 2444 52183
rect 1844 52059 2444 52127
rect 1844 52003 1868 52059
rect 1924 52003 1992 52059
rect 2048 52003 2116 52059
rect 2172 52003 2240 52059
rect 2296 52003 2364 52059
rect 2420 52003 2444 52059
rect 1844 51935 2444 52003
rect 1844 51879 1868 51935
rect 1924 51879 1992 51935
rect 2048 51879 2116 51935
rect 2172 51879 2240 51935
rect 2296 51879 2364 51935
rect 2420 51879 2444 51935
rect 1844 51811 2444 51879
rect 1844 51755 1868 51811
rect 1924 51755 1992 51811
rect 2048 51755 2116 51811
rect 2172 51755 2240 51811
rect 2296 51755 2364 51811
rect 2420 51755 2444 51811
rect 1844 51687 2444 51755
rect 1844 51631 1868 51687
rect 1924 51631 1992 51687
rect 2048 51631 2116 51687
rect 2172 51631 2240 51687
rect 2296 51631 2364 51687
rect 2420 51631 2444 51687
rect 1844 51563 2444 51631
rect 1844 51507 1868 51563
rect 1924 51507 1992 51563
rect 2048 51507 2116 51563
rect 2172 51507 2240 51563
rect 2296 51507 2364 51563
rect 2420 51507 2444 51563
rect 1844 34614 2444 51507
rect 1844 34558 1930 34614
rect 1986 34558 2054 34614
rect 2110 34558 2178 34614
rect 2234 34558 2302 34614
rect 2358 34558 2444 34614
rect 1844 34490 2444 34558
rect 1844 34434 1930 34490
rect 1986 34434 2054 34490
rect 2110 34434 2178 34490
rect 2234 34434 2302 34490
rect 2358 34434 2444 34490
rect 1844 34366 2444 34434
rect 1844 34310 1930 34366
rect 1986 34310 2054 34366
rect 2110 34310 2178 34366
rect 2234 34310 2302 34366
rect 2358 34310 2444 34366
rect 1844 34242 2444 34310
rect 1844 34186 1930 34242
rect 1986 34186 2054 34242
rect 2110 34186 2178 34242
rect 2234 34186 2302 34242
rect 2358 34186 2444 34242
rect 1844 32240 2444 34186
rect 1844 32184 1930 32240
rect 1986 32184 2054 32240
rect 2110 32184 2178 32240
rect 2234 32184 2302 32240
rect 2358 32184 2444 32240
rect 1844 32116 2444 32184
rect 1844 32060 1930 32116
rect 1986 32060 2054 32116
rect 2110 32060 2178 32116
rect 2234 32060 2302 32116
rect 2358 32060 2444 32116
rect 1844 30440 2444 32060
rect 1844 30384 1930 30440
rect 1986 30384 2054 30440
rect 2110 30384 2178 30440
rect 2234 30384 2302 30440
rect 2358 30384 2444 30440
rect 1844 30316 2444 30384
rect 1844 30260 1930 30316
rect 1986 30260 2054 30316
rect 2110 30260 2178 30316
rect 2234 30260 2302 30316
rect 2358 30260 2444 30316
rect 1844 28640 2444 30260
rect 1844 28584 1930 28640
rect 1986 28584 2054 28640
rect 2110 28584 2178 28640
rect 2234 28584 2302 28640
rect 2358 28584 2444 28640
rect 1844 28516 2444 28584
rect 1844 28460 1930 28516
rect 1986 28460 2054 28516
rect 2110 28460 2178 28516
rect 2234 28460 2302 28516
rect 2358 28460 2444 28516
rect 1844 26840 2444 28460
rect 1844 26784 1930 26840
rect 1986 26784 2054 26840
rect 2110 26784 2178 26840
rect 2234 26784 2302 26840
rect 2358 26784 2444 26840
rect 1844 26716 2444 26784
rect 1844 26660 1930 26716
rect 1986 26660 2054 26716
rect 2110 26660 2178 26716
rect 2234 26660 2302 26716
rect 2358 26660 2444 26716
rect 1844 25040 2444 26660
rect 1844 24984 1930 25040
rect 1986 24984 2054 25040
rect 2110 24984 2178 25040
rect 2234 24984 2302 25040
rect 2358 24984 2444 25040
rect 1844 24916 2444 24984
rect 1844 24860 1930 24916
rect 1986 24860 2054 24916
rect 2110 24860 2178 24916
rect 2234 24860 2302 24916
rect 2358 24860 2444 24916
rect 1844 23240 2444 24860
rect 1844 23184 1930 23240
rect 1986 23184 2054 23240
rect 2110 23184 2178 23240
rect 2234 23184 2302 23240
rect 2358 23184 2444 23240
rect 1844 23116 2444 23184
rect 1844 23060 1930 23116
rect 1986 23060 2054 23116
rect 2110 23060 2178 23116
rect 2234 23060 2302 23116
rect 2358 23060 2444 23116
rect 1844 21440 2444 23060
rect 1844 21384 1930 21440
rect 1986 21384 2054 21440
rect 2110 21384 2178 21440
rect 2234 21384 2302 21440
rect 2358 21384 2444 21440
rect 1844 21316 2444 21384
rect 1844 21260 1930 21316
rect 1986 21260 2054 21316
rect 2110 21260 2178 21316
rect 2234 21260 2302 21316
rect 2358 21260 2444 21316
rect 1844 19640 2444 21260
rect 1844 19584 1930 19640
rect 1986 19584 2054 19640
rect 2110 19584 2178 19640
rect 2234 19584 2302 19640
rect 2358 19584 2444 19640
rect 1844 19516 2444 19584
rect 1844 19460 1930 19516
rect 1986 19460 2054 19516
rect 2110 19460 2178 19516
rect 2234 19460 2302 19516
rect 2358 19460 2444 19516
rect 1844 17840 2444 19460
rect 1844 17784 1930 17840
rect 1986 17784 2054 17840
rect 2110 17784 2178 17840
rect 2234 17784 2302 17840
rect 2358 17784 2444 17840
rect 1844 17716 2444 17784
rect 1844 17660 1930 17716
rect 1986 17660 2054 17716
rect 2110 17660 2178 17716
rect 2234 17660 2302 17716
rect 2358 17660 2444 17716
rect 1844 16040 2444 17660
rect 1844 15984 1930 16040
rect 1986 15984 2054 16040
rect 2110 15984 2178 16040
rect 2234 15984 2302 16040
rect 2358 15984 2444 16040
rect 1844 15916 2444 15984
rect 1844 15860 1930 15916
rect 1986 15860 2054 15916
rect 2110 15860 2178 15916
rect 2234 15860 2302 15916
rect 2358 15860 2444 15916
rect 1844 14240 2444 15860
rect 1844 14184 1930 14240
rect 1986 14184 2054 14240
rect 2110 14184 2178 14240
rect 2234 14184 2302 14240
rect 2358 14184 2444 14240
rect 1844 14116 2444 14184
rect 1844 14060 1930 14116
rect 1986 14060 2054 14116
rect 2110 14060 2178 14116
rect 2234 14060 2302 14116
rect 2358 14060 2444 14116
rect 1844 12440 2444 14060
rect 1844 12384 1930 12440
rect 1986 12384 2054 12440
rect 2110 12384 2178 12440
rect 2234 12384 2302 12440
rect 2358 12384 2444 12440
rect 1844 12316 2444 12384
rect 1844 12260 1930 12316
rect 1986 12260 2054 12316
rect 2110 12260 2178 12316
rect 2234 12260 2302 12316
rect 2358 12260 2444 12316
rect 1844 10640 2444 12260
rect 1844 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2444 10640
rect 1844 10516 2444 10584
rect 1844 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2444 10516
rect 1844 8840 2444 10460
rect 1844 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2444 8840
rect 1844 8716 2444 8784
rect 1844 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2444 8716
rect 1844 7040 2444 8660
rect 1844 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2444 7040
rect 1844 6916 2444 6984
rect 1844 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2444 6916
rect 1844 5240 2444 6860
rect 1844 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2444 5240
rect 1844 5116 2444 5184
rect 1844 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2444 5116
rect 1844 3440 2444 5060
rect 1844 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2444 3440
rect 1844 3316 2444 3384
rect 1844 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2444 3316
rect 1844 3136 2444 3260
rect 85726 60991 86326 66640
rect 85726 60935 85750 60991
rect 85806 60935 85874 60991
rect 85930 60935 85998 60991
rect 86054 60935 86122 60991
rect 86178 60935 86246 60991
rect 86302 60935 86326 60991
rect 85726 60867 86326 60935
rect 85726 60811 85750 60867
rect 85806 60811 85874 60867
rect 85930 60811 85998 60867
rect 86054 60811 86122 60867
rect 86178 60811 86246 60867
rect 86302 60811 86326 60867
rect 85726 60743 86326 60811
rect 85726 60687 85750 60743
rect 85806 60687 85874 60743
rect 85930 60687 85998 60743
rect 86054 60687 86122 60743
rect 86178 60687 86246 60743
rect 86302 60687 86326 60743
rect 85726 60619 86326 60687
rect 85726 60563 85750 60619
rect 85806 60563 85874 60619
rect 85930 60563 85998 60619
rect 86054 60563 86122 60619
rect 86178 60563 86246 60619
rect 86302 60563 86326 60619
rect 85726 60495 86326 60563
rect 85726 60439 85750 60495
rect 85806 60439 85874 60495
rect 85930 60439 85998 60495
rect 86054 60439 86122 60495
rect 86178 60439 86246 60495
rect 86302 60439 86326 60495
rect 85726 60371 86326 60439
rect 85726 60315 85750 60371
rect 85806 60315 85874 60371
rect 85930 60315 85998 60371
rect 86054 60315 86122 60371
rect 86178 60315 86246 60371
rect 86302 60315 86326 60371
rect 85726 60247 86326 60315
rect 85726 60191 85750 60247
rect 85806 60191 85874 60247
rect 85930 60191 85998 60247
rect 86054 60191 86122 60247
rect 86178 60191 86246 60247
rect 86302 60191 86326 60247
rect 85726 60123 86326 60191
rect 85726 60067 85750 60123
rect 85806 60067 85874 60123
rect 85930 60067 85998 60123
rect 86054 60067 86122 60123
rect 86178 60067 86246 60123
rect 86302 60067 86326 60123
rect 85726 59999 86326 60067
rect 85726 59943 85750 59999
rect 85806 59943 85874 59999
rect 85930 59943 85998 59999
rect 86054 59943 86122 59999
rect 86178 59943 86246 59999
rect 86302 59943 86326 59999
rect 85726 59875 86326 59943
rect 85726 59819 85750 59875
rect 85806 59819 85874 59875
rect 85930 59819 85998 59875
rect 86054 59819 86122 59875
rect 86178 59819 86246 59875
rect 86302 59819 86326 59875
rect 85726 59751 86326 59819
rect 85726 59695 85750 59751
rect 85806 59695 85874 59751
rect 85930 59695 85998 59751
rect 86054 59695 86122 59751
rect 86178 59695 86246 59751
rect 86302 59695 86326 59751
rect 85726 57089 86326 59695
rect 85726 57033 85750 57089
rect 85806 57033 85874 57089
rect 85930 57033 85998 57089
rect 86054 57033 86122 57089
rect 86178 57033 86246 57089
rect 86302 57033 86326 57089
rect 85726 56965 86326 57033
rect 85726 56909 85750 56965
rect 85806 56909 85874 56965
rect 85930 56909 85998 56965
rect 86054 56909 86122 56965
rect 86178 56909 86246 56965
rect 86302 56909 86326 56965
rect 85726 56841 86326 56909
rect 85726 56785 85750 56841
rect 85806 56785 85874 56841
rect 85930 56785 85998 56841
rect 86054 56785 86122 56841
rect 86178 56785 86246 56841
rect 86302 56785 86326 56841
rect 85726 56717 86326 56785
rect 85726 56661 85750 56717
rect 85806 56661 85874 56717
rect 85930 56661 85998 56717
rect 86054 56661 86122 56717
rect 86178 56661 86246 56717
rect 86302 56661 86326 56717
rect 85726 56593 86326 56661
rect 85726 56537 85750 56593
rect 85806 56537 85874 56593
rect 85930 56537 85998 56593
rect 86054 56537 86122 56593
rect 86178 56537 86246 56593
rect 86302 56537 86326 56593
rect 85726 56469 86326 56537
rect 85726 56413 85750 56469
rect 85806 56413 85874 56469
rect 85930 56413 85998 56469
rect 86054 56413 86122 56469
rect 86178 56413 86246 56469
rect 86302 56413 86326 56469
rect 85726 56345 86326 56413
rect 85726 56289 85750 56345
rect 85806 56289 85874 56345
rect 85930 56289 85998 56345
rect 86054 56289 86122 56345
rect 86178 56289 86246 56345
rect 86302 56289 86326 56345
rect 85726 56221 86326 56289
rect 85726 56165 85750 56221
rect 85806 56165 85874 56221
rect 85930 56165 85998 56221
rect 86054 56165 86122 56221
rect 86178 56165 86246 56221
rect 86302 56165 86326 56221
rect 85726 56097 86326 56165
rect 85726 56041 85750 56097
rect 85806 56041 85874 56097
rect 85930 56041 85998 56097
rect 86054 56041 86122 56097
rect 86178 56041 86246 56097
rect 86302 56041 86326 56097
rect 85726 55973 86326 56041
rect 85726 55917 85750 55973
rect 85806 55917 85874 55973
rect 85930 55917 85998 55973
rect 86054 55917 86122 55973
rect 86178 55917 86246 55973
rect 86302 55917 86326 55973
rect 85726 55849 86326 55917
rect 85726 55793 85750 55849
rect 85806 55793 85874 55849
rect 85930 55793 85998 55849
rect 86054 55793 86122 55849
rect 86178 55793 86246 55849
rect 86302 55793 86326 55849
rect 85726 55725 86326 55793
rect 85726 55669 85750 55725
rect 85806 55669 85874 55725
rect 85930 55669 85998 55725
rect 86054 55669 86122 55725
rect 86178 55669 86246 55725
rect 86302 55669 86326 55725
rect 85726 55601 86326 55669
rect 85726 55545 85750 55601
rect 85806 55545 85874 55601
rect 85930 55545 85998 55601
rect 86054 55545 86122 55601
rect 86178 55545 86246 55601
rect 86302 55545 86326 55601
rect 85726 55477 86326 55545
rect 85726 55421 85750 55477
rect 85806 55421 85874 55477
rect 85930 55421 85998 55477
rect 86054 55421 86122 55477
rect 86178 55421 86246 55477
rect 86302 55421 86326 55477
rect 85726 55353 86326 55421
rect 85726 55297 85750 55353
rect 85806 55297 85874 55353
rect 85930 55297 85998 55353
rect 86054 55297 86122 55353
rect 86178 55297 86246 55353
rect 86302 55297 86326 55353
rect 85726 55229 86326 55297
rect 85726 55173 85750 55229
rect 85806 55173 85874 55229
rect 85930 55173 85998 55229
rect 86054 55173 86122 55229
rect 86178 55173 86246 55229
rect 86302 55173 86326 55229
rect 85726 55105 86326 55173
rect 85726 55049 85750 55105
rect 85806 55049 85874 55105
rect 85930 55049 85998 55105
rect 86054 55049 86122 55105
rect 86178 55049 86246 55105
rect 86302 55049 86326 55105
rect 85726 46200 86326 55049
rect 85726 46144 85750 46200
rect 85806 46144 85874 46200
rect 85930 46144 85998 46200
rect 86054 46144 86122 46200
rect 86178 46144 86246 46200
rect 86302 46144 86326 46200
rect 85726 46076 86326 46144
rect 85726 46020 85750 46076
rect 85806 46020 85874 46076
rect 85930 46020 85998 46076
rect 86054 46020 86122 46076
rect 86178 46020 86246 46076
rect 86302 46020 86326 46076
rect 85726 45952 86326 46020
rect 85726 45896 85750 45952
rect 85806 45896 85874 45952
rect 85930 45896 85998 45952
rect 86054 45896 86122 45952
rect 86178 45896 86246 45952
rect 86302 45896 86326 45952
rect 85726 45828 86326 45896
rect 85726 45772 85750 45828
rect 85806 45772 85874 45828
rect 85930 45772 85998 45828
rect 86054 45772 86122 45828
rect 86178 45772 86246 45828
rect 86302 45772 86326 45828
rect 85726 45704 86326 45772
rect 85726 45648 85750 45704
rect 85806 45648 85874 45704
rect 85930 45648 85998 45704
rect 86054 45648 86122 45704
rect 86178 45648 86246 45704
rect 86302 45648 86326 45704
rect 85726 45580 86326 45648
rect 85726 45524 85750 45580
rect 85806 45524 85874 45580
rect 85930 45524 85998 45580
rect 86054 45524 86122 45580
rect 86178 45524 86246 45580
rect 86302 45524 86326 45580
rect 85726 45456 86326 45524
rect 85726 45400 85750 45456
rect 85806 45400 85874 45456
rect 85930 45400 85998 45456
rect 86054 45400 86122 45456
rect 86178 45400 86246 45456
rect 86302 45400 86326 45456
rect 85726 45332 86326 45400
rect 85726 45276 85750 45332
rect 85806 45276 85874 45332
rect 85930 45276 85998 45332
rect 86054 45276 86122 45332
rect 86178 45276 86246 45332
rect 86302 45276 86326 45332
rect 85726 33264 86326 45276
rect 85726 33208 85812 33264
rect 85868 33208 85936 33264
rect 85992 33208 86060 33264
rect 86116 33208 86184 33264
rect 86240 33208 86326 33264
rect 85726 33140 86326 33208
rect 85726 33084 85812 33140
rect 85868 33084 85936 33140
rect 85992 33084 86060 33140
rect 86116 33084 86184 33140
rect 86240 33084 86326 33140
rect 85726 33016 86326 33084
rect 85726 32960 85812 33016
rect 85868 32960 85936 33016
rect 85992 32960 86060 33016
rect 86116 32960 86184 33016
rect 86240 32960 86326 33016
rect 85726 32892 86326 32960
rect 85726 32836 85812 32892
rect 85868 32836 85936 32892
rect 85992 32836 86060 32892
rect 86116 32836 86184 32892
rect 86240 32836 86326 32892
rect 85726 31464 86326 32836
rect 85726 31408 85812 31464
rect 85868 31408 85936 31464
rect 85992 31408 86060 31464
rect 86116 31408 86184 31464
rect 86240 31408 86326 31464
rect 85726 31340 86326 31408
rect 85726 31284 85812 31340
rect 85868 31284 85936 31340
rect 85992 31284 86060 31340
rect 86116 31284 86184 31340
rect 86240 31284 86326 31340
rect 85726 31216 86326 31284
rect 85726 31160 85812 31216
rect 85868 31160 85936 31216
rect 85992 31160 86060 31216
rect 86116 31160 86184 31216
rect 86240 31160 86326 31216
rect 85726 31092 86326 31160
rect 85726 31036 85812 31092
rect 85868 31036 85936 31092
rect 85992 31036 86060 31092
rect 86116 31036 86184 31092
rect 86240 31036 86326 31092
rect 85726 29664 86326 31036
rect 85726 29608 85812 29664
rect 85868 29608 85936 29664
rect 85992 29608 86060 29664
rect 86116 29608 86184 29664
rect 86240 29608 86326 29664
rect 85726 29540 86326 29608
rect 85726 29484 85812 29540
rect 85868 29484 85936 29540
rect 85992 29484 86060 29540
rect 86116 29484 86184 29540
rect 86240 29484 86326 29540
rect 85726 29416 86326 29484
rect 85726 29360 85812 29416
rect 85868 29360 85936 29416
rect 85992 29360 86060 29416
rect 86116 29360 86184 29416
rect 86240 29360 86326 29416
rect 85726 29292 86326 29360
rect 85726 29236 85812 29292
rect 85868 29236 85936 29292
rect 85992 29236 86060 29292
rect 86116 29236 86184 29292
rect 86240 29236 86326 29292
rect 85726 27864 86326 29236
rect 85726 27808 85812 27864
rect 85868 27808 85936 27864
rect 85992 27808 86060 27864
rect 86116 27808 86184 27864
rect 86240 27808 86326 27864
rect 85726 27740 86326 27808
rect 85726 27684 85812 27740
rect 85868 27684 85936 27740
rect 85992 27684 86060 27740
rect 86116 27684 86184 27740
rect 86240 27684 86326 27740
rect 85726 27616 86326 27684
rect 85726 27560 85812 27616
rect 85868 27560 85936 27616
rect 85992 27560 86060 27616
rect 86116 27560 86184 27616
rect 86240 27560 86326 27616
rect 85726 27492 86326 27560
rect 85726 27436 85812 27492
rect 85868 27436 85936 27492
rect 85992 27436 86060 27492
rect 86116 27436 86184 27492
rect 86240 27436 86326 27492
rect 85726 26064 86326 27436
rect 85726 26008 85812 26064
rect 85868 26008 85936 26064
rect 85992 26008 86060 26064
rect 86116 26008 86184 26064
rect 86240 26008 86326 26064
rect 85726 25940 86326 26008
rect 85726 25884 85812 25940
rect 85868 25884 85936 25940
rect 85992 25884 86060 25940
rect 86116 25884 86184 25940
rect 86240 25884 86326 25940
rect 85726 25816 86326 25884
rect 85726 25760 85812 25816
rect 85868 25760 85936 25816
rect 85992 25760 86060 25816
rect 86116 25760 86184 25816
rect 86240 25760 86326 25816
rect 85726 25692 86326 25760
rect 85726 25636 85812 25692
rect 85868 25636 85936 25692
rect 85992 25636 86060 25692
rect 86116 25636 86184 25692
rect 86240 25636 86326 25692
rect 85726 24264 86326 25636
rect 85726 24208 85812 24264
rect 85868 24208 85936 24264
rect 85992 24208 86060 24264
rect 86116 24208 86184 24264
rect 86240 24208 86326 24264
rect 85726 24140 86326 24208
rect 85726 24084 85812 24140
rect 85868 24084 85936 24140
rect 85992 24084 86060 24140
rect 86116 24084 86184 24140
rect 86240 24084 86326 24140
rect 85726 24016 86326 24084
rect 85726 23960 85812 24016
rect 85868 23960 85936 24016
rect 85992 23960 86060 24016
rect 86116 23960 86184 24016
rect 86240 23960 86326 24016
rect 85726 23892 86326 23960
rect 85726 23836 85812 23892
rect 85868 23836 85936 23892
rect 85992 23836 86060 23892
rect 86116 23836 86184 23892
rect 86240 23836 86326 23892
rect 85726 22464 86326 23836
rect 85726 22408 85812 22464
rect 85868 22408 85936 22464
rect 85992 22408 86060 22464
rect 86116 22408 86184 22464
rect 86240 22408 86326 22464
rect 85726 22340 86326 22408
rect 85726 22284 85812 22340
rect 85868 22284 85936 22340
rect 85992 22284 86060 22340
rect 86116 22284 86184 22340
rect 86240 22284 86326 22340
rect 85726 22216 86326 22284
rect 85726 22160 85812 22216
rect 85868 22160 85936 22216
rect 85992 22160 86060 22216
rect 86116 22160 86184 22216
rect 86240 22160 86326 22216
rect 85726 22092 86326 22160
rect 85726 22036 85812 22092
rect 85868 22036 85936 22092
rect 85992 22036 86060 22092
rect 86116 22036 86184 22092
rect 86240 22036 86326 22092
rect 85726 20664 86326 22036
rect 85726 20608 85812 20664
rect 85868 20608 85936 20664
rect 85992 20608 86060 20664
rect 86116 20608 86184 20664
rect 86240 20608 86326 20664
rect 85726 20540 86326 20608
rect 85726 20484 85812 20540
rect 85868 20484 85936 20540
rect 85992 20484 86060 20540
rect 86116 20484 86184 20540
rect 86240 20484 86326 20540
rect 85726 20416 86326 20484
rect 85726 20360 85812 20416
rect 85868 20360 85936 20416
rect 85992 20360 86060 20416
rect 86116 20360 86184 20416
rect 86240 20360 86326 20416
rect 85726 20292 86326 20360
rect 85726 20236 85812 20292
rect 85868 20236 85936 20292
rect 85992 20236 86060 20292
rect 86116 20236 86184 20292
rect 86240 20236 86326 20292
rect 85726 18864 86326 20236
rect 85726 18808 85812 18864
rect 85868 18808 85936 18864
rect 85992 18808 86060 18864
rect 86116 18808 86184 18864
rect 86240 18808 86326 18864
rect 85726 18740 86326 18808
rect 85726 18684 85812 18740
rect 85868 18684 85936 18740
rect 85992 18684 86060 18740
rect 86116 18684 86184 18740
rect 86240 18684 86326 18740
rect 85726 18616 86326 18684
rect 85726 18560 85812 18616
rect 85868 18560 85936 18616
rect 85992 18560 86060 18616
rect 86116 18560 86184 18616
rect 86240 18560 86326 18616
rect 85726 18492 86326 18560
rect 85726 18436 85812 18492
rect 85868 18436 85936 18492
rect 85992 18436 86060 18492
rect 86116 18436 86184 18492
rect 86240 18436 86326 18492
rect 85726 17064 86326 18436
rect 85726 17008 85812 17064
rect 85868 17008 85936 17064
rect 85992 17008 86060 17064
rect 86116 17008 86184 17064
rect 86240 17008 86326 17064
rect 85726 16940 86326 17008
rect 85726 16884 85812 16940
rect 85868 16884 85936 16940
rect 85992 16884 86060 16940
rect 86116 16884 86184 16940
rect 86240 16884 86326 16940
rect 85726 16816 86326 16884
rect 85726 16760 85812 16816
rect 85868 16760 85936 16816
rect 85992 16760 86060 16816
rect 86116 16760 86184 16816
rect 86240 16760 86326 16816
rect 85726 16692 86326 16760
rect 85726 16636 85812 16692
rect 85868 16636 85936 16692
rect 85992 16636 86060 16692
rect 86116 16636 86184 16692
rect 86240 16636 86326 16692
rect 85726 15264 86326 16636
rect 85726 15208 85812 15264
rect 85868 15208 85936 15264
rect 85992 15208 86060 15264
rect 86116 15208 86184 15264
rect 86240 15208 86326 15264
rect 85726 15140 86326 15208
rect 85726 15084 85812 15140
rect 85868 15084 85936 15140
rect 85992 15084 86060 15140
rect 86116 15084 86184 15140
rect 86240 15084 86326 15140
rect 85726 15016 86326 15084
rect 85726 14960 85812 15016
rect 85868 14960 85936 15016
rect 85992 14960 86060 15016
rect 86116 14960 86184 15016
rect 86240 14960 86326 15016
rect 85726 14892 86326 14960
rect 85726 14836 85812 14892
rect 85868 14836 85936 14892
rect 85992 14836 86060 14892
rect 86116 14836 86184 14892
rect 86240 14836 86326 14892
rect 85726 13464 86326 14836
rect 85726 13408 85812 13464
rect 85868 13408 85936 13464
rect 85992 13408 86060 13464
rect 86116 13408 86184 13464
rect 86240 13408 86326 13464
rect 85726 13340 86326 13408
rect 85726 13284 85812 13340
rect 85868 13284 85936 13340
rect 85992 13284 86060 13340
rect 86116 13284 86184 13340
rect 86240 13284 86326 13340
rect 85726 13216 86326 13284
rect 85726 13160 85812 13216
rect 85868 13160 85936 13216
rect 85992 13160 86060 13216
rect 86116 13160 86184 13216
rect 86240 13160 86326 13216
rect 85726 13092 86326 13160
rect 85726 13036 85812 13092
rect 85868 13036 85936 13092
rect 85992 13036 86060 13092
rect 86116 13036 86184 13092
rect 86240 13036 86326 13092
rect 85726 11664 86326 13036
rect 85726 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86326 11664
rect 85726 11540 86326 11608
rect 85726 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86326 11540
rect 85726 11416 86326 11484
rect 85726 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86326 11416
rect 85726 11292 86326 11360
rect 85726 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86326 11292
rect 85726 9864 86326 11236
rect 85726 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86326 9864
rect 85726 9740 86326 9808
rect 85726 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86326 9740
rect 85726 9616 86326 9684
rect 85726 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86326 9616
rect 85726 9492 86326 9560
rect 85726 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86326 9492
rect 85726 8064 86326 9436
rect 85726 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86326 8064
rect 85726 7940 86326 8008
rect 85726 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86326 7940
rect 85726 7816 86326 7884
rect 85726 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86326 7816
rect 85726 7692 86326 7760
rect 85726 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86326 7692
rect 85726 6264 86326 7636
rect 85726 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86326 6264
rect 85726 6140 86326 6208
rect 85726 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86326 6140
rect 85726 6016 86326 6084
rect 85726 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86326 6016
rect 85726 5892 86326 5960
rect 85726 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86326 5892
rect 85726 4464 86326 5836
rect 85726 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86326 4464
rect 85726 4340 86326 4408
rect 85726 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86326 4340
rect 85726 4216 86326 4284
rect 85726 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86326 4216
rect 85726 4092 86326 4160
rect 85726 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86326 4092
rect 85726 3136 86326 4036
rect 86526 66608 87126 66640
rect 86526 66552 86550 66608
rect 86606 66552 86674 66608
rect 86730 66552 86798 66608
rect 86854 66552 86922 66608
rect 86978 66552 87046 66608
rect 87102 66552 87126 66608
rect 86526 66484 87126 66552
rect 86526 66428 86550 66484
rect 86606 66428 86674 66484
rect 86730 66428 86798 66484
rect 86854 66428 86922 66484
rect 86978 66428 87046 66484
rect 87102 66428 87126 66484
rect 86526 66360 87126 66428
rect 86526 66304 86550 66360
rect 86606 66304 86674 66360
rect 86730 66304 86798 66360
rect 86854 66304 86922 66360
rect 86978 66304 87046 66360
rect 87102 66304 87126 66360
rect 86526 66236 87126 66304
rect 86526 66180 86550 66236
rect 86606 66180 86674 66236
rect 86730 66180 86798 66236
rect 86854 66180 86922 66236
rect 86978 66180 87046 66236
rect 87102 66180 87126 66236
rect 86526 66112 87126 66180
rect 86526 66056 86550 66112
rect 86606 66056 86674 66112
rect 86730 66056 86798 66112
rect 86854 66056 86922 66112
rect 86978 66056 87046 66112
rect 87102 66056 87126 66112
rect 86526 65988 87126 66056
rect 86526 65932 86550 65988
rect 86606 65932 86674 65988
rect 86730 65932 86798 65988
rect 86854 65932 86922 65988
rect 86978 65932 87046 65988
rect 87102 65932 87126 65988
rect 86526 65864 87126 65932
rect 86526 65808 86550 65864
rect 86606 65808 86674 65864
rect 86730 65808 86798 65864
rect 86854 65808 86922 65864
rect 86978 65808 87046 65864
rect 87102 65808 87126 65864
rect 86526 65740 87126 65808
rect 86526 65684 86550 65740
rect 86606 65684 86674 65740
rect 86730 65684 86798 65740
rect 86854 65684 86922 65740
rect 86978 65684 87046 65740
rect 87102 65684 87126 65740
rect 86526 65616 87126 65684
rect 86526 65560 86550 65616
rect 86606 65560 86674 65616
rect 86730 65560 86798 65616
rect 86854 65560 86922 65616
rect 86978 65560 87046 65616
rect 87102 65560 87126 65616
rect 86526 65492 87126 65560
rect 86526 65436 86550 65492
rect 86606 65436 86674 65492
rect 86730 65436 86798 65492
rect 86854 65436 86922 65492
rect 86978 65436 87046 65492
rect 87102 65436 87126 65492
rect 86526 63391 87126 65436
rect 86526 63335 86550 63391
rect 86606 63335 86674 63391
rect 86730 63335 86798 63391
rect 86854 63335 86922 63391
rect 86978 63335 87046 63391
rect 87102 63335 87126 63391
rect 86526 63267 87126 63335
rect 86526 63211 86550 63267
rect 86606 63211 86674 63267
rect 86730 63211 86798 63267
rect 86854 63211 86922 63267
rect 86978 63211 87046 63267
rect 87102 63211 87126 63267
rect 86526 63143 87126 63211
rect 86526 63087 86550 63143
rect 86606 63087 86674 63143
rect 86730 63087 86798 63143
rect 86854 63087 86922 63143
rect 86978 63087 87046 63143
rect 87102 63087 87126 63143
rect 86526 63019 87126 63087
rect 86526 62963 86550 63019
rect 86606 62963 86674 63019
rect 86730 62963 86798 63019
rect 86854 62963 86922 63019
rect 86978 62963 87046 63019
rect 87102 62963 87126 63019
rect 86526 62895 87126 62963
rect 86526 62839 86550 62895
rect 86606 62839 86674 62895
rect 86730 62839 86798 62895
rect 86854 62839 86922 62895
rect 86978 62839 87046 62895
rect 87102 62839 87126 62895
rect 86526 62771 87126 62839
rect 86526 62715 86550 62771
rect 86606 62715 86674 62771
rect 86730 62715 86798 62771
rect 86854 62715 86922 62771
rect 86978 62715 87046 62771
rect 87102 62715 87126 62771
rect 86526 62647 87126 62715
rect 86526 62591 86550 62647
rect 86606 62591 86674 62647
rect 86730 62591 86798 62647
rect 86854 62591 86922 62647
rect 86978 62591 87046 62647
rect 87102 62591 87126 62647
rect 86526 62523 87126 62591
rect 86526 62467 86550 62523
rect 86606 62467 86674 62523
rect 86730 62467 86798 62523
rect 86854 62467 86922 62523
rect 86978 62467 87046 62523
rect 87102 62467 87126 62523
rect 86526 62399 87126 62467
rect 86526 62343 86550 62399
rect 86606 62343 86674 62399
rect 86730 62343 86798 62399
rect 86854 62343 86922 62399
rect 86978 62343 87046 62399
rect 87102 62343 87126 62399
rect 86526 62275 87126 62343
rect 86526 62219 86550 62275
rect 86606 62219 86674 62275
rect 86730 62219 86798 62275
rect 86854 62219 86922 62275
rect 86978 62219 87046 62275
rect 87102 62219 87126 62275
rect 86526 62151 87126 62219
rect 86526 62095 86550 62151
rect 86606 62095 86674 62151
rect 86730 62095 86798 62151
rect 86854 62095 86922 62151
rect 86978 62095 87046 62151
rect 87102 62095 87126 62151
rect 86526 62027 87126 62095
rect 86526 61971 86550 62027
rect 86606 61971 86674 62027
rect 86730 61971 86798 62027
rect 86854 61971 86922 62027
rect 86978 61971 87046 62027
rect 87102 61971 87126 62027
rect 86526 61903 87126 61971
rect 86526 61847 86550 61903
rect 86606 61847 86674 61903
rect 86730 61847 86798 61903
rect 86854 61847 86922 61903
rect 86978 61847 87046 61903
rect 87102 61847 87126 61903
rect 86526 61779 87126 61847
rect 86526 61723 86550 61779
rect 86606 61723 86674 61779
rect 86730 61723 86798 61779
rect 86854 61723 86922 61779
rect 86978 61723 87046 61779
rect 87102 61723 87126 61779
rect 86526 61655 87126 61723
rect 86526 61599 86550 61655
rect 86606 61599 86674 61655
rect 86730 61599 86798 61655
rect 86854 61599 86922 61655
rect 86978 61599 87046 61655
rect 87102 61599 87126 61655
rect 86526 54787 87126 61599
rect 86526 54731 86550 54787
rect 86606 54731 86674 54787
rect 86730 54731 86798 54787
rect 86854 54731 86922 54787
rect 86978 54731 87046 54787
rect 87102 54731 87126 54787
rect 86526 54663 87126 54731
rect 86526 54607 86550 54663
rect 86606 54607 86674 54663
rect 86730 54607 86798 54663
rect 86854 54607 86922 54663
rect 86978 54607 87046 54663
rect 87102 54607 87126 54663
rect 86526 54539 87126 54607
rect 86526 54483 86550 54539
rect 86606 54483 86674 54539
rect 86730 54483 86798 54539
rect 86854 54483 86922 54539
rect 86978 54483 87046 54539
rect 87102 54483 87126 54539
rect 86526 54415 87126 54483
rect 86526 54359 86550 54415
rect 86606 54359 86674 54415
rect 86730 54359 86798 54415
rect 86854 54359 86922 54415
rect 86978 54359 87046 54415
rect 87102 54359 87126 54415
rect 86526 54291 87126 54359
rect 86526 54235 86550 54291
rect 86606 54235 86674 54291
rect 86730 54235 86798 54291
rect 86854 54235 86922 54291
rect 86978 54235 87046 54291
rect 87102 54235 87126 54291
rect 86526 54167 87126 54235
rect 86526 54111 86550 54167
rect 86606 54111 86674 54167
rect 86730 54111 86798 54167
rect 86854 54111 86922 54167
rect 86978 54111 87046 54167
rect 87102 54111 87126 54167
rect 86526 54043 87126 54111
rect 86526 53987 86550 54043
rect 86606 53987 86674 54043
rect 86730 53987 86798 54043
rect 86854 53987 86922 54043
rect 86978 53987 87046 54043
rect 87102 53987 87126 54043
rect 86526 53919 87126 53987
rect 86526 53863 86550 53919
rect 86606 53863 86674 53919
rect 86730 53863 86798 53919
rect 86854 53863 86922 53919
rect 86978 53863 87046 53919
rect 87102 53863 87126 53919
rect 86526 53795 87126 53863
rect 86526 53739 86550 53795
rect 86606 53739 86674 53795
rect 86730 53739 86798 53795
rect 86854 53739 86922 53795
rect 86978 53739 87046 53795
rect 87102 53739 87126 53795
rect 86526 53671 87126 53739
rect 86526 53615 86550 53671
rect 86606 53615 86674 53671
rect 86730 53615 86798 53671
rect 86854 53615 86922 53671
rect 86978 53615 87046 53671
rect 87102 53615 87126 53671
rect 86526 53547 87126 53615
rect 86526 53491 86550 53547
rect 86606 53491 86674 53547
rect 86730 53491 86798 53547
rect 86854 53491 86922 53547
rect 86978 53491 87046 53547
rect 87102 53491 87126 53547
rect 86526 53423 87126 53491
rect 86526 53367 86550 53423
rect 86606 53367 86674 53423
rect 86730 53367 86798 53423
rect 86854 53367 86922 53423
rect 86978 53367 87046 53423
rect 87102 53367 87126 53423
rect 86526 53299 87126 53367
rect 86526 53243 86550 53299
rect 86606 53243 86674 53299
rect 86730 53243 86798 53299
rect 86854 53243 86922 53299
rect 86978 53243 87046 53299
rect 87102 53243 87126 53299
rect 86526 53175 87126 53243
rect 86526 53119 86550 53175
rect 86606 53119 86674 53175
rect 86730 53119 86798 53175
rect 86854 53119 86922 53175
rect 86978 53119 87046 53175
rect 87102 53119 87126 53175
rect 86526 53051 87126 53119
rect 86526 52995 86550 53051
rect 86606 52995 86674 53051
rect 86730 52995 86798 53051
rect 86854 52995 86922 53051
rect 86978 52995 87046 53051
rect 87102 52995 87126 53051
rect 86526 52927 87126 52995
rect 86526 52871 86550 52927
rect 86606 52871 86674 52927
rect 86730 52871 86798 52927
rect 86854 52871 86922 52927
rect 86978 52871 87046 52927
rect 87102 52871 87126 52927
rect 86526 52803 87126 52871
rect 86526 52747 86550 52803
rect 86606 52747 86674 52803
rect 86730 52747 86798 52803
rect 86854 52747 86922 52803
rect 86978 52747 87046 52803
rect 87102 52747 87126 52803
rect 86526 52679 87126 52747
rect 86526 52623 86550 52679
rect 86606 52623 86674 52679
rect 86730 52623 86798 52679
rect 86854 52623 86922 52679
rect 86978 52623 87046 52679
rect 87102 52623 87126 52679
rect 86526 52555 87126 52623
rect 86526 52499 86550 52555
rect 86606 52499 86674 52555
rect 86730 52499 86798 52555
rect 86854 52499 86922 52555
rect 86978 52499 87046 52555
rect 87102 52499 87126 52555
rect 86526 52431 87126 52499
rect 86526 52375 86550 52431
rect 86606 52375 86674 52431
rect 86730 52375 86798 52431
rect 86854 52375 86922 52431
rect 86978 52375 87046 52431
rect 87102 52375 87126 52431
rect 86526 52307 87126 52375
rect 86526 52251 86550 52307
rect 86606 52251 86674 52307
rect 86730 52251 86798 52307
rect 86854 52251 86922 52307
rect 86978 52251 87046 52307
rect 87102 52251 87126 52307
rect 86526 52183 87126 52251
rect 86526 52127 86550 52183
rect 86606 52127 86674 52183
rect 86730 52127 86798 52183
rect 86854 52127 86922 52183
rect 86978 52127 87046 52183
rect 87102 52127 87126 52183
rect 86526 52059 87126 52127
rect 86526 52003 86550 52059
rect 86606 52003 86674 52059
rect 86730 52003 86798 52059
rect 86854 52003 86922 52059
rect 86978 52003 87046 52059
rect 87102 52003 87126 52059
rect 86526 51935 87126 52003
rect 86526 51879 86550 51935
rect 86606 51879 86674 51935
rect 86730 51879 86798 51935
rect 86854 51879 86922 51935
rect 86978 51879 87046 51935
rect 87102 51879 87126 51935
rect 86526 51811 87126 51879
rect 86526 51755 86550 51811
rect 86606 51755 86674 51811
rect 86730 51755 86798 51811
rect 86854 51755 86922 51811
rect 86978 51755 87046 51811
rect 87102 51755 87126 51811
rect 86526 51687 87126 51755
rect 86526 51631 86550 51687
rect 86606 51631 86674 51687
rect 86730 51631 86798 51687
rect 86854 51631 86922 51687
rect 86978 51631 87046 51687
rect 87102 51631 87126 51687
rect 86526 51563 87126 51631
rect 86526 51507 86550 51563
rect 86606 51507 86674 51563
rect 86730 51507 86798 51563
rect 86854 51507 86922 51563
rect 86978 51507 87046 51563
rect 87102 51507 87126 51563
rect 86526 47856 87126 51507
rect 86526 47800 86550 47856
rect 86606 47800 86674 47856
rect 86730 47800 86798 47856
rect 86854 47800 86922 47856
rect 86978 47800 87046 47856
rect 87102 47800 87126 47856
rect 86526 47732 87126 47800
rect 86526 47676 86550 47732
rect 86606 47676 86674 47732
rect 86730 47676 86798 47732
rect 86854 47676 86922 47732
rect 86978 47676 87046 47732
rect 87102 47676 87126 47732
rect 86526 47608 87126 47676
rect 86526 47552 86550 47608
rect 86606 47552 86674 47608
rect 86730 47552 86798 47608
rect 86854 47552 86922 47608
rect 86978 47552 87046 47608
rect 87102 47552 87126 47608
rect 86526 47484 87126 47552
rect 86526 47428 86550 47484
rect 86606 47428 86674 47484
rect 86730 47428 86798 47484
rect 86854 47428 86922 47484
rect 86978 47428 87046 47484
rect 87102 47428 87126 47484
rect 86526 47360 87126 47428
rect 86526 47304 86550 47360
rect 86606 47304 86674 47360
rect 86730 47304 86798 47360
rect 86854 47304 86922 47360
rect 86978 47304 87046 47360
rect 87102 47304 87126 47360
rect 86526 47236 87126 47304
rect 86526 47180 86550 47236
rect 86606 47180 86674 47236
rect 86730 47180 86798 47236
rect 86854 47180 86922 47236
rect 86978 47180 87046 47236
rect 87102 47180 87126 47236
rect 86526 47112 87126 47180
rect 86526 47056 86550 47112
rect 86606 47056 86674 47112
rect 86730 47056 86798 47112
rect 86854 47056 86922 47112
rect 86978 47056 87046 47112
rect 87102 47056 87126 47112
rect 86526 46988 87126 47056
rect 86526 46932 86550 46988
rect 86606 46932 86674 46988
rect 86730 46932 86798 46988
rect 86854 46932 86922 46988
rect 86978 46932 87046 46988
rect 87102 46932 87126 46988
rect 86526 34459 87126 46932
rect 86526 34403 86612 34459
rect 86668 34403 86736 34459
rect 86792 34403 86860 34459
rect 86916 34403 86984 34459
rect 87040 34403 87126 34459
rect 86526 34335 87126 34403
rect 86526 34279 86612 34335
rect 86668 34279 86736 34335
rect 86792 34279 86860 34335
rect 86916 34279 86984 34335
rect 87040 34279 87126 34335
rect 86526 34211 87126 34279
rect 86526 34155 86612 34211
rect 86668 34155 86736 34211
rect 86792 34155 86860 34211
rect 86916 34155 86984 34211
rect 87040 34155 87126 34211
rect 86526 34087 87126 34155
rect 86526 34031 86612 34087
rect 86668 34031 86736 34087
rect 86792 34031 86860 34087
rect 86916 34031 86984 34087
rect 87040 34031 87126 34087
rect 86526 32364 87126 34031
rect 86526 32308 86612 32364
rect 86668 32308 86736 32364
rect 86792 32308 86860 32364
rect 86916 32308 86984 32364
rect 87040 32308 87126 32364
rect 86526 32240 87126 32308
rect 86526 32184 86612 32240
rect 86668 32184 86736 32240
rect 86792 32184 86860 32240
rect 86916 32184 86984 32240
rect 87040 32184 87126 32240
rect 86526 32116 87126 32184
rect 86526 32060 86612 32116
rect 86668 32060 86736 32116
rect 86792 32060 86860 32116
rect 86916 32060 86984 32116
rect 87040 32060 87126 32116
rect 86526 31992 87126 32060
rect 86526 31936 86612 31992
rect 86668 31936 86736 31992
rect 86792 31936 86860 31992
rect 86916 31936 86984 31992
rect 87040 31936 87126 31992
rect 86526 30564 87126 31936
rect 86526 30508 86612 30564
rect 86668 30508 86736 30564
rect 86792 30508 86860 30564
rect 86916 30508 86984 30564
rect 87040 30508 87126 30564
rect 86526 30440 87126 30508
rect 86526 30384 86612 30440
rect 86668 30384 86736 30440
rect 86792 30384 86860 30440
rect 86916 30384 86984 30440
rect 87040 30384 87126 30440
rect 86526 30316 87126 30384
rect 86526 30260 86612 30316
rect 86668 30260 86736 30316
rect 86792 30260 86860 30316
rect 86916 30260 86984 30316
rect 87040 30260 87126 30316
rect 86526 30192 87126 30260
rect 86526 30136 86612 30192
rect 86668 30136 86736 30192
rect 86792 30136 86860 30192
rect 86916 30136 86984 30192
rect 87040 30136 87126 30192
rect 86526 28764 87126 30136
rect 86526 28708 86612 28764
rect 86668 28708 86736 28764
rect 86792 28708 86860 28764
rect 86916 28708 86984 28764
rect 87040 28708 87126 28764
rect 86526 28640 87126 28708
rect 86526 28584 86612 28640
rect 86668 28584 86736 28640
rect 86792 28584 86860 28640
rect 86916 28584 86984 28640
rect 87040 28584 87126 28640
rect 86526 28516 87126 28584
rect 86526 28460 86612 28516
rect 86668 28460 86736 28516
rect 86792 28460 86860 28516
rect 86916 28460 86984 28516
rect 87040 28460 87126 28516
rect 86526 28392 87126 28460
rect 86526 28336 86612 28392
rect 86668 28336 86736 28392
rect 86792 28336 86860 28392
rect 86916 28336 86984 28392
rect 87040 28336 87126 28392
rect 86526 26964 87126 28336
rect 86526 26908 86612 26964
rect 86668 26908 86736 26964
rect 86792 26908 86860 26964
rect 86916 26908 86984 26964
rect 87040 26908 87126 26964
rect 86526 26840 87126 26908
rect 86526 26784 86612 26840
rect 86668 26784 86736 26840
rect 86792 26784 86860 26840
rect 86916 26784 86984 26840
rect 87040 26784 87126 26840
rect 86526 26716 87126 26784
rect 86526 26660 86612 26716
rect 86668 26660 86736 26716
rect 86792 26660 86860 26716
rect 86916 26660 86984 26716
rect 87040 26660 87126 26716
rect 86526 26592 87126 26660
rect 86526 26536 86612 26592
rect 86668 26536 86736 26592
rect 86792 26536 86860 26592
rect 86916 26536 86984 26592
rect 87040 26536 87126 26592
rect 86526 25164 87126 26536
rect 86526 25108 86612 25164
rect 86668 25108 86736 25164
rect 86792 25108 86860 25164
rect 86916 25108 86984 25164
rect 87040 25108 87126 25164
rect 86526 25040 87126 25108
rect 86526 24984 86612 25040
rect 86668 24984 86736 25040
rect 86792 24984 86860 25040
rect 86916 24984 86984 25040
rect 87040 24984 87126 25040
rect 86526 24916 87126 24984
rect 86526 24860 86612 24916
rect 86668 24860 86736 24916
rect 86792 24860 86860 24916
rect 86916 24860 86984 24916
rect 87040 24860 87126 24916
rect 86526 24792 87126 24860
rect 86526 24736 86612 24792
rect 86668 24736 86736 24792
rect 86792 24736 86860 24792
rect 86916 24736 86984 24792
rect 87040 24736 87126 24792
rect 86526 23364 87126 24736
rect 86526 23308 86612 23364
rect 86668 23308 86736 23364
rect 86792 23308 86860 23364
rect 86916 23308 86984 23364
rect 87040 23308 87126 23364
rect 86526 23240 87126 23308
rect 86526 23184 86612 23240
rect 86668 23184 86736 23240
rect 86792 23184 86860 23240
rect 86916 23184 86984 23240
rect 87040 23184 87126 23240
rect 86526 23116 87126 23184
rect 86526 23060 86612 23116
rect 86668 23060 86736 23116
rect 86792 23060 86860 23116
rect 86916 23060 86984 23116
rect 87040 23060 87126 23116
rect 86526 22992 87126 23060
rect 86526 22936 86612 22992
rect 86668 22936 86736 22992
rect 86792 22936 86860 22992
rect 86916 22936 86984 22992
rect 87040 22936 87126 22992
rect 86526 21564 87126 22936
rect 86526 21508 86612 21564
rect 86668 21508 86736 21564
rect 86792 21508 86860 21564
rect 86916 21508 86984 21564
rect 87040 21508 87126 21564
rect 86526 21440 87126 21508
rect 86526 21384 86612 21440
rect 86668 21384 86736 21440
rect 86792 21384 86860 21440
rect 86916 21384 86984 21440
rect 87040 21384 87126 21440
rect 86526 21316 87126 21384
rect 86526 21260 86612 21316
rect 86668 21260 86736 21316
rect 86792 21260 86860 21316
rect 86916 21260 86984 21316
rect 87040 21260 87126 21316
rect 86526 21192 87126 21260
rect 86526 21136 86612 21192
rect 86668 21136 86736 21192
rect 86792 21136 86860 21192
rect 86916 21136 86984 21192
rect 87040 21136 87126 21192
rect 86526 19764 87126 21136
rect 86526 19708 86612 19764
rect 86668 19708 86736 19764
rect 86792 19708 86860 19764
rect 86916 19708 86984 19764
rect 87040 19708 87126 19764
rect 86526 19640 87126 19708
rect 86526 19584 86612 19640
rect 86668 19584 86736 19640
rect 86792 19584 86860 19640
rect 86916 19584 86984 19640
rect 87040 19584 87126 19640
rect 86526 19516 87126 19584
rect 86526 19460 86612 19516
rect 86668 19460 86736 19516
rect 86792 19460 86860 19516
rect 86916 19460 86984 19516
rect 87040 19460 87126 19516
rect 86526 19392 87126 19460
rect 86526 19336 86612 19392
rect 86668 19336 86736 19392
rect 86792 19336 86860 19392
rect 86916 19336 86984 19392
rect 87040 19336 87126 19392
rect 86526 17964 87126 19336
rect 86526 17908 86612 17964
rect 86668 17908 86736 17964
rect 86792 17908 86860 17964
rect 86916 17908 86984 17964
rect 87040 17908 87126 17964
rect 86526 17840 87126 17908
rect 86526 17784 86612 17840
rect 86668 17784 86736 17840
rect 86792 17784 86860 17840
rect 86916 17784 86984 17840
rect 87040 17784 87126 17840
rect 86526 17716 87126 17784
rect 86526 17660 86612 17716
rect 86668 17660 86736 17716
rect 86792 17660 86860 17716
rect 86916 17660 86984 17716
rect 87040 17660 87126 17716
rect 86526 17592 87126 17660
rect 86526 17536 86612 17592
rect 86668 17536 86736 17592
rect 86792 17536 86860 17592
rect 86916 17536 86984 17592
rect 87040 17536 87126 17592
rect 86526 16164 87126 17536
rect 86526 16108 86612 16164
rect 86668 16108 86736 16164
rect 86792 16108 86860 16164
rect 86916 16108 86984 16164
rect 87040 16108 87126 16164
rect 86526 16040 87126 16108
rect 86526 15984 86612 16040
rect 86668 15984 86736 16040
rect 86792 15984 86860 16040
rect 86916 15984 86984 16040
rect 87040 15984 87126 16040
rect 86526 15916 87126 15984
rect 86526 15860 86612 15916
rect 86668 15860 86736 15916
rect 86792 15860 86860 15916
rect 86916 15860 86984 15916
rect 87040 15860 87126 15916
rect 86526 15792 87126 15860
rect 86526 15736 86612 15792
rect 86668 15736 86736 15792
rect 86792 15736 86860 15792
rect 86916 15736 86984 15792
rect 87040 15736 87126 15792
rect 86526 14364 87126 15736
rect 86526 14308 86612 14364
rect 86668 14308 86736 14364
rect 86792 14308 86860 14364
rect 86916 14308 86984 14364
rect 87040 14308 87126 14364
rect 86526 14240 87126 14308
rect 86526 14184 86612 14240
rect 86668 14184 86736 14240
rect 86792 14184 86860 14240
rect 86916 14184 86984 14240
rect 87040 14184 87126 14240
rect 86526 14116 87126 14184
rect 86526 14060 86612 14116
rect 86668 14060 86736 14116
rect 86792 14060 86860 14116
rect 86916 14060 86984 14116
rect 87040 14060 87126 14116
rect 86526 13992 87126 14060
rect 86526 13936 86612 13992
rect 86668 13936 86736 13992
rect 86792 13936 86860 13992
rect 86916 13936 86984 13992
rect 87040 13936 87126 13992
rect 86526 12564 87126 13936
rect 86526 12508 86612 12564
rect 86668 12508 86736 12564
rect 86792 12508 86860 12564
rect 86916 12508 86984 12564
rect 87040 12508 87126 12564
rect 86526 12440 87126 12508
rect 86526 12384 86612 12440
rect 86668 12384 86736 12440
rect 86792 12384 86860 12440
rect 86916 12384 86984 12440
rect 87040 12384 87126 12440
rect 86526 12316 87126 12384
rect 86526 12260 86612 12316
rect 86668 12260 86736 12316
rect 86792 12260 86860 12316
rect 86916 12260 86984 12316
rect 87040 12260 87126 12316
rect 86526 12192 87126 12260
rect 86526 12136 86612 12192
rect 86668 12136 86736 12192
rect 86792 12136 86860 12192
rect 86916 12136 86984 12192
rect 87040 12136 87126 12192
rect 86526 10764 87126 12136
rect 86526 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87126 10764
rect 86526 10640 87126 10708
rect 86526 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87126 10640
rect 86526 10516 87126 10584
rect 86526 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87126 10516
rect 86526 10392 87126 10460
rect 86526 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87126 10392
rect 86526 8964 87126 10336
rect 86526 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87126 8964
rect 86526 8840 87126 8908
rect 86526 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87126 8840
rect 86526 8716 87126 8784
rect 86526 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87126 8716
rect 86526 8592 87126 8660
rect 86526 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87126 8592
rect 86526 7164 87126 8536
rect 86526 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87126 7164
rect 86526 7040 87126 7108
rect 86526 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87126 7040
rect 86526 6916 87126 6984
rect 86526 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87126 6916
rect 86526 6792 87126 6860
rect 86526 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87126 6792
rect 86526 5364 87126 6736
rect 86526 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87126 5364
rect 86526 5240 87126 5308
rect 86526 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87126 5240
rect 86526 5116 87126 5184
rect 86526 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87126 5116
rect 86526 4992 87126 5060
rect 86526 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87126 4992
rect 86526 3632 87126 4936
rect 86526 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87126 3632
rect 86526 3508 87126 3576
rect 86526 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87126 3508
rect 86526 3384 87126 3452
rect 86526 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87126 3384
rect 86526 3260 87126 3328
rect 86526 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87126 3260
rect 86526 3136 87126 3204
use gf180mcu_fd_ip_sram__sram256x8m8wm1  RAM
timestamp 0
transform -1 0 87372 0 -1 69176
box 0 0 86372 68176
<< labels >>
flabel metal2 s 52944 69576 53056 70376 0 FreeSans 448 90 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 54644 69576 54756 70376 0 FreeSans 448 90 0 0 A[1]
port 1 nsew signal input
flabel metal2 s 56344 69576 56456 70376 0 FreeSans 448 90 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 30944 69576 31056 70376 0 FreeSans 448 90 0 0 A[3]
port 3 nsew signal input
flabel metal2 s 31944 69576 32056 70376 0 FreeSans 448 90 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 32744 69576 32856 70376 0 FreeSans 448 90 0 0 A[5]
port 5 nsew signal input
flabel metal2 s 33344 69576 33456 70376 0 FreeSans 448 90 0 0 A[6]
port 6 nsew signal input
flabel metal2 s 57444 69576 57556 70376 0 FreeSans 448 90 0 0 A[7]
port 7 nsew signal input
flabel metal2 s 36844 69576 36956 70376 0 FreeSans 448 90 0 0 CEN
port 8 nsew signal input
flabel metal2 s 59244 69576 59356 70376 0 FreeSans 448 90 0 0 CLK
port 9 nsew signal input
flabel metal2 s 85344 69576 85456 70376 0 FreeSans 448 90 0 0 D[0]
port 10 nsew signal input
flabel metal2 s 74944 69576 75056 70376 0 FreeSans 448 90 0 0 D[1]
port 11 nsew signal input
flabel metal2 s 73744 69576 73856 70376 0 FreeSans 448 90 0 0 D[2]
port 12 nsew signal input
flabel metal2 s 63344 69576 63456 70376 0 FreeSans 448 90 0 0 D[3]
port 13 nsew signal input
flabel metal2 s 25744 69576 25856 70376 0 FreeSans 448 90 0 0 D[4]
port 14 nsew signal input
flabel metal2 s 15444 69576 15556 70376 0 FreeSans 448 90 0 0 D[5]
port 15 nsew signal input
flabel metal2 s 14144 69576 14256 70376 0 FreeSans 448 90 0 0 D[6]
port 16 nsew signal input
flabel metal2 s 3744 69576 3856 70376 0 FreeSans 448 90 0 0 D[7]
port 17 nsew signal input
flabel metal2 s 46568 69576 46680 70376 0 FreeSans 448 90 0 0 GWEN
port 18 nsew signal input
flabel metal2 s 83844 69576 83956 70376 0 FreeSans 448 90 0 0 Q[0]
port 19 nsew signal tristate
flabel metal2 s 75644 69576 75756 70376 0 FreeSans 448 90 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 73044 69576 73156 70376 0 FreeSans 448 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal2 s 64944 69576 65056 70376 0 FreeSans 448 90 0 0 Q[3]
port 22 nsew signal tristate
flabel metal2 s 24244 69576 24356 70376 0 FreeSans 448 90 0 0 Q[4]
port 23 nsew signal tristate
flabel metal2 s 16044 69576 16156 70376 0 FreeSans 448 90 0 0 Q[5]
port 24 nsew signal tristate
flabel metal2 s 13444 69576 13556 70376 0 FreeSans 448 90 0 0 Q[6]
port 25 nsew signal tristate
flabel metal2 s 5344 69576 5456 70376 0 FreeSans 448 90 0 0 Q[7]
port 26 nsew signal tristate
flabel metal4 s 1044 3136 1644 66640 0 FreeSans 2560 90 0 0 VDD
port 27 nsew power bidirectional
flabel metal4 s 85726 3136 86326 66640 0 FreeSans 2560 90 0 0 VDD
port 27 nsew power bidirectional
flabel metal4 s 1844 3136 2444 66640 0 FreeSans 2560 90 0 0 VSS
port 28 nsew ground bidirectional
flabel metal4 s 86526 3136 87126 66640 0 FreeSans 2560 90 0 0 VSS
port 28 nsew ground bidirectional
flabel metal2 s 84644 69576 84756 70376 0 FreeSans 448 90 0 0 WEN[0]
port 29 nsew signal input
flabel metal2 s 74544 69576 74656 70376 0 FreeSans 448 90 0 0 WEN[1]
port 30 nsew signal input
flabel metal2 s 74144 69576 74256 70376 0 FreeSans 448 90 0 0 WEN[2]
port 31 nsew signal input
flabel metal2 s 63744 69576 63856 70376 0 FreeSans 448 90 0 0 WEN[3]
port 32 nsew signal input
flabel metal2 s 25044 69576 25156 70376 0 FreeSans 448 90 0 0 WEN[4]
port 33 nsew signal input
flabel metal2 s 14994 69576 15106 70376 0 FreeSans 448 90 0 0 WEN[5]
port 34 nsew signal input
flabel metal2 s 14544 69576 14656 70376 0 FreeSans 448 90 0 0 WEN[6]
port 35 nsew signal input
flabel metal2 s 4444 69576 4556 70376 0 FreeSans 448 90 0 0 WEN[7]
port 36 nsew signal input
rlabel via3 86274 60963 86274 60963 0 VDD
rlabel via3 87074 66580 87074 66580 0 VSS
rlabel metal2 53032 69328 53032 69328 0 A[0]
rlabel metal2 54712 69328 54712 69328 0 A[1]
rlabel metal2 56392 69328 56392 69328 0 A[2]
rlabel metal2 30968 69328 30968 69328 0 A[3]
rlabel metal2 32088 69174 32088 69174 0 A[4]
rlabel metal2 32816 69342 32816 69342 0 A[5]
rlabel metal2 33432 69328 33432 69328 0 A[6]
rlabel metal2 57512 69328 57512 69328 0 A[7]
rlabel metal2 36904 69328 36904 69328 0 CEN
rlabel metal2 59304 69328 59304 69328 0 CLK
rlabel metal2 85400 69328 85400 69328 0 D[0]
rlabel metal2 74984 69328 74984 69328 0 D[1]
rlabel metal2 73808 69342 73808 69342 0 D[2]
rlabel metal2 63392 69342 63392 69342 0 D[3]
rlabel metal2 25816 69328 25816 69328 0 D[4]
rlabel metal2 15512 69328 15512 69328 0 D[5]
rlabel metal2 14168 69328 14168 69328 0 D[6]
rlabel metal2 3808 69342 3808 69342 0 D[7]
rlabel metal2 46648 69328 46648 69328 0 GWEN
rlabel metal2 83888 69342 83888 69342 0 Q[0]
rlabel metal2 75712 69342 75712 69342 0 Q[1]
rlabel metal2 73080 69328 73080 69328 0 Q[2]
rlabel metal2 65016 69328 65016 69328 0 Q[3]
rlabel metal2 24304 69342 24304 69342 0 Q[4]
rlabel metal2 16072 69328 16072 69328 0 Q[5]
rlabel metal2 13496 69328 13496 69328 0 Q[6]
rlabel metal2 5432 69328 5432 69328 0 Q[7]
rlabel metal2 84728 69328 84728 69328 0 WEN[0]
rlabel metal2 74592 69342 74592 69342 0 WEN[1]
rlabel metal2 74200 69328 74200 69328 0 WEN[2]
rlabel metal2 63784 69328 63784 69328 0 WEN[3]
rlabel metal2 25088 69342 25088 69342 0 WEN[4]
rlabel metal2 15064 69328 15064 69328 0 WEN[5]
rlabel metal2 14616 69328 14616 69328 0 WEN[6]
rlabel metal2 4536 69328 4536 69328 0 WEN[7]
<< properties >>
string FIXED_BBOX 0 0 88972 70376
<< end >>
