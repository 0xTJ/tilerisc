VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO risc16
  CLASS BLOCK ;
  FOREIGN risc16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END clk
  PIN dmem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END dmem_addr[0]
  PIN dmem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 4.000 68.880 ;
    END
  END dmem_addr[10]
  PIN dmem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END dmem_addr[11]
  PIN dmem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END dmem_addr[12]
  PIN dmem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 4.000 31.920 ;
    END
  END dmem_addr[13]
  PIN dmem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 4.000 19.600 ;
    END
  END dmem_addr[14]
  PIN dmem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.720 4.000 7.280 ;
    END
  END dmem_addr[15]
  PIN dmem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END dmem_addr[1]
  PIN dmem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END dmem_addr[2]
  PIN dmem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END dmem_addr[3]
  PIN dmem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 4.000 142.800 ;
    END
  END dmem_addr[4]
  PIN dmem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END dmem_addr[5]
  PIN dmem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END dmem_addr[6]
  PIN dmem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END dmem_addr[7]
  PIN dmem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 4.000 93.520 ;
    END
  END dmem_addr[8]
  PIN dmem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END dmem_addr[9]
  PIN dmem_data_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 6.720 400.000 7.280 ;
    END
  END dmem_data_in[0]
  PIN dmem_data_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 129.920 400.000 130.480 ;
    END
  END dmem_data_in[10]
  PIN dmem_data_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 142.240 400.000 142.800 ;
    END
  END dmem_data_in[11]
  PIN dmem_data_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 154.560 400.000 155.120 ;
    END
  END dmem_data_in[12]
  PIN dmem_data_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 166.880 400.000 167.440 ;
    END
  END dmem_data_in[13]
  PIN dmem_data_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 179.200 400.000 179.760 ;
    END
  END dmem_data_in[14]
  PIN dmem_data_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 191.520 400.000 192.080 ;
    END
  END dmem_data_in[15]
  PIN dmem_data_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 19.040 400.000 19.600 ;
    END
  END dmem_data_in[1]
  PIN dmem_data_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 31.360 400.000 31.920 ;
    END
  END dmem_data_in[2]
  PIN dmem_data_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 43.680 400.000 44.240 ;
    END
  END dmem_data_in[3]
  PIN dmem_data_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 56.000 400.000 56.560 ;
    END
  END dmem_data_in[4]
  PIN dmem_data_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 68.320 400.000 68.880 ;
    END
  END dmem_data_in[5]
  PIN dmem_data_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 80.640 400.000 81.200 ;
    END
  END dmem_data_in[6]
  PIN dmem_data_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 92.960 400.000 93.520 ;
    END
  END dmem_data_in[7]
  PIN dmem_data_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 105.280 400.000 105.840 ;
    END
  END dmem_data_in[8]
  PIN dmem_data_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 117.600 400.000 118.160 ;
    END
  END dmem_data_in[9]
  PIN dmem_data_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 0.000 18.480 4.000 ;
    END
  END dmem_data_out[0]
  PIN dmem_data_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 0.000 220.080 4.000 ;
    END
  END dmem_data_out[10]
  PIN dmem_data_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END dmem_data_out[11]
  PIN dmem_data_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END dmem_data_out[12]
  PIN dmem_data_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END dmem_data_out[13]
  PIN dmem_data_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 0.000 300.720 4.000 ;
    END
  END dmem_data_out[14]
  PIN dmem_data_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END dmem_data_out[15]
  PIN dmem_data_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END dmem_data_out[1]
  PIN dmem_data_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END dmem_data_out[2]
  PIN dmem_data_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END dmem_data_out[3]
  PIN dmem_data_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END dmem_data_out[4]
  PIN dmem_data_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END dmem_data_out[5]
  PIN dmem_data_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END dmem_data_out[6]
  PIN dmem_data_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END dmem_data_out[7]
  PIN dmem_data_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END dmem_data_out[8]
  PIN dmem_data_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END dmem_data_out[9]
  PIN dmem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END dmem_we
  PIN instr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 196.000 193.200 200.000 ;
    END
  END instr[0]
  PIN instr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 196.000 70.000 200.000 ;
    END
  END instr[10]
  PIN instr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 196.000 57.680 200.000 ;
    END
  END instr[11]
  PIN instr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 196.000 45.360 200.000 ;
    END
  END instr[12]
  PIN instr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 196.000 33.040 200.000 ;
    END
  END instr[13]
  PIN instr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 196.000 20.720 200.000 ;
    END
  END instr[14]
  PIN instr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 196.000 8.400 200.000 ;
    END
  END instr[15]
  PIN instr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 196.000 180.880 200.000 ;
    END
  END instr[1]
  PIN instr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 196.000 168.560 200.000 ;
    END
  END instr[2]
  PIN instr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 196.000 156.240 200.000 ;
    END
  END instr[3]
  PIN instr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 196.000 143.920 200.000 ;
    END
  END instr[4]
  PIN instr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 196.000 131.600 200.000 ;
    END
  END instr[5]
  PIN instr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 196.000 119.280 200.000 ;
    END
  END instr[6]
  PIN instr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 196.000 106.960 200.000 ;
    END
  END instr[7]
  PIN instr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 196.000 94.640 200.000 ;
    END
  END instr[8]
  PIN instr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 196.000 82.320 200.000 ;
    END
  END instr[9]
  PIN pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 196.000 390.320 200.000 ;
    END
  END pc[0]
  PIN pc[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 196.000 267.120 200.000 ;
    END
  END pc[10]
  PIN pc[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 196.000 254.800 200.000 ;
    END
  END pc[11]
  PIN pc[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 196.000 242.480 200.000 ;
    END
  END pc[12]
  PIN pc[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 196.000 230.160 200.000 ;
    END
  END pc[13]
  PIN pc[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 196.000 217.840 200.000 ;
    END
  END pc[14]
  PIN pc[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 196.000 205.520 200.000 ;
    END
  END pc[15]
  PIN pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 196.000 378.000 200.000 ;
    END
  END pc[1]
  PIN pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 196.000 365.680 200.000 ;
    END
  END pc[2]
  PIN pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 196.000 353.360 200.000 ;
    END
  END pc[3]
  PIN pc[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 196.000 341.040 200.000 ;
    END
  END pc[4]
  PIN pc[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 196.000 328.720 200.000 ;
    END
  END pc[5]
  PIN pc[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 196.000 316.400 200.000 ;
    END
  END pc[6]
  PIN pc[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 196.000 304.080 200.000 ;
    END
  END pc[7]
  PIN pc[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 196.000 291.760 200.000 ;
    END
  END pc[8]
  PIN pc[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 196.000 279.440 200.000 ;
    END
  END pc[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 54.220 15.380 55.820 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.820 15.380 152.420 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 247.420 15.380 249.020 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 344.020 15.380 345.620 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 102.520 15.380 104.120 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 199.120 15.380 200.720 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 295.720 15.380 297.320 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.320 15.380 393.920 184.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 393.920 184.540 ;
      LAYER Metal2 ;
        RECT 8.700 195.700 19.860 196.420 ;
        RECT 21.020 195.700 32.180 196.420 ;
        RECT 33.340 195.700 44.500 196.420 ;
        RECT 45.660 195.700 56.820 196.420 ;
        RECT 57.980 195.700 69.140 196.420 ;
        RECT 70.300 195.700 81.460 196.420 ;
        RECT 82.620 195.700 93.780 196.420 ;
        RECT 94.940 195.700 106.100 196.420 ;
        RECT 107.260 195.700 118.420 196.420 ;
        RECT 119.580 195.700 130.740 196.420 ;
        RECT 131.900 195.700 143.060 196.420 ;
        RECT 144.220 195.700 155.380 196.420 ;
        RECT 156.540 195.700 167.700 196.420 ;
        RECT 168.860 195.700 180.020 196.420 ;
        RECT 181.180 195.700 192.340 196.420 ;
        RECT 193.500 195.700 204.660 196.420 ;
        RECT 205.820 195.700 216.980 196.420 ;
        RECT 218.140 195.700 229.300 196.420 ;
        RECT 230.460 195.700 241.620 196.420 ;
        RECT 242.780 195.700 253.940 196.420 ;
        RECT 255.100 195.700 266.260 196.420 ;
        RECT 267.420 195.700 278.580 196.420 ;
        RECT 279.740 195.700 290.900 196.420 ;
        RECT 292.060 195.700 303.220 196.420 ;
        RECT 304.380 195.700 315.540 196.420 ;
        RECT 316.700 195.700 327.860 196.420 ;
        RECT 329.020 195.700 340.180 196.420 ;
        RECT 341.340 195.700 352.500 196.420 ;
        RECT 353.660 195.700 364.820 196.420 ;
        RECT 365.980 195.700 377.140 196.420 ;
        RECT 378.300 195.700 389.460 196.420 ;
        RECT 390.620 195.700 393.780 196.420 ;
        RECT 7.980 4.300 393.780 195.700 ;
        RECT 7.980 3.500 17.620 4.300 ;
        RECT 18.780 3.500 37.780 4.300 ;
        RECT 38.940 3.500 57.940 4.300 ;
        RECT 59.100 3.500 78.100 4.300 ;
        RECT 79.260 3.500 98.260 4.300 ;
        RECT 99.420 3.500 118.420 4.300 ;
        RECT 119.580 3.500 138.580 4.300 ;
        RECT 139.740 3.500 158.740 4.300 ;
        RECT 159.900 3.500 178.900 4.300 ;
        RECT 180.060 3.500 199.060 4.300 ;
        RECT 200.220 3.500 219.220 4.300 ;
        RECT 220.380 3.500 239.380 4.300 ;
        RECT 240.540 3.500 259.540 4.300 ;
        RECT 260.700 3.500 279.700 4.300 ;
        RECT 280.860 3.500 299.860 4.300 ;
        RECT 301.020 3.500 320.020 4.300 ;
        RECT 321.180 3.500 340.180 4.300 ;
        RECT 341.340 3.500 360.340 4.300 ;
        RECT 361.500 3.500 380.500 4.300 ;
        RECT 381.660 3.500 393.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 191.220 395.700 191.940 ;
        RECT 4.000 180.060 396.000 191.220 ;
        RECT 4.300 178.900 395.700 180.060 ;
        RECT 4.000 167.740 396.000 178.900 ;
        RECT 4.300 166.580 395.700 167.740 ;
        RECT 4.000 155.420 396.000 166.580 ;
        RECT 4.300 154.260 395.700 155.420 ;
        RECT 4.000 143.100 396.000 154.260 ;
        RECT 4.300 141.940 395.700 143.100 ;
        RECT 4.000 130.780 396.000 141.940 ;
        RECT 4.300 129.620 395.700 130.780 ;
        RECT 4.000 118.460 396.000 129.620 ;
        RECT 4.300 117.300 395.700 118.460 ;
        RECT 4.000 106.140 396.000 117.300 ;
        RECT 4.300 104.980 395.700 106.140 ;
        RECT 4.000 93.820 396.000 104.980 ;
        RECT 4.300 92.660 395.700 93.820 ;
        RECT 4.000 81.500 396.000 92.660 ;
        RECT 4.300 80.340 395.700 81.500 ;
        RECT 4.000 69.180 396.000 80.340 ;
        RECT 4.300 68.020 395.700 69.180 ;
        RECT 4.000 56.860 396.000 68.020 ;
        RECT 4.300 55.700 395.700 56.860 ;
        RECT 4.000 44.540 396.000 55.700 ;
        RECT 4.300 43.380 395.700 44.540 ;
        RECT 4.000 32.220 396.000 43.380 ;
        RECT 4.300 31.060 395.700 32.220 ;
        RECT 4.000 19.900 396.000 31.060 ;
        RECT 4.300 18.740 395.700 19.900 ;
        RECT 4.000 7.580 396.000 18.740 ;
        RECT 4.300 6.860 395.700 7.580 ;
  END
END risc16
END LIBRARY

