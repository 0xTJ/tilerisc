VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tinyrv
  CLASS BLOCK ;
  FOREIGN tinyrv ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 0.000 6.160 4.000 ;
    END
  END clk
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 11.200 0.000 11.760 4.000 ;
    END
  END inst[0]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END inst[10]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END inst[11]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END inst[12]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END inst[13]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END inst[14]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END inst[15]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END inst[16]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END inst[17]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END inst[18]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END inst[19]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END inst[1]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END inst[20]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END inst[21]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END inst[22]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END inst[23]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END inst[24]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END inst[25]
  PIN inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 0.000 157.360 4.000 ;
    END
  END inst[26]
  PIN inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END inst[27]
  PIN inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END inst[28]
  PIN inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END inst[29]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 0.000 22.960 4.000 ;
    END
  END inst[2]
  PIN inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END inst[30]
  PIN inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END inst[31]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 4.000 ;
    END
  END inst[3]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END inst[4]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 4.000 ;
    END
  END inst[5]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END inst[6]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END inst[7]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END inst[8]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END inst[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 596.000 510.160 600.000 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 596.000 465.360 600.000 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 596.000 460.880 600.000 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 596.000 456.400 600.000 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 596.000 451.920 600.000 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 596.000 447.440 600.000 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 596.000 442.960 600.000 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 596.000 438.480 600.000 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 596.000 434.000 600.000 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 596.000 429.520 600.000 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 596.000 425.040 600.000 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 596.000 505.680 600.000 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 596.000 420.560 600.000 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 596.000 416.080 600.000 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 596.000 411.600 600.000 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 596.000 407.120 600.000 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 596.000 402.640 600.000 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 596.000 398.160 600.000 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 596.000 393.680 600.000 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 596.000 389.200 600.000 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 596.000 384.720 600.000 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 596.000 380.240 600.000 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 596.000 501.200 600.000 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 596.000 375.760 600.000 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 596.000 371.280 600.000 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 596.000 496.720 600.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 596.000 492.240 600.000 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 596.000 487.760 600.000 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 482.720 596.000 483.280 600.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 596.000 478.800 600.000 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 596.000 474.320 600.000 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 596.000 469.840 600.000 ;
    END
  END mem_addr[9]
  PIN mem_ld_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 596.000 344.400 600.000 ;
    END
  END mem_ld_dat[0]
  PIN mem_ld_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 596.000 299.600 600.000 ;
    END
  END mem_ld_dat[10]
  PIN mem_ld_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 596.000 295.120 600.000 ;
    END
  END mem_ld_dat[11]
  PIN mem_ld_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 596.000 290.640 600.000 ;
    END
  END mem_ld_dat[12]
  PIN mem_ld_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 596.000 286.160 600.000 ;
    END
  END mem_ld_dat[13]
  PIN mem_ld_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 596.000 281.680 600.000 ;
    END
  END mem_ld_dat[14]
  PIN mem_ld_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 596.000 277.200 600.000 ;
    END
  END mem_ld_dat[15]
  PIN mem_ld_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 596.000 272.720 600.000 ;
    END
  END mem_ld_dat[16]
  PIN mem_ld_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 596.000 268.240 600.000 ;
    END
  END mem_ld_dat[17]
  PIN mem_ld_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 596.000 263.760 600.000 ;
    END
  END mem_ld_dat[18]
  PIN mem_ld_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 596.000 259.280 600.000 ;
    END
  END mem_ld_dat[19]
  PIN mem_ld_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 596.000 339.920 600.000 ;
    END
  END mem_ld_dat[1]
  PIN mem_ld_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 596.000 254.800 600.000 ;
    END
  END mem_ld_dat[20]
  PIN mem_ld_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 596.000 250.320 600.000 ;
    END
  END mem_ld_dat[21]
  PIN mem_ld_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 596.000 245.840 600.000 ;
    END
  END mem_ld_dat[22]
  PIN mem_ld_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 596.000 241.360 600.000 ;
    END
  END mem_ld_dat[23]
  PIN mem_ld_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 596.000 236.880 600.000 ;
    END
  END mem_ld_dat[24]
  PIN mem_ld_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 596.000 232.400 600.000 ;
    END
  END mem_ld_dat[25]
  PIN mem_ld_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 596.000 227.920 600.000 ;
    END
  END mem_ld_dat[26]
  PIN mem_ld_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 596.000 223.440 600.000 ;
    END
  END mem_ld_dat[27]
  PIN mem_ld_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 596.000 218.960 600.000 ;
    END
  END mem_ld_dat[28]
  PIN mem_ld_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 596.000 214.480 600.000 ;
    END
  END mem_ld_dat[29]
  PIN mem_ld_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 596.000 335.440 600.000 ;
    END
  END mem_ld_dat[2]
  PIN mem_ld_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 596.000 210.000 600.000 ;
    END
  END mem_ld_dat[30]
  PIN mem_ld_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 596.000 205.520 600.000 ;
    END
  END mem_ld_dat[31]
  PIN mem_ld_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 596.000 330.960 600.000 ;
    END
  END mem_ld_dat[3]
  PIN mem_ld_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 596.000 326.480 600.000 ;
    END
  END mem_ld_dat[4]
  PIN mem_ld_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 596.000 322.000 600.000 ;
    END
  END mem_ld_dat[5]
  PIN mem_ld_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 596.000 317.520 600.000 ;
    END
  END mem_ld_dat[6]
  PIN mem_ld_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 596.000 313.040 600.000 ;
    END
  END mem_ld_dat[7]
  PIN mem_ld_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 596.000 308.560 600.000 ;
    END
  END mem_ld_dat[8]
  PIN mem_ld_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 596.000 304.080 600.000 ;
    END
  END mem_ld_dat[9]
  PIN mem_ld_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 596.000 366.800 600.000 ;
    END
  END mem_ld_en
  PIN mem_ld_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 596.000 362.320 600.000 ;
    END
  END mem_ld_mask[0]
  PIN mem_ld_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 596.000 357.840 600.000 ;
    END
  END mem_ld_mask[1]
  PIN mem_ld_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 596.000 353.360 600.000 ;
    END
  END mem_ld_mask[2]
  PIN mem_ld_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 596.000 348.880 600.000 ;
    END
  END mem_ld_mask[3]
  PIN mem_st_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 596.000 178.640 600.000 ;
    END
  END mem_st_dat[0]
  PIN mem_st_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 596.000 133.840 600.000 ;
    END
  END mem_st_dat[10]
  PIN mem_st_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 596.000 129.360 600.000 ;
    END
  END mem_st_dat[11]
  PIN mem_st_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 596.000 124.880 600.000 ;
    END
  END mem_st_dat[12]
  PIN mem_st_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 596.000 120.400 600.000 ;
    END
  END mem_st_dat[13]
  PIN mem_st_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 596.000 115.920 600.000 ;
    END
  END mem_st_dat[14]
  PIN mem_st_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 596.000 111.440 600.000 ;
    END
  END mem_st_dat[15]
  PIN mem_st_dat[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 596.000 106.960 600.000 ;
    END
  END mem_st_dat[16]
  PIN mem_st_dat[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 596.000 102.480 600.000 ;
    END
  END mem_st_dat[17]
  PIN mem_st_dat[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 596.000 98.000 600.000 ;
    END
  END mem_st_dat[18]
  PIN mem_st_dat[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 596.000 93.520 600.000 ;
    END
  END mem_st_dat[19]
  PIN mem_st_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 596.000 174.160 600.000 ;
    END
  END mem_st_dat[1]
  PIN mem_st_dat[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 596.000 89.040 600.000 ;
    END
  END mem_st_dat[20]
  PIN mem_st_dat[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 596.000 84.560 600.000 ;
    END
  END mem_st_dat[21]
  PIN mem_st_dat[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 596.000 80.080 600.000 ;
    END
  END mem_st_dat[22]
  PIN mem_st_dat[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 596.000 75.600 600.000 ;
    END
  END mem_st_dat[23]
  PIN mem_st_dat[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 596.000 71.120 600.000 ;
    END
  END mem_st_dat[24]
  PIN mem_st_dat[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 596.000 66.640 600.000 ;
    END
  END mem_st_dat[25]
  PIN mem_st_dat[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 596.000 62.160 600.000 ;
    END
  END mem_st_dat[26]
  PIN mem_st_dat[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 596.000 57.680 600.000 ;
    END
  END mem_st_dat[27]
  PIN mem_st_dat[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 596.000 53.200 600.000 ;
    END
  END mem_st_dat[28]
  PIN mem_st_dat[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 596.000 48.720 600.000 ;
    END
  END mem_st_dat[29]
  PIN mem_st_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 596.000 169.680 600.000 ;
    END
  END mem_st_dat[2]
  PIN mem_st_dat[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 596.000 44.240 600.000 ;
    END
  END mem_st_dat[30]
  PIN mem_st_dat[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 596.000 39.760 600.000 ;
    END
  END mem_st_dat[31]
  PIN mem_st_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 596.000 165.200 600.000 ;
    END
  END mem_st_dat[3]
  PIN mem_st_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 596.000 160.720 600.000 ;
    END
  END mem_st_dat[4]
  PIN mem_st_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 596.000 156.240 600.000 ;
    END
  END mem_st_dat[5]
  PIN mem_st_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 596.000 151.760 600.000 ;
    END
  END mem_st_dat[6]
  PIN mem_st_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 596.000 147.280 600.000 ;
    END
  END mem_st_dat[7]
  PIN mem_st_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 596.000 142.800 600.000 ;
    END
  END mem_st_dat[8]
  PIN mem_st_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 596.000 138.320 600.000 ;
    END
  END mem_st_dat[9]
  PIN mem_st_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 596.000 201.040 600.000 ;
    END
  END mem_st_en
  PIN mem_st_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 596.000 196.560 600.000 ;
    END
  END mem_st_mask[0]
  PIN mem_st_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 596.000 192.080 600.000 ;
    END
  END mem_st_mask[1]
  PIN mem_st_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 596.000 187.600 600.000 ;
    END
  END mem_st_mask[2]
  PIN mem_st_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 596.000 183.120 600.000 ;
    END
  END mem_st_mask[3]
  PIN pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END pc[0]
  PIN pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END pc[10]
  PIN pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END pc[11]
  PIN pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END pc[12]
  PIN pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END pc[13]
  PIN pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 0.000 269.360 4.000 ;
    END
  END pc[14]
  PIN pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 4.000 ;
    END
  END pc[15]
  PIN pc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END pc[16]
  PIN pc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END pc[17]
  PIN pc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 0.000 291.760 4.000 ;
    END
  END pc[18]
  PIN pc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END pc[19]
  PIN pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END pc[1]
  PIN pc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END pc[20]
  PIN pc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END pc[21]
  PIN pc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END pc[22]
  PIN pc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 0.000 319.760 4.000 ;
    END
  END pc[23]
  PIN pc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END pc[24]
  PIN pc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END pc[25]
  PIN pc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 0.000 336.560 4.000 ;
    END
  END pc[26]
  PIN pc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 0.000 342.160 4.000 ;
    END
  END pc[27]
  PIN pc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END pc[28]
  PIN pc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END pc[29]
  PIN pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 0.000 202.160 4.000 ;
    END
  END pc[2]
  PIN pc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 358.400 0.000 358.960 4.000 ;
    END
  END pc[30]
  PIN pc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END pc[31]
  PIN pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END pc[3]
  PIN pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END pc[4]
  PIN pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END pc[5]
  PIN pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 0.000 224.560 4.000 ;
    END
  END pc[6]
  PIN pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END pc[7]
  PIN pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END pc[8]
  PIN pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 4.000 ;
    END
  END pc[9]
  PIN pc_next[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END pc_next[0]
  PIN pc_next[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 0.000 426.160 4.000 ;
    END
  END pc_next[10]
  PIN pc_next[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 0.000 431.760 4.000 ;
    END
  END pc_next[11]
  PIN pc_next[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 0.000 437.360 4.000 ;
    END
  END pc_next[12]
  PIN pc_next[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 0.000 442.960 4.000 ;
    END
  END pc_next[13]
  PIN pc_next[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 0.000 448.560 4.000 ;
    END
  END pc_next[14]
  PIN pc_next[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END pc_next[15]
  PIN pc_next[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END pc_next[16]
  PIN pc_next[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END pc_next[17]
  PIN pc_next[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 0.000 470.960 4.000 ;
    END
  END pc_next[18]
  PIN pc_next[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 0.000 476.560 4.000 ;
    END
  END pc_next[19]
  PIN pc_next[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END pc_next[1]
  PIN pc_next[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END pc_next[20]
  PIN pc_next[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 0.000 487.760 4.000 ;
    END
  END pc_next[21]
  PIN pc_next[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 492.800 0.000 493.360 4.000 ;
    END
  END pc_next[22]
  PIN pc_next[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 0.000 498.960 4.000 ;
    END
  END pc_next[23]
  PIN pc_next[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 0.000 504.560 4.000 ;
    END
  END pc_next[24]
  PIN pc_next[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END pc_next[25]
  PIN pc_next[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END pc_next[26]
  PIN pc_next[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 0.000 521.360 4.000 ;
    END
  END pc_next[27]
  PIN pc_next[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 0.000 526.960 4.000 ;
    END
  END pc_next[28]
  PIN pc_next[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END pc_next[29]
  PIN pc_next[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END pc_next[2]
  PIN pc_next[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 0.000 538.160 4.000 ;
    END
  END pc_next[30]
  PIN pc_next[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 0.000 543.760 4.000 ;
    END
  END pc_next[31]
  PIN pc_next[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END pc_next[3]
  PIN pc_next[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 4.000 ;
    END
  END pc_next[4]
  PIN pc_next[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END pc_next[5]
  PIN pc_next[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END pc_next[6]
  PIN pc_next[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END pc_next[7]
  PIN pc_next[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END pc_next[8]
  PIN pc_next[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 0.000 420.560 4.000 ;
    END
  END pc_next[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 543.200 585.610 ;
      LAYER Metal2 ;
        RECT 5.740 595.700 38.900 596.820 ;
        RECT 40.060 595.700 43.380 596.820 ;
        RECT 44.540 595.700 47.860 596.820 ;
        RECT 49.020 595.700 52.340 596.820 ;
        RECT 53.500 595.700 56.820 596.820 ;
        RECT 57.980 595.700 61.300 596.820 ;
        RECT 62.460 595.700 65.780 596.820 ;
        RECT 66.940 595.700 70.260 596.820 ;
        RECT 71.420 595.700 74.740 596.820 ;
        RECT 75.900 595.700 79.220 596.820 ;
        RECT 80.380 595.700 83.700 596.820 ;
        RECT 84.860 595.700 88.180 596.820 ;
        RECT 89.340 595.700 92.660 596.820 ;
        RECT 93.820 595.700 97.140 596.820 ;
        RECT 98.300 595.700 101.620 596.820 ;
        RECT 102.780 595.700 106.100 596.820 ;
        RECT 107.260 595.700 110.580 596.820 ;
        RECT 111.740 595.700 115.060 596.820 ;
        RECT 116.220 595.700 119.540 596.820 ;
        RECT 120.700 595.700 124.020 596.820 ;
        RECT 125.180 595.700 128.500 596.820 ;
        RECT 129.660 595.700 132.980 596.820 ;
        RECT 134.140 595.700 137.460 596.820 ;
        RECT 138.620 595.700 141.940 596.820 ;
        RECT 143.100 595.700 146.420 596.820 ;
        RECT 147.580 595.700 150.900 596.820 ;
        RECT 152.060 595.700 155.380 596.820 ;
        RECT 156.540 595.700 159.860 596.820 ;
        RECT 161.020 595.700 164.340 596.820 ;
        RECT 165.500 595.700 168.820 596.820 ;
        RECT 169.980 595.700 173.300 596.820 ;
        RECT 174.460 595.700 177.780 596.820 ;
        RECT 178.940 595.700 182.260 596.820 ;
        RECT 183.420 595.700 186.740 596.820 ;
        RECT 187.900 595.700 191.220 596.820 ;
        RECT 192.380 595.700 195.700 596.820 ;
        RECT 196.860 595.700 200.180 596.820 ;
        RECT 201.340 595.700 204.660 596.820 ;
        RECT 205.820 595.700 209.140 596.820 ;
        RECT 210.300 595.700 213.620 596.820 ;
        RECT 214.780 595.700 218.100 596.820 ;
        RECT 219.260 595.700 222.580 596.820 ;
        RECT 223.740 595.700 227.060 596.820 ;
        RECT 228.220 595.700 231.540 596.820 ;
        RECT 232.700 595.700 236.020 596.820 ;
        RECT 237.180 595.700 240.500 596.820 ;
        RECT 241.660 595.700 244.980 596.820 ;
        RECT 246.140 595.700 249.460 596.820 ;
        RECT 250.620 595.700 253.940 596.820 ;
        RECT 255.100 595.700 258.420 596.820 ;
        RECT 259.580 595.700 262.900 596.820 ;
        RECT 264.060 595.700 267.380 596.820 ;
        RECT 268.540 595.700 271.860 596.820 ;
        RECT 273.020 595.700 276.340 596.820 ;
        RECT 277.500 595.700 280.820 596.820 ;
        RECT 281.980 595.700 285.300 596.820 ;
        RECT 286.460 595.700 289.780 596.820 ;
        RECT 290.940 595.700 294.260 596.820 ;
        RECT 295.420 595.700 298.740 596.820 ;
        RECT 299.900 595.700 303.220 596.820 ;
        RECT 304.380 595.700 307.700 596.820 ;
        RECT 308.860 595.700 312.180 596.820 ;
        RECT 313.340 595.700 316.660 596.820 ;
        RECT 317.820 595.700 321.140 596.820 ;
        RECT 322.300 595.700 325.620 596.820 ;
        RECT 326.780 595.700 330.100 596.820 ;
        RECT 331.260 595.700 334.580 596.820 ;
        RECT 335.740 595.700 339.060 596.820 ;
        RECT 340.220 595.700 343.540 596.820 ;
        RECT 344.700 595.700 348.020 596.820 ;
        RECT 349.180 595.700 352.500 596.820 ;
        RECT 353.660 595.700 356.980 596.820 ;
        RECT 358.140 595.700 361.460 596.820 ;
        RECT 362.620 595.700 365.940 596.820 ;
        RECT 367.100 595.700 370.420 596.820 ;
        RECT 371.580 595.700 374.900 596.820 ;
        RECT 376.060 595.700 379.380 596.820 ;
        RECT 380.540 595.700 383.860 596.820 ;
        RECT 385.020 595.700 388.340 596.820 ;
        RECT 389.500 595.700 392.820 596.820 ;
        RECT 393.980 595.700 397.300 596.820 ;
        RECT 398.460 595.700 401.780 596.820 ;
        RECT 402.940 595.700 406.260 596.820 ;
        RECT 407.420 595.700 410.740 596.820 ;
        RECT 411.900 595.700 415.220 596.820 ;
        RECT 416.380 595.700 419.700 596.820 ;
        RECT 420.860 595.700 424.180 596.820 ;
        RECT 425.340 595.700 428.660 596.820 ;
        RECT 429.820 595.700 433.140 596.820 ;
        RECT 434.300 595.700 437.620 596.820 ;
        RECT 438.780 595.700 442.100 596.820 ;
        RECT 443.260 595.700 446.580 596.820 ;
        RECT 447.740 595.700 451.060 596.820 ;
        RECT 452.220 595.700 455.540 596.820 ;
        RECT 456.700 595.700 460.020 596.820 ;
        RECT 461.180 595.700 464.500 596.820 ;
        RECT 465.660 595.700 468.980 596.820 ;
        RECT 470.140 595.700 473.460 596.820 ;
        RECT 474.620 595.700 477.940 596.820 ;
        RECT 479.100 595.700 482.420 596.820 ;
        RECT 483.580 595.700 486.900 596.820 ;
        RECT 488.060 595.700 491.380 596.820 ;
        RECT 492.540 595.700 495.860 596.820 ;
        RECT 497.020 595.700 500.340 596.820 ;
        RECT 501.500 595.700 504.820 596.820 ;
        RECT 505.980 595.700 509.300 596.820 ;
        RECT 510.460 595.700 544.180 596.820 ;
        RECT 5.740 4.300 544.180 595.700 ;
        RECT 6.460 3.500 10.900 4.300 ;
        RECT 12.060 3.500 16.500 4.300 ;
        RECT 17.660 3.500 22.100 4.300 ;
        RECT 23.260 3.500 27.700 4.300 ;
        RECT 28.860 3.500 33.300 4.300 ;
        RECT 34.460 3.500 38.900 4.300 ;
        RECT 40.060 3.500 44.500 4.300 ;
        RECT 45.660 3.500 50.100 4.300 ;
        RECT 51.260 3.500 55.700 4.300 ;
        RECT 56.860 3.500 61.300 4.300 ;
        RECT 62.460 3.500 66.900 4.300 ;
        RECT 68.060 3.500 72.500 4.300 ;
        RECT 73.660 3.500 78.100 4.300 ;
        RECT 79.260 3.500 83.700 4.300 ;
        RECT 84.860 3.500 89.300 4.300 ;
        RECT 90.460 3.500 94.900 4.300 ;
        RECT 96.060 3.500 100.500 4.300 ;
        RECT 101.660 3.500 106.100 4.300 ;
        RECT 107.260 3.500 111.700 4.300 ;
        RECT 112.860 3.500 117.300 4.300 ;
        RECT 118.460 3.500 122.900 4.300 ;
        RECT 124.060 3.500 128.500 4.300 ;
        RECT 129.660 3.500 134.100 4.300 ;
        RECT 135.260 3.500 139.700 4.300 ;
        RECT 140.860 3.500 145.300 4.300 ;
        RECT 146.460 3.500 150.900 4.300 ;
        RECT 152.060 3.500 156.500 4.300 ;
        RECT 157.660 3.500 162.100 4.300 ;
        RECT 163.260 3.500 167.700 4.300 ;
        RECT 168.860 3.500 173.300 4.300 ;
        RECT 174.460 3.500 178.900 4.300 ;
        RECT 180.060 3.500 184.500 4.300 ;
        RECT 185.660 3.500 190.100 4.300 ;
        RECT 191.260 3.500 195.700 4.300 ;
        RECT 196.860 3.500 201.300 4.300 ;
        RECT 202.460 3.500 206.900 4.300 ;
        RECT 208.060 3.500 212.500 4.300 ;
        RECT 213.660 3.500 218.100 4.300 ;
        RECT 219.260 3.500 223.700 4.300 ;
        RECT 224.860 3.500 229.300 4.300 ;
        RECT 230.460 3.500 234.900 4.300 ;
        RECT 236.060 3.500 240.500 4.300 ;
        RECT 241.660 3.500 246.100 4.300 ;
        RECT 247.260 3.500 251.700 4.300 ;
        RECT 252.860 3.500 257.300 4.300 ;
        RECT 258.460 3.500 262.900 4.300 ;
        RECT 264.060 3.500 268.500 4.300 ;
        RECT 269.660 3.500 274.100 4.300 ;
        RECT 275.260 3.500 279.700 4.300 ;
        RECT 280.860 3.500 285.300 4.300 ;
        RECT 286.460 3.500 290.900 4.300 ;
        RECT 292.060 3.500 296.500 4.300 ;
        RECT 297.660 3.500 302.100 4.300 ;
        RECT 303.260 3.500 307.700 4.300 ;
        RECT 308.860 3.500 313.300 4.300 ;
        RECT 314.460 3.500 318.900 4.300 ;
        RECT 320.060 3.500 324.500 4.300 ;
        RECT 325.660 3.500 330.100 4.300 ;
        RECT 331.260 3.500 335.700 4.300 ;
        RECT 336.860 3.500 341.300 4.300 ;
        RECT 342.460 3.500 346.900 4.300 ;
        RECT 348.060 3.500 352.500 4.300 ;
        RECT 353.660 3.500 358.100 4.300 ;
        RECT 359.260 3.500 363.700 4.300 ;
        RECT 364.860 3.500 369.300 4.300 ;
        RECT 370.460 3.500 374.900 4.300 ;
        RECT 376.060 3.500 380.500 4.300 ;
        RECT 381.660 3.500 386.100 4.300 ;
        RECT 387.260 3.500 391.700 4.300 ;
        RECT 392.860 3.500 397.300 4.300 ;
        RECT 398.460 3.500 402.900 4.300 ;
        RECT 404.060 3.500 408.500 4.300 ;
        RECT 409.660 3.500 414.100 4.300 ;
        RECT 415.260 3.500 419.700 4.300 ;
        RECT 420.860 3.500 425.300 4.300 ;
        RECT 426.460 3.500 430.900 4.300 ;
        RECT 432.060 3.500 436.500 4.300 ;
        RECT 437.660 3.500 442.100 4.300 ;
        RECT 443.260 3.500 447.700 4.300 ;
        RECT 448.860 3.500 453.300 4.300 ;
        RECT 454.460 3.500 458.900 4.300 ;
        RECT 460.060 3.500 464.500 4.300 ;
        RECT 465.660 3.500 470.100 4.300 ;
        RECT 471.260 3.500 475.700 4.300 ;
        RECT 476.860 3.500 481.300 4.300 ;
        RECT 482.460 3.500 486.900 4.300 ;
        RECT 488.060 3.500 492.500 4.300 ;
        RECT 493.660 3.500 498.100 4.300 ;
        RECT 499.260 3.500 503.700 4.300 ;
        RECT 504.860 3.500 509.300 4.300 ;
        RECT 510.460 3.500 514.900 4.300 ;
        RECT 516.060 3.500 520.500 4.300 ;
        RECT 521.660 3.500 526.100 4.300 ;
        RECT 527.260 3.500 531.700 4.300 ;
        RECT 532.860 3.500 537.300 4.300 ;
        RECT 538.460 3.500 542.900 4.300 ;
        RECT 544.060 3.500 544.180 4.300 ;
      LAYER Metal3 ;
        RECT 5.690 6.860 544.230 588.980 ;
      LAYER Metal4 ;
        RECT 46.620 584.680 541.940 588.470 ;
        RECT 46.620 15.080 98.740 584.680 ;
        RECT 100.940 15.080 175.540 584.680 ;
        RECT 177.740 15.080 252.340 584.680 ;
        RECT 254.540 15.080 329.140 584.680 ;
        RECT 331.340 15.080 405.940 584.680 ;
        RECT 408.140 15.080 482.740 584.680 ;
        RECT 484.940 15.080 541.940 584.680 ;
        RECT 46.620 6.810 541.940 15.080 ;
  END
END tinyrv
END LIBRARY

