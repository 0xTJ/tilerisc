// This is the unpowered netlist.
module tinyrv (clk,
    alu_out_out,
    inst_in,
    mem_load_out);
 input clk;
 output [31:0] alu_out_out;
 input [31:0] inst_in;
 input [31:0] mem_load_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \pc[0] ;
 wire \pc[10] ;
 wire \pc[11] ;
 wire \pc[12] ;
 wire \pc[13] ;
 wire \pc[14] ;
 wire \pc[15] ;
 wire \pc[16] ;
 wire \pc[17] ;
 wire \pc[18] ;
 wire \pc[19] ;
 wire \pc[1] ;
 wire \pc[20] ;
 wire \pc[21] ;
 wire \pc[22] ;
 wire \pc[23] ;
 wire \pc[24] ;
 wire \pc[25] ;
 wire \pc[26] ;
 wire \pc[27] ;
 wire \pc[28] ;
 wire \pc[29] ;
 wire \pc[2] ;
 wire \pc[30] ;
 wire \pc[31] ;
 wire \pc[3] ;
 wire \pc[4] ;
 wire \pc[5] ;
 wire \pc[6] ;
 wire \pc[7] ;
 wire \pc[8] ;
 wire \pc[9] ;
 wire \pc_next[10] ;
 wire \pc_next[11] ;
 wire \pc_next[12] ;
 wire \pc_next[13] ;
 wire \pc_next[14] ;
 wire \pc_next[15] ;
 wire \pc_next[16] ;
 wire \pc_next[17] ;
 wire \pc_next[18] ;
 wire \pc_next[19] ;
 wire \pc_next[20] ;
 wire \pc_next[21] ;
 wire \pc_next[22] ;
 wire \pc_next[23] ;
 wire \pc_next[24] ;
 wire \pc_next[25] ;
 wire \pc_next[26] ;
 wire \pc_next[27] ;
 wire \pc_next[28] ;
 wire \pc_next[29] ;
 wire \pc_next[2] ;
 wire \pc_next[30] ;
 wire \pc_next[31] ;
 wire \pc_next[3] ;
 wire \pc_next[4] ;
 wire \pc_next[5] ;
 wire \pc_next[6] ;
 wire \pc_next[7] ;
 wire \pc_next[8] ;
 wire \pc_next[9] ;
 wire \reg_file.reg_storage[10][0] ;
 wire \reg_file.reg_storage[10][10] ;
 wire \reg_file.reg_storage[10][11] ;
 wire \reg_file.reg_storage[10][12] ;
 wire \reg_file.reg_storage[10][13] ;
 wire \reg_file.reg_storage[10][14] ;
 wire \reg_file.reg_storage[10][15] ;
 wire \reg_file.reg_storage[10][16] ;
 wire \reg_file.reg_storage[10][17] ;
 wire \reg_file.reg_storage[10][18] ;
 wire \reg_file.reg_storage[10][19] ;
 wire \reg_file.reg_storage[10][1] ;
 wire \reg_file.reg_storage[10][20] ;
 wire \reg_file.reg_storage[10][21] ;
 wire \reg_file.reg_storage[10][22] ;
 wire \reg_file.reg_storage[10][23] ;
 wire \reg_file.reg_storage[10][24] ;
 wire \reg_file.reg_storage[10][25] ;
 wire \reg_file.reg_storage[10][26] ;
 wire \reg_file.reg_storage[10][27] ;
 wire \reg_file.reg_storage[10][28] ;
 wire \reg_file.reg_storage[10][29] ;
 wire \reg_file.reg_storage[10][2] ;
 wire \reg_file.reg_storage[10][30] ;
 wire \reg_file.reg_storage[10][31] ;
 wire \reg_file.reg_storage[10][3] ;
 wire \reg_file.reg_storage[10][4] ;
 wire \reg_file.reg_storage[10][5] ;
 wire \reg_file.reg_storage[10][6] ;
 wire \reg_file.reg_storage[10][7] ;
 wire \reg_file.reg_storage[10][8] ;
 wire \reg_file.reg_storage[10][9] ;
 wire \reg_file.reg_storage[11][0] ;
 wire \reg_file.reg_storage[11][10] ;
 wire \reg_file.reg_storage[11][11] ;
 wire \reg_file.reg_storage[11][12] ;
 wire \reg_file.reg_storage[11][13] ;
 wire \reg_file.reg_storage[11][14] ;
 wire \reg_file.reg_storage[11][15] ;
 wire \reg_file.reg_storage[11][16] ;
 wire \reg_file.reg_storage[11][17] ;
 wire \reg_file.reg_storage[11][18] ;
 wire \reg_file.reg_storage[11][19] ;
 wire \reg_file.reg_storage[11][1] ;
 wire \reg_file.reg_storage[11][20] ;
 wire \reg_file.reg_storage[11][21] ;
 wire \reg_file.reg_storage[11][22] ;
 wire \reg_file.reg_storage[11][23] ;
 wire \reg_file.reg_storage[11][24] ;
 wire \reg_file.reg_storage[11][25] ;
 wire \reg_file.reg_storage[11][26] ;
 wire \reg_file.reg_storage[11][27] ;
 wire \reg_file.reg_storage[11][28] ;
 wire \reg_file.reg_storage[11][29] ;
 wire \reg_file.reg_storage[11][2] ;
 wire \reg_file.reg_storage[11][30] ;
 wire \reg_file.reg_storage[11][31] ;
 wire \reg_file.reg_storage[11][3] ;
 wire \reg_file.reg_storage[11][4] ;
 wire \reg_file.reg_storage[11][5] ;
 wire \reg_file.reg_storage[11][6] ;
 wire \reg_file.reg_storage[11][7] ;
 wire \reg_file.reg_storage[11][8] ;
 wire \reg_file.reg_storage[11][9] ;
 wire \reg_file.reg_storage[12][0] ;
 wire \reg_file.reg_storage[12][10] ;
 wire \reg_file.reg_storage[12][11] ;
 wire \reg_file.reg_storage[12][12] ;
 wire \reg_file.reg_storage[12][13] ;
 wire \reg_file.reg_storage[12][14] ;
 wire \reg_file.reg_storage[12][15] ;
 wire \reg_file.reg_storage[12][16] ;
 wire \reg_file.reg_storage[12][17] ;
 wire \reg_file.reg_storage[12][18] ;
 wire \reg_file.reg_storage[12][19] ;
 wire \reg_file.reg_storage[12][1] ;
 wire \reg_file.reg_storage[12][20] ;
 wire \reg_file.reg_storage[12][21] ;
 wire \reg_file.reg_storage[12][22] ;
 wire \reg_file.reg_storage[12][23] ;
 wire \reg_file.reg_storage[12][24] ;
 wire \reg_file.reg_storage[12][25] ;
 wire \reg_file.reg_storage[12][26] ;
 wire \reg_file.reg_storage[12][27] ;
 wire \reg_file.reg_storage[12][28] ;
 wire \reg_file.reg_storage[12][29] ;
 wire \reg_file.reg_storage[12][2] ;
 wire \reg_file.reg_storage[12][30] ;
 wire \reg_file.reg_storage[12][31] ;
 wire \reg_file.reg_storage[12][3] ;
 wire \reg_file.reg_storage[12][4] ;
 wire \reg_file.reg_storage[12][5] ;
 wire \reg_file.reg_storage[12][6] ;
 wire \reg_file.reg_storage[12][7] ;
 wire \reg_file.reg_storage[12][8] ;
 wire \reg_file.reg_storage[12][9] ;
 wire \reg_file.reg_storage[13][0] ;
 wire \reg_file.reg_storage[13][10] ;
 wire \reg_file.reg_storage[13][11] ;
 wire \reg_file.reg_storage[13][12] ;
 wire \reg_file.reg_storage[13][13] ;
 wire \reg_file.reg_storage[13][14] ;
 wire \reg_file.reg_storage[13][15] ;
 wire \reg_file.reg_storage[13][16] ;
 wire \reg_file.reg_storage[13][17] ;
 wire \reg_file.reg_storage[13][18] ;
 wire \reg_file.reg_storage[13][19] ;
 wire \reg_file.reg_storage[13][1] ;
 wire \reg_file.reg_storage[13][20] ;
 wire \reg_file.reg_storage[13][21] ;
 wire \reg_file.reg_storage[13][22] ;
 wire \reg_file.reg_storage[13][23] ;
 wire \reg_file.reg_storage[13][24] ;
 wire \reg_file.reg_storage[13][25] ;
 wire \reg_file.reg_storage[13][26] ;
 wire \reg_file.reg_storage[13][27] ;
 wire \reg_file.reg_storage[13][28] ;
 wire \reg_file.reg_storage[13][29] ;
 wire \reg_file.reg_storage[13][2] ;
 wire \reg_file.reg_storage[13][30] ;
 wire \reg_file.reg_storage[13][31] ;
 wire \reg_file.reg_storage[13][3] ;
 wire \reg_file.reg_storage[13][4] ;
 wire \reg_file.reg_storage[13][5] ;
 wire \reg_file.reg_storage[13][6] ;
 wire \reg_file.reg_storage[13][7] ;
 wire \reg_file.reg_storage[13][8] ;
 wire \reg_file.reg_storage[13][9] ;
 wire \reg_file.reg_storage[14][0] ;
 wire \reg_file.reg_storage[14][10] ;
 wire \reg_file.reg_storage[14][11] ;
 wire \reg_file.reg_storage[14][12] ;
 wire \reg_file.reg_storage[14][13] ;
 wire \reg_file.reg_storage[14][14] ;
 wire \reg_file.reg_storage[14][15] ;
 wire \reg_file.reg_storage[14][16] ;
 wire \reg_file.reg_storage[14][17] ;
 wire \reg_file.reg_storage[14][18] ;
 wire \reg_file.reg_storage[14][19] ;
 wire \reg_file.reg_storage[14][1] ;
 wire \reg_file.reg_storage[14][20] ;
 wire \reg_file.reg_storage[14][21] ;
 wire \reg_file.reg_storage[14][22] ;
 wire \reg_file.reg_storage[14][23] ;
 wire \reg_file.reg_storage[14][24] ;
 wire \reg_file.reg_storage[14][25] ;
 wire \reg_file.reg_storage[14][26] ;
 wire \reg_file.reg_storage[14][27] ;
 wire \reg_file.reg_storage[14][28] ;
 wire \reg_file.reg_storage[14][29] ;
 wire \reg_file.reg_storage[14][2] ;
 wire \reg_file.reg_storage[14][30] ;
 wire \reg_file.reg_storage[14][31] ;
 wire \reg_file.reg_storage[14][3] ;
 wire \reg_file.reg_storage[14][4] ;
 wire \reg_file.reg_storage[14][5] ;
 wire \reg_file.reg_storage[14][6] ;
 wire \reg_file.reg_storage[14][7] ;
 wire \reg_file.reg_storage[14][8] ;
 wire \reg_file.reg_storage[14][9] ;
 wire \reg_file.reg_storage[15][0] ;
 wire \reg_file.reg_storage[15][10] ;
 wire \reg_file.reg_storage[15][11] ;
 wire \reg_file.reg_storage[15][12] ;
 wire \reg_file.reg_storage[15][13] ;
 wire \reg_file.reg_storage[15][14] ;
 wire \reg_file.reg_storage[15][15] ;
 wire \reg_file.reg_storage[15][16] ;
 wire \reg_file.reg_storage[15][17] ;
 wire \reg_file.reg_storage[15][18] ;
 wire \reg_file.reg_storage[15][19] ;
 wire \reg_file.reg_storage[15][1] ;
 wire \reg_file.reg_storage[15][20] ;
 wire \reg_file.reg_storage[15][21] ;
 wire \reg_file.reg_storage[15][22] ;
 wire \reg_file.reg_storage[15][23] ;
 wire \reg_file.reg_storage[15][24] ;
 wire \reg_file.reg_storage[15][25] ;
 wire \reg_file.reg_storage[15][26] ;
 wire \reg_file.reg_storage[15][27] ;
 wire \reg_file.reg_storage[15][28] ;
 wire \reg_file.reg_storage[15][29] ;
 wire \reg_file.reg_storage[15][2] ;
 wire \reg_file.reg_storage[15][30] ;
 wire \reg_file.reg_storage[15][31] ;
 wire \reg_file.reg_storage[15][3] ;
 wire \reg_file.reg_storage[15][4] ;
 wire \reg_file.reg_storage[15][5] ;
 wire \reg_file.reg_storage[15][6] ;
 wire \reg_file.reg_storage[15][7] ;
 wire \reg_file.reg_storage[15][8] ;
 wire \reg_file.reg_storage[15][9] ;
 wire \reg_file.reg_storage[1][0] ;
 wire \reg_file.reg_storage[1][10] ;
 wire \reg_file.reg_storage[1][11] ;
 wire \reg_file.reg_storage[1][12] ;
 wire \reg_file.reg_storage[1][13] ;
 wire \reg_file.reg_storage[1][14] ;
 wire \reg_file.reg_storage[1][15] ;
 wire \reg_file.reg_storage[1][16] ;
 wire \reg_file.reg_storage[1][17] ;
 wire \reg_file.reg_storage[1][18] ;
 wire \reg_file.reg_storage[1][19] ;
 wire \reg_file.reg_storage[1][1] ;
 wire \reg_file.reg_storage[1][20] ;
 wire \reg_file.reg_storage[1][21] ;
 wire \reg_file.reg_storage[1][22] ;
 wire \reg_file.reg_storage[1][23] ;
 wire \reg_file.reg_storage[1][24] ;
 wire \reg_file.reg_storage[1][25] ;
 wire \reg_file.reg_storage[1][26] ;
 wire \reg_file.reg_storage[1][27] ;
 wire \reg_file.reg_storage[1][28] ;
 wire \reg_file.reg_storage[1][29] ;
 wire \reg_file.reg_storage[1][2] ;
 wire \reg_file.reg_storage[1][30] ;
 wire \reg_file.reg_storage[1][31] ;
 wire \reg_file.reg_storage[1][3] ;
 wire \reg_file.reg_storage[1][4] ;
 wire \reg_file.reg_storage[1][5] ;
 wire \reg_file.reg_storage[1][6] ;
 wire \reg_file.reg_storage[1][7] ;
 wire \reg_file.reg_storage[1][8] ;
 wire \reg_file.reg_storage[1][9] ;
 wire \reg_file.reg_storage[2][0] ;
 wire \reg_file.reg_storage[2][10] ;
 wire \reg_file.reg_storage[2][11] ;
 wire \reg_file.reg_storage[2][12] ;
 wire \reg_file.reg_storage[2][13] ;
 wire \reg_file.reg_storage[2][14] ;
 wire \reg_file.reg_storage[2][15] ;
 wire \reg_file.reg_storage[2][16] ;
 wire \reg_file.reg_storage[2][17] ;
 wire \reg_file.reg_storage[2][18] ;
 wire \reg_file.reg_storage[2][19] ;
 wire \reg_file.reg_storage[2][1] ;
 wire \reg_file.reg_storage[2][20] ;
 wire \reg_file.reg_storage[2][21] ;
 wire \reg_file.reg_storage[2][22] ;
 wire \reg_file.reg_storage[2][23] ;
 wire \reg_file.reg_storage[2][24] ;
 wire \reg_file.reg_storage[2][25] ;
 wire \reg_file.reg_storage[2][26] ;
 wire \reg_file.reg_storage[2][27] ;
 wire \reg_file.reg_storage[2][28] ;
 wire \reg_file.reg_storage[2][29] ;
 wire \reg_file.reg_storage[2][2] ;
 wire \reg_file.reg_storage[2][30] ;
 wire \reg_file.reg_storage[2][31] ;
 wire \reg_file.reg_storage[2][3] ;
 wire \reg_file.reg_storage[2][4] ;
 wire \reg_file.reg_storage[2][5] ;
 wire \reg_file.reg_storage[2][6] ;
 wire \reg_file.reg_storage[2][7] ;
 wire \reg_file.reg_storage[2][8] ;
 wire \reg_file.reg_storage[2][9] ;
 wire \reg_file.reg_storage[3][0] ;
 wire \reg_file.reg_storage[3][10] ;
 wire \reg_file.reg_storage[3][11] ;
 wire \reg_file.reg_storage[3][12] ;
 wire \reg_file.reg_storage[3][13] ;
 wire \reg_file.reg_storage[3][14] ;
 wire \reg_file.reg_storage[3][15] ;
 wire \reg_file.reg_storage[3][16] ;
 wire \reg_file.reg_storage[3][17] ;
 wire \reg_file.reg_storage[3][18] ;
 wire \reg_file.reg_storage[3][19] ;
 wire \reg_file.reg_storage[3][1] ;
 wire \reg_file.reg_storage[3][20] ;
 wire \reg_file.reg_storage[3][21] ;
 wire \reg_file.reg_storage[3][22] ;
 wire \reg_file.reg_storage[3][23] ;
 wire \reg_file.reg_storage[3][24] ;
 wire \reg_file.reg_storage[3][25] ;
 wire \reg_file.reg_storage[3][26] ;
 wire \reg_file.reg_storage[3][27] ;
 wire \reg_file.reg_storage[3][28] ;
 wire \reg_file.reg_storage[3][29] ;
 wire \reg_file.reg_storage[3][2] ;
 wire \reg_file.reg_storage[3][30] ;
 wire \reg_file.reg_storage[3][31] ;
 wire \reg_file.reg_storage[3][3] ;
 wire \reg_file.reg_storage[3][4] ;
 wire \reg_file.reg_storage[3][5] ;
 wire \reg_file.reg_storage[3][6] ;
 wire \reg_file.reg_storage[3][7] ;
 wire \reg_file.reg_storage[3][8] ;
 wire \reg_file.reg_storage[3][9] ;
 wire \reg_file.reg_storage[4][0] ;
 wire \reg_file.reg_storage[4][10] ;
 wire \reg_file.reg_storage[4][11] ;
 wire \reg_file.reg_storage[4][12] ;
 wire \reg_file.reg_storage[4][13] ;
 wire \reg_file.reg_storage[4][14] ;
 wire \reg_file.reg_storage[4][15] ;
 wire \reg_file.reg_storage[4][16] ;
 wire \reg_file.reg_storage[4][17] ;
 wire \reg_file.reg_storage[4][18] ;
 wire \reg_file.reg_storage[4][19] ;
 wire \reg_file.reg_storage[4][1] ;
 wire \reg_file.reg_storage[4][20] ;
 wire \reg_file.reg_storage[4][21] ;
 wire \reg_file.reg_storage[4][22] ;
 wire \reg_file.reg_storage[4][23] ;
 wire \reg_file.reg_storage[4][24] ;
 wire \reg_file.reg_storage[4][25] ;
 wire \reg_file.reg_storage[4][26] ;
 wire \reg_file.reg_storage[4][27] ;
 wire \reg_file.reg_storage[4][28] ;
 wire \reg_file.reg_storage[4][29] ;
 wire \reg_file.reg_storage[4][2] ;
 wire \reg_file.reg_storage[4][30] ;
 wire \reg_file.reg_storage[4][31] ;
 wire \reg_file.reg_storage[4][3] ;
 wire \reg_file.reg_storage[4][4] ;
 wire \reg_file.reg_storage[4][5] ;
 wire \reg_file.reg_storage[4][6] ;
 wire \reg_file.reg_storage[4][7] ;
 wire \reg_file.reg_storage[4][8] ;
 wire \reg_file.reg_storage[4][9] ;
 wire \reg_file.reg_storage[5][0] ;
 wire \reg_file.reg_storage[5][10] ;
 wire \reg_file.reg_storage[5][11] ;
 wire \reg_file.reg_storage[5][12] ;
 wire \reg_file.reg_storage[5][13] ;
 wire \reg_file.reg_storage[5][14] ;
 wire \reg_file.reg_storage[5][15] ;
 wire \reg_file.reg_storage[5][16] ;
 wire \reg_file.reg_storage[5][17] ;
 wire \reg_file.reg_storage[5][18] ;
 wire \reg_file.reg_storage[5][19] ;
 wire \reg_file.reg_storage[5][1] ;
 wire \reg_file.reg_storage[5][20] ;
 wire \reg_file.reg_storage[5][21] ;
 wire \reg_file.reg_storage[5][22] ;
 wire \reg_file.reg_storage[5][23] ;
 wire \reg_file.reg_storage[5][24] ;
 wire \reg_file.reg_storage[5][25] ;
 wire \reg_file.reg_storage[5][26] ;
 wire \reg_file.reg_storage[5][27] ;
 wire \reg_file.reg_storage[5][28] ;
 wire \reg_file.reg_storage[5][29] ;
 wire \reg_file.reg_storage[5][2] ;
 wire \reg_file.reg_storage[5][30] ;
 wire \reg_file.reg_storage[5][31] ;
 wire \reg_file.reg_storage[5][3] ;
 wire \reg_file.reg_storage[5][4] ;
 wire \reg_file.reg_storage[5][5] ;
 wire \reg_file.reg_storage[5][6] ;
 wire \reg_file.reg_storage[5][7] ;
 wire \reg_file.reg_storage[5][8] ;
 wire \reg_file.reg_storage[5][9] ;
 wire \reg_file.reg_storage[6][0] ;
 wire \reg_file.reg_storage[6][10] ;
 wire \reg_file.reg_storage[6][11] ;
 wire \reg_file.reg_storage[6][12] ;
 wire \reg_file.reg_storage[6][13] ;
 wire \reg_file.reg_storage[6][14] ;
 wire \reg_file.reg_storage[6][15] ;
 wire \reg_file.reg_storage[6][16] ;
 wire \reg_file.reg_storage[6][17] ;
 wire \reg_file.reg_storage[6][18] ;
 wire \reg_file.reg_storage[6][19] ;
 wire \reg_file.reg_storage[6][1] ;
 wire \reg_file.reg_storage[6][20] ;
 wire \reg_file.reg_storage[6][21] ;
 wire \reg_file.reg_storage[6][22] ;
 wire \reg_file.reg_storage[6][23] ;
 wire \reg_file.reg_storage[6][24] ;
 wire \reg_file.reg_storage[6][25] ;
 wire \reg_file.reg_storage[6][26] ;
 wire \reg_file.reg_storage[6][27] ;
 wire \reg_file.reg_storage[6][28] ;
 wire \reg_file.reg_storage[6][29] ;
 wire \reg_file.reg_storage[6][2] ;
 wire \reg_file.reg_storage[6][30] ;
 wire \reg_file.reg_storage[6][31] ;
 wire \reg_file.reg_storage[6][3] ;
 wire \reg_file.reg_storage[6][4] ;
 wire \reg_file.reg_storage[6][5] ;
 wire \reg_file.reg_storage[6][6] ;
 wire \reg_file.reg_storage[6][7] ;
 wire \reg_file.reg_storage[6][8] ;
 wire \reg_file.reg_storage[6][9] ;
 wire \reg_file.reg_storage[7][0] ;
 wire \reg_file.reg_storage[7][10] ;
 wire \reg_file.reg_storage[7][11] ;
 wire \reg_file.reg_storage[7][12] ;
 wire \reg_file.reg_storage[7][13] ;
 wire \reg_file.reg_storage[7][14] ;
 wire \reg_file.reg_storage[7][15] ;
 wire \reg_file.reg_storage[7][16] ;
 wire \reg_file.reg_storage[7][17] ;
 wire \reg_file.reg_storage[7][18] ;
 wire \reg_file.reg_storage[7][19] ;
 wire \reg_file.reg_storage[7][1] ;
 wire \reg_file.reg_storage[7][20] ;
 wire \reg_file.reg_storage[7][21] ;
 wire \reg_file.reg_storage[7][22] ;
 wire \reg_file.reg_storage[7][23] ;
 wire \reg_file.reg_storage[7][24] ;
 wire \reg_file.reg_storage[7][25] ;
 wire \reg_file.reg_storage[7][26] ;
 wire \reg_file.reg_storage[7][27] ;
 wire \reg_file.reg_storage[7][28] ;
 wire \reg_file.reg_storage[7][29] ;
 wire \reg_file.reg_storage[7][2] ;
 wire \reg_file.reg_storage[7][30] ;
 wire \reg_file.reg_storage[7][31] ;
 wire \reg_file.reg_storage[7][3] ;
 wire \reg_file.reg_storage[7][4] ;
 wire \reg_file.reg_storage[7][5] ;
 wire \reg_file.reg_storage[7][6] ;
 wire \reg_file.reg_storage[7][7] ;
 wire \reg_file.reg_storage[7][8] ;
 wire \reg_file.reg_storage[7][9] ;
 wire \reg_file.reg_storage[8][0] ;
 wire \reg_file.reg_storage[8][10] ;
 wire \reg_file.reg_storage[8][11] ;
 wire \reg_file.reg_storage[8][12] ;
 wire \reg_file.reg_storage[8][13] ;
 wire \reg_file.reg_storage[8][14] ;
 wire \reg_file.reg_storage[8][15] ;
 wire \reg_file.reg_storage[8][16] ;
 wire \reg_file.reg_storage[8][17] ;
 wire \reg_file.reg_storage[8][18] ;
 wire \reg_file.reg_storage[8][19] ;
 wire \reg_file.reg_storage[8][1] ;
 wire \reg_file.reg_storage[8][20] ;
 wire \reg_file.reg_storage[8][21] ;
 wire \reg_file.reg_storage[8][22] ;
 wire \reg_file.reg_storage[8][23] ;
 wire \reg_file.reg_storage[8][24] ;
 wire \reg_file.reg_storage[8][25] ;
 wire \reg_file.reg_storage[8][26] ;
 wire \reg_file.reg_storage[8][27] ;
 wire \reg_file.reg_storage[8][28] ;
 wire \reg_file.reg_storage[8][29] ;
 wire \reg_file.reg_storage[8][2] ;
 wire \reg_file.reg_storage[8][30] ;
 wire \reg_file.reg_storage[8][31] ;
 wire \reg_file.reg_storage[8][3] ;
 wire \reg_file.reg_storage[8][4] ;
 wire \reg_file.reg_storage[8][5] ;
 wire \reg_file.reg_storage[8][6] ;
 wire \reg_file.reg_storage[8][7] ;
 wire \reg_file.reg_storage[8][8] ;
 wire \reg_file.reg_storage[8][9] ;
 wire \reg_file.reg_storage[9][0] ;
 wire \reg_file.reg_storage[9][10] ;
 wire \reg_file.reg_storage[9][11] ;
 wire \reg_file.reg_storage[9][12] ;
 wire \reg_file.reg_storage[9][13] ;
 wire \reg_file.reg_storage[9][14] ;
 wire \reg_file.reg_storage[9][15] ;
 wire \reg_file.reg_storage[9][16] ;
 wire \reg_file.reg_storage[9][17] ;
 wire \reg_file.reg_storage[9][18] ;
 wire \reg_file.reg_storage[9][19] ;
 wire \reg_file.reg_storage[9][1] ;
 wire \reg_file.reg_storage[9][20] ;
 wire \reg_file.reg_storage[9][21] ;
 wire \reg_file.reg_storage[9][22] ;
 wire \reg_file.reg_storage[9][23] ;
 wire \reg_file.reg_storage[9][24] ;
 wire \reg_file.reg_storage[9][25] ;
 wire \reg_file.reg_storage[9][26] ;
 wire \reg_file.reg_storage[9][27] ;
 wire \reg_file.reg_storage[9][28] ;
 wire \reg_file.reg_storage[9][29] ;
 wire \reg_file.reg_storage[9][2] ;
 wire \reg_file.reg_storage[9][30] ;
 wire \reg_file.reg_storage[9][31] ;
 wire \reg_file.reg_storage[9][3] ;
 wire \reg_file.reg_storage[9][4] ;
 wire \reg_file.reg_storage[9][5] ;
 wire \reg_file.reg_storage[9][6] ;
 wire \reg_file.reg_storage[9][7] ;
 wire \reg_file.reg_storage[9][8] ;
 wire \reg_file.reg_storage[9][9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__B2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A3 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__S0 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__S1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__S (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__S (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__S0 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__S1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__S0 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__S1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__S0 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__S1 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A3 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A3 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__I (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__S1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__S (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__S0 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__S1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(\pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__B2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__S (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I3 (.I(\reg_file.reg_storage[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__S0 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__S1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__S0 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__S1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__S0 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__S1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__S (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I3 (.I(\reg_file.reg_storage[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__S0 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__S0 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__S1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__S0 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__S1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__S0 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__S1 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A3 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__B (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A3 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__S1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__S (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__S (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__S1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__S1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__S0 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__S1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__B1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__B2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__S0 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__S1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__S (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__S (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__S0 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__S1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__S0 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__S1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__S0 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__S1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A3 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A3 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__I (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I3 (.I(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__S0 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__S1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__B (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__S0 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__S1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__S0 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__S1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I0 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I3 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__S0 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__S1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(\pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__I (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__I (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__S0 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__S1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__I (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__B (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__S0 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__S1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__I0 (.I(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__S0 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__S1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__S0 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__S1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__B1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__B2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__S0 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__S1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__I (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(\reg_file.reg_storage[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__B (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__S0 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__S1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S0 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I0 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I3 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__S0 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__S1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__B1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__B2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__I (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I2 (.I(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I3 (.I(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__S0 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__S1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(\reg_file.reg_storage[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__I1 (.I(\reg_file.reg_storage[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__I2 (.I(\reg_file.reg_storage[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__S0 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__S1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__S0 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__S1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I3 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__S0 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__S1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__B1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__B2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__S0 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__S1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__I (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__B (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__S0 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__S1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__S0 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__S1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__S0 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__S1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__B1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__B2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__S0 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__S1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__B (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__I (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__S0 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__S1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__S0 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__S1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__B (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__S0 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__S1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__S0 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__S1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__S0 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__S1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__B1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__B2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__C (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__S0 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__S1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__C (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__B (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__B (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__S1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__S0 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__S1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__B (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A3 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__B2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__C (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I0 (.I(\reg_file.reg_storage[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__S0 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__S1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__S0 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__S1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__S0 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__S1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__S0 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__S1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(\pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__B2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I0 (.I(\reg_file.reg_storage[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__S0 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__S1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__B (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__S0 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__S1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__S0 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__S1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__I1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__S0 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__S1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__I (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__I (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__I3 (.I(\reg_file.reg_storage[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__S0 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__S1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__B (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__S0 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__S1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__I3 (.I(\reg_file.reg_storage[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__S0 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__S1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__I1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__S0 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__S1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__B2 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I1 (.I(\reg_file.reg_storage[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I2 (.I(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I3 (.I(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__S0 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__S1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__B (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I0 (.I(\reg_file.reg_storage[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I2 (.I(\reg_file.reg_storage[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I3 (.I(\reg_file.reg_storage[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__S0 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__S1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I0 (.I(\reg_file.reg_storage[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I1 (.I(\reg_file.reg_storage[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I2 (.I(\reg_file.reg_storage[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I3 (.I(\reg_file.reg_storage[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__S0 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__S1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__S0 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(\pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__B1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__B2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__S1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__S1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__S1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__I3 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__S0 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__S1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(\pc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__B2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__I (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__S0 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__S1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__B (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__S0 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__S1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__S0 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__S1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__S0 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__S1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__B1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__B2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__I3 (.I(\reg_file.reg_storage[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__S0 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__S1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__B (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__S0 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__S1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__S0 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__S1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__I1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__S0 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__S1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(\pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__B1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__I0 (.I(\reg_file.reg_storage[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__S0 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__S1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(\reg_file.reg_storage[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__B (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__S0 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__S1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__I0 (.I(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__S0 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__S1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__S0 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__S1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__B (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I0 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__S1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__S (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__S0 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__S1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__S0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__S1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__S0 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__S1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__B2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__I2 (.I(\reg_file.reg_storage[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__S0 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__S1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__I (.I(\reg_file.reg_storage[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__I (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__B (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__S0 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__S1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__S0 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__S1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I0 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I3 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__S0 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__S1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(\pc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__B2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__I (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I1 (.I(\reg_file.reg_storage[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I2 (.I(\reg_file.reg_storage[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I3 (.I(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__S0 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__S1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(\reg_file.reg_storage[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__B (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I1 (.I(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I2 (.I(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__S0 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__S1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I2 (.I(\reg_file.reg_storage[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I3 (.I(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__S0 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__S1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__S0 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__S1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(\pc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__B1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__B2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__S0 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__S1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__S0 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__S1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__S (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__C (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(\reg_file.reg_storage[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__B (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__S (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(\reg_file.reg_storage[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__C (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__C (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I3 (.I(\reg_file.reg_storage[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__S0 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__S1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__S0 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__S1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__I3 (.I(\reg_file.reg_storage[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__S0 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__S1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__S0 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__S1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__I3 (.I(\reg_file.reg_storage[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__S0 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__S0 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__S1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__S0 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__S0 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I3 (.I(\reg_file.reg_storage[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__S0 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__S1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__B (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__S0 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__S1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__S0 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__S1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I3 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__S0 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__S0 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__S1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A2 (.I(\reg_file.reg_storage[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__B (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__S0 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__S1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__I1 (.I(\reg_file.reg_storage[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__I2 (.I(\reg_file.reg_storage[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__S0 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__S1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__S0 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__B1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__B2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__S0 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__S1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__B (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__S0 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__S1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__S0 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__S1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__S0 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__S1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__B2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__I1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__S (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I3 (.I(\reg_file.reg_storage[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__S0 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__S1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__B (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__S0 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__S1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__S0 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__S1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I3 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__S0 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__S1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(\pc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__B2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(\pc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__S0 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__S1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__S0 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__S1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__S (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I2 (.I(\reg_file.reg_storage[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I3 (.I(\reg_file.reg_storage[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__S0 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__S1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__B (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__B (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__C (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I2 (.I(\reg_file.reg_storage[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__S0 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__S1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I (.I(\reg_file.reg_storage[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I1 (.I(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I2 (.I(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__S0 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__S1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__S0 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__S1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__S0 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__S1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__B1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__B2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I2 (.I(\reg_file.reg_storage[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__S0 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__S1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__I (.I(\reg_file.reg_storage[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__B (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I1 (.I(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__S0 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__S1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__S0 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__S1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__S0 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(\pc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__B1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__B2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I2 (.I(\reg_file.reg_storage[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I3 (.I(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__S1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__B (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I1 (.I(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I2 (.I(\reg_file.reg_storage[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__S0 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__S1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I2 (.I(\reg_file.reg_storage[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__S0 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__S1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__I3 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__S0 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__S1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(\pc[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__B1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I2 (.I(\reg_file.reg_storage[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I3 (.I(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__S0 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__S1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__B (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I1 (.I(\reg_file.reg_storage[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I2 (.I(\reg_file.reg_storage[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__S0 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__S1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__I1 (.I(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__I2 (.I(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__S0 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__S1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__S0 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__S1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__B1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__B1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__C (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A3 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__I (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__B1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__B2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A3 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__S (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__S (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__I (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__B2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__S (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__S (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__S (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__I (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__C (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__C (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__B (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__B (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__S (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__B2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__S (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__S (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__S (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__B (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__I0 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__S (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__I (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__S (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__C (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__C (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__S0 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__S1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__S (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I0 (.I(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__S (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__S0 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__S1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S0 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__S0 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__S1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__B1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__B (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__S (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__S (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__S (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I0 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__S (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__S (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__I1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__S (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__S (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__I0 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__S (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__B (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__C (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__C (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__S (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__I (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__B (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__B2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__C (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__S (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A2 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__B (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I2 (.I(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I3 (.I(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__S0 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__S1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I0 (.I(\reg_file.reg_storage[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__S (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__I1 (.I(\reg_file.reg_storage[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__I2 (.I(\reg_file.reg_storage[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__S0 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__S1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__S0 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__S1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__S0 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__S1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__B1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__B (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__S (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__B (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__C (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__B2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__S0 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__S1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__I0 (.I(\reg_file.reg_storage[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__S (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__S0 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__S1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__S0 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__S1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__S0 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__S1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__B1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__B (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__B (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__I (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__S (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__C (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__C (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__B (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__S (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__S (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__S0 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__S1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__S (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__S (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__S0 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__S1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I0 (.I(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__S0 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__S1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__S0 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__S1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__I (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__S (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I0 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__S (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I0 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__B2 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__S (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__I0 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__I1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__C (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__I1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__I3 (.I(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__S0 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__S1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__S (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__S (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__S0 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__S1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__S0 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__S1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__S0 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__S1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__B (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__B (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__B2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__S (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__I0 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__S (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__B1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__B2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I1 (.I(\reg_file.reg_storage[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I2 (.I(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I3 (.I(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__S0 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__S1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__S (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__S (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I0 (.I(\reg_file.reg_storage[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I2 (.I(\reg_file.reg_storage[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I3 (.I(\reg_file.reg_storage[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__S0 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__S1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I0 (.I(\reg_file.reg_storage[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I1 (.I(\reg_file.reg_storage[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I2 (.I(\reg_file.reg_storage[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I3 (.I(\reg_file.reg_storage[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__S0 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__S1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__S0 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__S1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__B (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__S (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__B2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__B1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__B2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__I (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__B2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__C2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__I3 (.I(\reg_file.reg_storage[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__S0 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__S1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__S (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__S (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__S0 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__S1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__I3 (.I(\reg_file.reg_storage[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__S0 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__S1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__S0 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__S1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__I (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__I (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A3 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A3 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__S (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__S (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__I (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__I (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__B (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__I1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__B (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__S (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__I (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I0 (.I(\reg_file.reg_storage[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__S0 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__S1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__I (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__S0 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__S1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__S0 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__S1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__I (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__I1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__B (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__B2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A3 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__I (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__I0 (.I(\reg_file.reg_storage[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__S0 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__S1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__I (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__S0 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__S1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__S0 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__S1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I0 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__S (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__B (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__B1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__B2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__B1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__B2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__I3 (.I(\reg_file.reg_storage[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__S0 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__S1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__S0 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__S1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__S0 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__S1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__I1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__B (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__B2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__B (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__S (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__I0 (.I(\reg_file.reg_storage[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__S0 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__S1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A2 (.I(\reg_file.reg_storage[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__S0 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__S1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__I0 (.I(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__S0 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__S1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__S1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__B2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I0 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__B2 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__B1 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__B2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__S0 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__S1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__S0 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__S1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__S0 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__S1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A3 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A4 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__B (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__S (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I0 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__B2 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__I (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__B (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__B2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__I (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__S0 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__B (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__S1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__S0 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__S0 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__S1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__B (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__I0 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__I0 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__S (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A2 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__B (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__B2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__I (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__S0 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__S1 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__S0 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__S1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__S0 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__S1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__I0 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__I1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__S0 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A4 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__B (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__B (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__B2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__S1 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(\reg_file.reg_storage[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__S0 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__S1 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__I1 (.I(\reg_file.reg_storage[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__I2 (.I(\reg_file.reg_storage[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__S1 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__S0 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__S1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__B (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__S (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I0 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__I (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__B (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__C (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__I (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__I3 (.I(\reg_file.reg_storage[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__S0 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__S1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__I (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__B (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__I (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__S0 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__S1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__S0 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__S1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__S0 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__S1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A2 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__I (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A4 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__B (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__S (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__B (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__B (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__B2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__I (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__I3 (.I(\reg_file.reg_storage[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__S0 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__S1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__B (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__S0 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__S1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S0 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__S0 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__S1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__I (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__C (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__B1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__C (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__I3 (.I(\reg_file.reg_storage[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__S0 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__S1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__B (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__S0 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__S1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__I3 (.I(\reg_file.reg_storage[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__S0 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__S1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__I (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__S1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__S (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__B (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__B2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__I (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__I (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__I (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__I (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__I2 (.I(\reg_file.reg_storage[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__I3 (.I(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__S1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__I (.I(\reg_file.reg_storage[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__I (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__S0 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__S1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__S0 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__S1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__S1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__B (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__S (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__I0 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__I (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I1 (.I(\reg_file.reg_storage[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I2 (.I(\reg_file.reg_storage[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I3 (.I(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__S0 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__S1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__I (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A1 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__B (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I1 (.I(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I2 (.I(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__S0 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__S1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I2 (.I(\reg_file.reg_storage[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I3 (.I(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__S0 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__S1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__S1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__B (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__B (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__S (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__C (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__C (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__B2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__B1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__I (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__I2 (.I(\reg_file.reg_storage[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__I (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A1 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__S1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__S1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__I1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__S1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__B (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__I (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__S (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__S (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__C (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__B (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__B2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__I2 (.I(\reg_file.reg_storage[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__S0 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__I (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__I1 (.I(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__S0 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__S0 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__I1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__S0 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__B (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__S (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__S (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__C (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__B2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__I (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__I2 (.I(\reg_file.reg_storage[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__S0 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__S1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__I1 (.I(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__I2 (.I(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__S1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__S0 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__S1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__I (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__S0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__C (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__B (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__I (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__B (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__B (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__B2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I1 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__S (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__C (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__C (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__I (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I2 (.I(\reg_file.reg_storage[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I3 (.I(\reg_file.reg_storage[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__S0 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__I (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__S0 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__S1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__S0 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__S0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__S1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__I (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__B (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__B (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__B (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__B2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__B (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__C (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__I (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__I3 (.I(\reg_file.reg_storage[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__S0 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__S0 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__S0 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__I1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__S0 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__I (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__B (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__C (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__B2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__B (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__I (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A2 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I2 (.I(\reg_file.reg_storage[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I3 (.I(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__S0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__I1 (.I(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__I2 (.I(\reg_file.reg_storage[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__S0 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__I2 (.I(\reg_file.reg_storage[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__S0 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__S0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__S1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__I (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__C (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__B (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__C (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__B2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A2 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A1 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__I2 (.I(\reg_file.reg_storage[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__I3 (.I(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__S0 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__I1 (.I(\reg_file.reg_storage[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__I2 (.I(\reg_file.reg_storage[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__S0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__I1 (.I(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__I2 (.I(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__S0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__S0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__S1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__B (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__C (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A2 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__B (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__C (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A2 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__C (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__C2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__B (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A2 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A3 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A1 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__B (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__B2 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__B (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__B (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A3 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__C (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__C (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__B (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A2 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__B (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A2 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__C (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__C (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__B (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A2 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__B (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__B (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__I (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A2 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__I (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__I (.I(\pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__B1 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__I (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__I (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__I (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__I (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__I (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__B1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__I (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__B1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__I (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__I (.I(\pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__B1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__I (.I(\pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__I (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__B1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__I (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__A2 (.I(\pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(\pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A2 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__I (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__B2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__I (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__B1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__I (.I(\pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__B1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__I (.I(\pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__B (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__B2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__I (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A2 (.I(\pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A1 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__B1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__B1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(\pc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A3 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__I (.I(\pc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A1 (.I(\pc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__B1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A1 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__B1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__I (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__B1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A1 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__C (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__B1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__B1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__B1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__B1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__B1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(\pc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(\pc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__B1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A1 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__I (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__I (.I(\pc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__I (.I(\pc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A1 (.I(\pc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A3 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__B1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(\pc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__I (.I(\pc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__B (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A1 (.I(\pc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__I (.I(\pc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(\pc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__B1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I (.I(\pc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A1 (.I(\pc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__B1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I (.I(\pc[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A2 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__B (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(\pc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A2 (.I(\pc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__B2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__B1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__B2 (.I(\pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I0 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__B (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__I (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__I (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__S (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__B1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__I (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__S (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__I (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__I (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__B2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__I (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__S (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__B (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__I (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__S (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__I (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__I (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__B (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__I (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__I (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__B (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__B (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__I (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__B2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__I (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__I (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__I (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__I (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__B2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__I (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(\reg_file.reg_storage[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__B2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__I (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A1 (.I(\reg_file.reg_storage[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__B2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__I (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__I (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__B1 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__B2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__I (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__I (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__B1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__B2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__C (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__I (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__B1 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__B2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__C (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__B1 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__C (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__A1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__I (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__C (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__I (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__I (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__I (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__I (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__C (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(\reg_file.reg_storage[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A1 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__I (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__C (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__I (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A1 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__I (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__C (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__I (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__C (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__I (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__I (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__I (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__B1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__I (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__C (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__B2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__C (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__I (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__S (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__I0 (.I(\reg_file.reg_storage[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__S (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__S (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__S (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__I (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__I (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__I (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A1 (.I(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A1 (.I(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A1 (.I(\reg_file.reg_storage[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__I (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A1 (.I(\reg_file.reg_storage[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__I (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(\reg_file.reg_storage[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A1 (.I(\reg_file.reg_storage[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A2 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A1 (.I(\reg_file.reg_storage[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A2 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A2 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A1 (.I(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A1 (.I(\reg_file.reg_storage[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A1 (.I(\reg_file.reg_storage[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A1 (.I(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__I (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__S (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__S (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__S (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__S (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__I (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__I (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__I (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A1 (.I(\reg_file.reg_storage[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__I (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__I (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__A1 (.I(\reg_file.reg_storage[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__I (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__I (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__I (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__I (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A1 (.I(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__I (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__I (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__S (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__I (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__S (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__S (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__S (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__I (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__I (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__I (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A2 (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__A2 (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A2 (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A2 (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__I (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__I (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A1 (.I(\reg_file.reg_storage[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__I (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__I (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(\reg_file.reg_storage[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__I (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A2 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A2 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__A2 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A2 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__I (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__I (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A1 (.I(\reg_file.reg_storage[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__I (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__I (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A2 (.I(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A1 (.I(\reg_file.reg_storage[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A2 (.I(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A1 (.I(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A2 (.I(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__I (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__S (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__S (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__I (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__S (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__I (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__I1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__S (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__I (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__I (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__I (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__I (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__I (.I(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__I (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__I (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__I (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__I (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__I (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__I (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A1 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__I (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__I (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__I (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__I (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__I (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__I (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__I (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__I (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__I (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(\reg_file.reg_storage[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__I (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__I (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A1 (.I(\reg_file.reg_storage[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__I (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__I (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A1 (.I(\reg_file.reg_storage[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__I (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__I (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__I (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__I (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__I (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__I (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__I (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__I (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A2 (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A2 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__I (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A2 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__A2 (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A2 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__I (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A2 (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A1 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A2 (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__I (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__I (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__I (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__I (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A1 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__I (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__I (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__I (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__I (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__I (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__I (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A2 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__I (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A2 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A1 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A2 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__I (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__I (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__S (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__S (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__I1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__S (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__I (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__I (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__I (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A1 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__I (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__I (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A1 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A1 (.I(\reg_file.reg_storage[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__I (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__I (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A1 (.I(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__I (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__I (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__I (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__I (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__I (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__I (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A1 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__I (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__I (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A1 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__S (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__S (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__S (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__I1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__S (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__I (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__I (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__A1 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__I (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__I (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A1 (.I(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__I (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__I (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A1 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__I (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A1 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__I (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A1 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__S (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__S (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__S (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__I1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__S (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__I (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A2 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A1 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A2 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A2 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A1 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__I (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A1 (.I(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A1 (.I(\reg_file.reg_storage[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__I (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A1 (.I(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__I (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__I (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__I (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A2 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__A2 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A2 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A1 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__I (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A1 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__I (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__A1 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__I (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__S (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__I (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__I (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__I1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__S (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__I (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__I (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__I (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(\reg_file.reg_storage[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__I (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__I (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__I (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__I (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__I (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A1 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__I (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__I (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__I (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__I (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__I (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__I (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__I (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__I (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A1 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__I (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A1 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__I (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__I (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__I (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__I (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__I (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__I (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A1 (.I(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__I (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__I (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A1 (.I(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A1 (.I(\reg_file.reg_storage[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__I (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__S (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__S (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__S (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__I1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__S (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__I (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__I (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__I (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(\reg_file.reg_storage[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__I (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__I (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A1 (.I(\reg_file.reg_storage[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__I (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__A1 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__I (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__I (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A1 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__I (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__I (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__A1 (.I(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A1 (.I(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__I (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A1 (.I(\reg_file.reg_storage[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(\reg_file.reg_storage[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__S (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__S (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__S (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__I1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__S (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__I (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__I (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A1 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A1 (.I(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__I (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A1 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__I (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A1 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__I (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A2 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A2 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A2 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A1 (.I(\reg_file.reg_storage[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A2 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A1 (.I(\reg_file.reg_storage[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A1 (.I(\reg_file.reg_storage[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A1 (.I(\reg_file.reg_storage[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A1 (.I(\reg_file.reg_storage[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A1 (.I(\reg_file.reg_storage[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A1 (.I(\reg_file.reg_storage[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A1 (.I(\reg_file.reg_storage[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__B1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__B1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__S (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__S (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__S (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__I1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__S (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__I (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A1 (.I(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A1 (.I(\reg_file.reg_storage[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A1 (.I(\reg_file.reg_storage[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__I (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A1 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__I (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A1 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__I (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A1 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A1 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__I (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A2 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A2 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A1 (.I(\reg_file.reg_storage[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A1 (.I(\reg_file.reg_storage[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A1 (.I(\reg_file.reg_storage[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A1 (.I(\reg_file.reg_storage[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__A1 (.I(\reg_file.reg_storage[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__I (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__S (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__I1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__S (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__S (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__S (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__I (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A1 (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A1 (.I(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A1 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A1 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__I (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A1 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__I (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A1 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A1 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(\reg_file.reg_storage[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A1 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__I (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__I (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A1 (.I(\reg_file.reg_storage[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A1 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__I (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A1 (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__I (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A1 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A1 (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A1 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__I (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__S (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__I1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__S (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__S (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__S (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__I (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__I (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A1 (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A1 (.I(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__A1 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A1 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A1 (.I(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A1 (.I(\reg_file.reg_storage[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__A1 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__A1 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A1 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A1 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__A1 (.I(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A1 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A1 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__I (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__A1 (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__I (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__A2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A1 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A1 (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__A1 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__A2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__I (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__S (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__I1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__S (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__S (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__S (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__I (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__I (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__I (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A1 (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__A1 (.I(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__A1 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A1 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__I (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__I (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__A1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__A1 (.I(\reg_file.reg_storage[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__A1 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__I (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__I (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__A1 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__A1 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A1 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A1 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__I (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__I (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A1 (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A1 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__I (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__I (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A1 (.I(\reg_file.reg_storage[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8717__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__A1 (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__I (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A2 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__A2 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__A2 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__A1 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__A2 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A2 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A1 (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A2 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A2 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A1 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A2 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__CLK (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8881__CLK (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9215__CLK (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(inst_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(inst_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(inst_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(inst_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(inst_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(inst_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(inst_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(inst_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(inst_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(inst_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(inst_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(inst_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(inst_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(inst_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(inst_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(inst_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(inst_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(inst_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(inst_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(inst_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(inst_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(inst_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(inst_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(inst_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(inst_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(mem_load_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(mem_load_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(mem_load_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(mem_load_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(mem_load_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(mem_load_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(mem_load_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(inst_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(mem_load_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(mem_load_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(mem_load_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(mem_load_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(mem_load_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(mem_load_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(mem_load_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(mem_load_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(mem_load_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(mem_load_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(inst_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(mem_load_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(mem_load_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(mem_load_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(mem_load_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(mem_load_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(mem_load_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(mem_load_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(mem_load_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(mem_load_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(mem_load_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(inst_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(mem_load_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(mem_load_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(mem_load_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(mem_load_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(mem_load_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(inst_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(inst_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(inst_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(inst_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output85_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output87_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output88_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output89_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer14_I (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer16_I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer17_I (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer18_I (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer3_I (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer8_I (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4334_ (.I(net6),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _4335_ (.I(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4336_ (.I(net27),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4337_ (.I(net28),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4338_ (.I(net29),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4339_ (.A1(_0484_),
    .A2(_0485_),
    .A3(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4340_ (.I(net26),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4341_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4342_ (.I(net23),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4343_ (.I(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4344_ (.A1(_0489_),
    .A2(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4345_ (.I(net26),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4346_ (.I(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4347_ (.I(net23),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4348_ (.I(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4349_ (.A1(net28),
    .A2(net29),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _4350_ (.A1(_0494_),
    .A2(_0496_),
    .A3(_0484_),
    .A4(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4351_ (.I(net29),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4352_ (.I(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4353_ (.I(_0500_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4354_ (.I(net27),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4355_ (.A1(_0493_),
    .A2(_0490_),
    .A3(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4356_ (.A1(_0485_),
    .A2(_0501_),
    .B(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4357_ (.A1(_0487_),
    .A2(_0492_),
    .B(_0498_),
    .C(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4358_ (.A1(_0483_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4359_ (.I(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4360_ (.I(net27),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4361_ (.I(net28),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4362_ (.A1(_0508_),
    .A2(_0509_),
    .A3(_0499_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4363_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4364_ (.A1(_0493_),
    .A2(_0496_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4365_ (.A1(net26),
    .A2(_0495_),
    .A3(_0484_),
    .A4(_0497_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4366_ (.I(_0486_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4367_ (.A1(net26),
    .A2(net23),
    .A3(_0508_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4368_ (.I(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4369_ (.A1(_0509_),
    .A2(_0514_),
    .B(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4370_ (.A1(_0511_),
    .A2(_0512_),
    .B(net106),
    .C(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4371_ (.I(net5),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4372_ (.A1(_0485_),
    .A2(_0514_),
    .A3(_0503_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4373_ (.A1(_0519_),
    .A2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4374_ (.A1(net4),
    .A2(_0518_),
    .B1(_0521_),
    .B2(net6),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4375_ (.I(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4376_ (.A1(_0509_),
    .A2(_0501_),
    .A3(_0516_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4377_ (.A1(net5),
    .A2(_0518_),
    .B(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4378_ (.A1(_0523_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4379_ (.A1(net24),
    .A2(_0518_),
    .B1(_0524_),
    .B2(_0483_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4380_ (.A1(_0507_),
    .A2(_0526_),
    .B(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4381_ (.I(net24),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4382_ (.I(_0520_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4383_ (.A1(_0529_),
    .A2(_0505_),
    .B1(_0530_),
    .B2(_0482_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4384_ (.A1(_0482_),
    .A2(_0518_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4385_ (.A1(_0519_),
    .A2(_0505_),
    .B(_0530_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4386_ (.A1(_0531_),
    .A2(_0532_),
    .A3(_0523_),
    .A4(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4387_ (.I(net4),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4388_ (.A1(_0483_),
    .A2(_0519_),
    .A3(_0530_),
    .B1(_0505_),
    .B2(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4389_ (.I(_0525_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4390_ (.A1(_0507_),
    .A2(_0536_),
    .A3(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4391_ (.A1(_0528_),
    .A2(_0534_),
    .A3(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4392_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4393_ (.A1(_0502_),
    .A2(_0485_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4394_ (.A1(_0493_),
    .A2(_0490_),
    .A3(_0486_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4395_ (.A1(_0510_),
    .A2(_0512_),
    .B1(_0541_),
    .B2(_0542_),
    .C(_0513_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4396_ (.I(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4397_ (.I(net13),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4398_ (.I(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4399_ (.I(net114),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4400_ (.I(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4401_ (.A1(_0500_),
    .A2(_0515_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4402_ (.A1(_0490_),
    .A2(_0508_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4403_ (.A1(_0486_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4404_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4405_ (.A1(_0488_),
    .A2(_0508_),
    .A3(_0499_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _4406_ (.A1(_0548_),
    .A2(net108),
    .A3(_0552_),
    .A4(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4407_ (.A1(_0544_),
    .A2(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _4408_ (.I(net16),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4409_ (.I(net15),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4410_ (.I(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4411_ (.I(net14),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4412_ (.I(_0546_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4413_ (.A1(_0559_),
    .A2(_0560_),
    .A3(net17),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4414_ (.A1(_0556_),
    .A2(_0558_),
    .A3(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4415_ (.I(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4416_ (.I(_0545_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4417_ (.I(net14),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4418_ (.I(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4419_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(\reg_file.reg_storage[5][0] ),
    .I2(\reg_file.reg_storage[6][0] ),
    .I3(\reg_file.reg_storage[7][0] ),
    .S0(_0564_),
    .S1(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4420_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(\reg_file.reg_storage[3][0] ),
    .S(_0546_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4421_ (.I0(\reg_file.reg_storage[1][0] ),
    .I1(_0568_),
    .S(_0566_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4422_ (.I(_0565_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4423_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(\reg_file.reg_storage[13][0] ),
    .I2(\reg_file.reg_storage[14][0] ),
    .I3(\reg_file.reg_storage[15][0] ),
    .S0(_0564_),
    .S1(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4424_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(\reg_file.reg_storage[9][0] ),
    .I2(\reg_file.reg_storage[10][0] ),
    .I3(\reg_file.reg_storage[11][0] ),
    .S0(_0564_),
    .S1(_0570_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4425_ (.I(net16),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4426_ (.I0(_0567_),
    .I1(_0569_),
    .I2(_0571_),
    .I3(_0572_),
    .S0(_0558_),
    .S1(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _4427_ (.A1(_0544_),
    .A2(_0563_),
    .A3(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _4428_ (.A1(_0555_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4429_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4430_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4431_ (.A1(_0491_),
    .A2(_0514_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4432_ (.A1(_0511_),
    .A2(_0579_),
    .B(_0489_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4433_ (.I(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4434_ (.I(_0487_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4435_ (.A1(_0496_),
    .A2(_0501_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4436_ (.I(net10),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4437_ (.A1(_0584_),
    .A2(net9),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4438_ (.I(net8),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4439_ (.I(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4440_ (.I(net7),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4441_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4442_ (.A1(_0587_),
    .A2(_0589_),
    .A3(net11),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4443_ (.A1(_0582_),
    .A2(_0583_),
    .B1(_0585_),
    .B2(_0590_),
    .C(_0494_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4444_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4445_ (.I(net7),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4446_ (.I(_0593_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4447_ (.I(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4448_ (.I(_0587_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4449_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(\reg_file.reg_storage[5][0] ),
    .I2(\reg_file.reg_storage[6][0] ),
    .I3(\reg_file.reg_storage[7][0] ),
    .S0(_0595_),
    .S1(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4450_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(\reg_file.reg_storage[3][0] ),
    .S(_0589_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4451_ (.I(_0586_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4452_ (.I0(\reg_file.reg_storage[1][0] ),
    .I1(_0598_),
    .S(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4453_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(\reg_file.reg_storage[13][0] ),
    .I2(\reg_file.reg_storage[14][0] ),
    .I3(\reg_file.reg_storage[15][0] ),
    .S0(_0595_),
    .S1(_0599_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4454_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(\reg_file.reg_storage[9][0] ),
    .I2(\reg_file.reg_storage[10][0] ),
    .I3(\reg_file.reg_storage[11][0] ),
    .S0(_0595_),
    .S1(_0599_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4455_ (.I(net9),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4456_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4457_ (.I(_0584_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4458_ (.I0(_0597_),
    .I1(_0600_),
    .I2(_0601_),
    .I3(_0602_),
    .S0(_0604_),
    .S1(_0605_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4459_ (.A1(\pc[0] ),
    .A2(_0581_),
    .B1(_0592_),
    .B2(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4460_ (.A1(_0578_),
    .A2(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4461_ (.I(_0580_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4462_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4463_ (.I(_0584_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4464_ (.I(_0603_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4465_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4466_ (.I(_0586_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4467_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4468_ (.I0(\reg_file.reg_storage[2][1] ),
    .I1(\reg_file.reg_storage[3][1] ),
    .S(_0589_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4469_ (.I(net8),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4470_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4471_ (.A1(_0618_),
    .A2(\reg_file.reg_storage[1][1] ),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4472_ (.A1(_0615_),
    .A2(_0616_),
    .B(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4473_ (.I(_0586_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4474_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(\reg_file.reg_storage[5][1] ),
    .I2(\reg_file.reg_storage[6][1] ),
    .I3(\reg_file.reg_storage[7][1] ),
    .S0(_0594_),
    .S1(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4475_ (.A1(_0612_),
    .A2(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4476_ (.A1(_0613_),
    .A2(_0620_),
    .B(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4477_ (.A1(_0611_),
    .A2(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4478_ (.A1(_0582_),
    .A2(_0583_),
    .B(_0494_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4479_ (.A1(_0585_),
    .A2(_0590_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_0626_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4481_ (.I(net10),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4482_ (.I(_0593_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4483_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(\reg_file.reg_storage[13][1] ),
    .I2(\reg_file.reg_storage[14][1] ),
    .I3(\reg_file.reg_storage[15][1] ),
    .S0(_0630_),
    .S1(_0618_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4484_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(\reg_file.reg_storage[9][1] ),
    .I2(\reg_file.reg_storage[10][1] ),
    .I3(\reg_file.reg_storage[11][1] ),
    .S0(_0594_),
    .S1(_0621_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4485_ (.I0(_0631_),
    .I1(_0632_),
    .S(_0612_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4486_ (.A1(_0629_),
    .A2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4487_ (.A1(_0625_),
    .A2(_0628_),
    .A3(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4488_ (.A1(\pc[1] ),
    .A2(_0610_),
    .B(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4489_ (.I(_0543_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4490_ (.I0(_0516_),
    .I1(_0550_),
    .S(_0500_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4491_ (.I(_0565_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4492_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4493_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4494_ (.A1(net31),
    .A2(_0549_),
    .B1(_0638_),
    .B2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4495_ (.A1(_0637_),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4496_ (.I(net13),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4497_ (.I(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4498_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(\reg_file.reg_storage[5][1] ),
    .I2(\reg_file.reg_storage[6][1] ),
    .I3(\reg_file.reg_storage[7][1] ),
    .S0(_0645_),
    .S1(_0559_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4499_ (.I0(\reg_file.reg_storage[2][1] ),
    .I1(\reg_file.reg_storage[3][1] ),
    .S(net113),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4500_ (.I0(\reg_file.reg_storage[1][1] ),
    .I1(_0647_),
    .S(_0559_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4501_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(\reg_file.reg_storage[13][1] ),
    .I2(\reg_file.reg_storage[14][1] ),
    .I3(\reg_file.reg_storage[15][1] ),
    .S0(_0645_),
    .S1(_0566_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4502_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(\reg_file.reg_storage[9][1] ),
    .I2(\reg_file.reg_storage[10][1] ),
    .I3(\reg_file.reg_storage[11][1] ),
    .S0(_0645_),
    .S1(_0566_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4503_ (.I0(_0646_),
    .I1(_0648_),
    .I2(_0649_),
    .I3(_0650_),
    .S0(_0558_),
    .S1(_0573_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _4504_ (.A1(_0544_),
    .A2(_0563_),
    .A3(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4505_ (.A1(_0652_),
    .A2(_0643_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4506_ (.I(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4507_ (.A1(_0531_),
    .A2(_0532_),
    .A3(_0522_),
    .A4(_0525_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4508_ (.I(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4509_ (.A1(_0577_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4510_ (.A1(_0636_),
    .A2(_0654_),
    .A3(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4511_ (.I(_0656_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4512_ (.A1(_0577_),
    .A2(_0659_),
    .B(_0654_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4513_ (.I(_0655_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4514_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4515_ (.A1(_0654_),
    .A2(_0577_),
    .A3(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4516_ (.I(\pc[1] ),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4517_ (.A1(_0625_),
    .A2(_0628_),
    .A3(_0634_),
    .B1(_0626_),
    .B2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4518_ (.I(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4519_ (.A1(_0660_),
    .A2(_0663_),
    .B(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4520_ (.A1(_0608_),
    .A2(_0658_),
    .B(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4521_ (.I(\pc[2] ),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4522_ (.I(_0609_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4523_ (.I(_0591_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4524_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4525_ (.I(_0630_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4526_ (.I(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4527_ (.I(_0617_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4528_ (.I(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4529_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(\reg_file.reg_storage[5][2] ),
    .I2(\reg_file.reg_storage[6][2] ),
    .I3(\reg_file.reg_storage[7][2] ),
    .S0(_0674_),
    .S1(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4530_ (.I(_0593_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4531_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(\reg_file.reg_storage[3][2] ),
    .S(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4532_ (.I(_0599_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4533_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_0679_),
    .S(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4534_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(\reg_file.reg_storage[13][2] ),
    .I2(\reg_file.reg_storage[14][2] ),
    .I3(\reg_file.reg_storage[15][2] ),
    .S0(_0674_),
    .S1(_0680_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4535_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(\reg_file.reg_storage[9][2] ),
    .I2(\reg_file.reg_storage[10][2] ),
    .I3(\reg_file.reg_storage[11][2] ),
    .S0(_0674_),
    .S1(_0680_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4536_ (.I(_0604_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4537_ (.I(_0584_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4538_ (.I(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4539_ (.I0(_0677_),
    .I1(_0681_),
    .I2(_0682_),
    .I3(_0683_),
    .S0(_0684_),
    .S1(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4540_ (.A1(_0669_),
    .A2(_0670_),
    .B1(_0672_),
    .B2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4541_ (.A1(_0541_),
    .A2(_0542_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4542_ (.A1(_0487_),
    .A2(_0492_),
    .B(_0498_),
    .C(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4543_ (.I(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4544_ (.I(_0557_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4545_ (.I(_0549_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4546_ (.A1(net32),
    .A2(_0514_),
    .A3(_0503_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4547_ (.A1(_0692_),
    .A2(_0693_),
    .A3(_0552_),
    .B(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4548_ (.A1(_0691_),
    .A2(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4549_ (.I(_0544_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4550_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4551_ (.I(_0639_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4552_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(\reg_file.reg_storage[5][2] ),
    .I2(\reg_file.reg_storage[6][2] ),
    .I3(\reg_file.reg_storage[7][2] ),
    .S0(_0560_),
    .S1(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4553_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(\reg_file.reg_storage[3][2] ),
    .S(_0564_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4554_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_0701_),
    .S(_0699_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4555_ (.I(net14),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4556_ (.I(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4557_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(\reg_file.reg_storage[13][2] ),
    .I2(\reg_file.reg_storage[14][2] ),
    .I3(\reg_file.reg_storage[15][2] ),
    .S0(_0560_),
    .S1(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4558_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(\reg_file.reg_storage[9][2] ),
    .I2(\reg_file.reg_storage[10][2] ),
    .I3(\reg_file.reg_storage[11][2] ),
    .S0(_0560_),
    .S1(_0704_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4559_ (.I(_0557_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4560_ (.I(net16),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4561_ (.I0(_0700_),
    .I1(_0702_),
    .I2(_0705_),
    .I3(_0706_),
    .S0(_0707_),
    .S1(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4562_ (.A1(_0698_),
    .A2(_0563_),
    .A3(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4563_ (.A1(_0696_),
    .A2(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4564_ (.A1(_0653_),
    .A2(_0576_),
    .B(_0661_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4565_ (.A1(_0711_),
    .A2(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4566_ (.A1(_0688_),
    .A2(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4567_ (.A1(_0668_),
    .A2(_0714_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4568_ (.I(_0539_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4569_ (.A1(_0690_),
    .A2(_0695_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4570_ (.A1(_0637_),
    .A2(_0563_),
    .A3(_0709_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4571_ (.A1(_0718_),
    .A2(_0717_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4572_ (.I(_0719_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4573_ (.I(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4574_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4575_ (.I(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4576_ (.I(_0578_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4577_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4578_ (.I(_0671_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4579_ (.I(_0593_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4580_ (.I(_0621_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4581_ (.I0(\reg_file.reg_storage[4][9] ),
    .I1(\reg_file.reg_storage[5][9] ),
    .I2(\reg_file.reg_storage[6][9] ),
    .I3(\reg_file.reg_storage[7][9] ),
    .S0(_0727_),
    .S1(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4582_ (.I(_0614_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4583_ (.I(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4584_ (.I(\reg_file.reg_storage[1][9] ),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4585_ (.I(_0595_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4586_ (.A1(_0733_),
    .A2(\reg_file.reg_storage[3][9] ),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4587_ (.I(_0588_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4588_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4589_ (.A1(_0736_),
    .A2(\reg_file.reg_storage[2][9] ),
    .B(_0615_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4590_ (.A1(_0731_),
    .A2(_0732_),
    .B1(_0734_),
    .B2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4591_ (.I(_0594_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4592_ (.I(_0587_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4593_ (.I0(\reg_file.reg_storage[12][9] ),
    .I1(\reg_file.reg_storage[13][9] ),
    .I2(\reg_file.reg_storage[14][9] ),
    .I3(\reg_file.reg_storage[15][9] ),
    .S0(_0739_),
    .S1(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4594_ (.I0(\reg_file.reg_storage[8][9] ),
    .I1(\reg_file.reg_storage[9][9] ),
    .I2(\reg_file.reg_storage[10][9] ),
    .I3(\reg_file.reg_storage[11][9] ),
    .S0(_0739_),
    .S1(_0740_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4595_ (.I0(_0729_),
    .I1(_0738_),
    .I2(_0741_),
    .I3(_0742_),
    .S0(_0613_),
    .S1(_0611_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4596_ (.A1(\pc[9] ),
    .A2(_0610_),
    .B1(_0726_),
    .B2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4597_ (.I(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4598_ (.I(_0745_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4599_ (.A1(_0725_),
    .A2(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4600_ (.A1(_0555_),
    .A2(_0575_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4601_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4602_ (.I(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4603_ (.I(_0609_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4604_ (.I(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4605_ (.I(_0671_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4606_ (.I(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4607_ (.I(_0588_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4608_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4609_ (.I(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4610_ (.I(_0621_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4611_ (.I(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4612_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(\reg_file.reg_storage[5][8] ),
    .I2(\reg_file.reg_storage[6][8] ),
    .I3(\reg_file.reg_storage[7][8] ),
    .S0(_0757_),
    .S1(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4613_ (.I(_0730_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4614_ (.I(_0761_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4615_ (.I(\reg_file.reg_storage[1][8] ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4616_ (.I(_0630_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4617_ (.I(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4618_ (.I(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(_0766_),
    .A2(\reg_file.reg_storage[3][8] ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4620_ (.I(_0735_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4621_ (.I(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4622_ (.I(_0614_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4623_ (.I(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4624_ (.I(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4625_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][8] ),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4626_ (.A1(_0762_),
    .A2(_0763_),
    .B1(_0767_),
    .B2(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4627_ (.I(_0756_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4628_ (.I(_0728_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4629_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(\reg_file.reg_storage[13][8] ),
    .I2(\reg_file.reg_storage[14][8] ),
    .I3(\reg_file.reg_storage[15][8] ),
    .S0(_0775_),
    .S1(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4630_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(\reg_file.reg_storage[9][8] ),
    .I2(\reg_file.reg_storage[10][8] ),
    .I3(\reg_file.reg_storage[11][8] ),
    .S0(_0757_),
    .S1(_0759_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4631_ (.I(_0684_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4632_ (.I(_0611_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4633_ (.I0(_0760_),
    .I1(_0774_),
    .I2(_0777_),
    .I3(_0778_),
    .S0(_0779_),
    .S1(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4634_ (.A1(\pc[8] ),
    .A2(_0752_),
    .B1(_0754_),
    .B2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4635_ (.I(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4636_ (.A1(_0750_),
    .A2(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4637_ (.A1(_0747_),
    .A2(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4638_ (.I(_0578_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4639_ (.I(\pc[7] ),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4640_ (.I(_0751_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4641_ (.I(_0753_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4642_ (.I(_0676_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4643_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(\reg_file.reg_storage[5][7] ),
    .I2(\reg_file.reg_storage[6][7] ),
    .I3(\reg_file.reg_storage[7][7] ),
    .S0(_0766_),
    .S1(_0790_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4644_ (.I(_0772_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4645_ (.I(\reg_file.reg_storage[1][7] ),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4646_ (.I(_0733_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4647_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4648_ (.A1(_0795_),
    .A2(\reg_file.reg_storage[3][7] ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4649_ (.I(_0768_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4650_ (.A1(_0797_),
    .A2(\reg_file.reg_storage[2][7] ),
    .B(_0762_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4651_ (.A1(_0792_),
    .A2(_0793_),
    .B1(_0796_),
    .B2(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4652_ (.I(_0678_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4653_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(\reg_file.reg_storage[13][7] ),
    .I2(\reg_file.reg_storage[14][7] ),
    .I3(\reg_file.reg_storage[15][7] ),
    .S0(_0800_),
    .S1(_0790_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4654_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(\reg_file.reg_storage[9][7] ),
    .I2(\reg_file.reg_storage[10][7] ),
    .I3(\reg_file.reg_storage[11][7] ),
    .S0(_0766_),
    .S1(_0790_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4655_ (.I(_0603_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4656_ (.I(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4657_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4658_ (.I(_0686_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4659_ (.I0(_0791_),
    .I1(_0799_),
    .I2(_0801_),
    .I3(_0802_),
    .S0(_0805_),
    .S1(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4660_ (.A1(_0787_),
    .A2(_0788_),
    .B1(_0789_),
    .B2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4661_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_0786_),
    .A2(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4663_ (.I(_0749_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4664_ (.I(\pc[6] ),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4665_ (.I(_0674_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4666_ (.I(_0758_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4667_ (.I0(\reg_file.reg_storage[4][6] ),
    .I1(\reg_file.reg_storage[5][6] ),
    .I2(\reg_file.reg_storage[6][6] ),
    .I3(\reg_file.reg_storage[7][6] ),
    .S0(_0813_),
    .S1(_0814_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4668_ (.I(\reg_file.reg_storage[1][6] ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4669_ (.I(_0764_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4670_ (.A1(_0817_),
    .A2(\reg_file.reg_storage[3][6] ),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4671_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][6] ),
    .B(_0772_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4672_ (.A1(_0762_),
    .A2(_0816_),
    .B1(_0818_),
    .B2(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4673_ (.I0(\reg_file.reg_storage[12][6] ),
    .I1(\reg_file.reg_storage[13][6] ),
    .I2(\reg_file.reg_storage[14][6] ),
    .I3(\reg_file.reg_storage[15][6] ),
    .S0(_0757_),
    .S1(_0759_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4674_ (.I0(\reg_file.reg_storage[8][6] ),
    .I1(\reg_file.reg_storage[9][6] ),
    .I2(\reg_file.reg_storage[10][6] ),
    .I3(\reg_file.reg_storage[11][6] ),
    .S0(_0813_),
    .S1(_0759_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4675_ (.I0(_0815_),
    .I1(_0820_),
    .I2(_0821_),
    .I3(_0822_),
    .S0(_0779_),
    .S1(_0806_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4676_ (.A1(_0812_),
    .A2(_0752_),
    .B1(_0789_),
    .B2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4677_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4678_ (.A1(_0811_),
    .A2(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(_0810_),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4680_ (.A1(_0643_),
    .A2(_0652_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4681_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4682_ (.I(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4683_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4684_ (.I(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4685_ (.I(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4686_ (.I0(_0785_),
    .I1(_0827_),
    .S(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4687_ (.I(_0654_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4688_ (.I(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4689_ (.I(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4690_ (.I(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4691_ (.I(_0589_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4692_ (.I(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4693_ (.I(_0740_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4694_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(\reg_file.reg_storage[5][5] ),
    .I2(\reg_file.reg_storage[6][5] ),
    .I3(\reg_file.reg_storage[7][5] ),
    .S0(_0840_),
    .S1(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4695_ (.I(_0731_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4696_ (.I(\reg_file.reg_storage[1][5] ),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4697_ (.A1(_0800_),
    .A2(\reg_file.reg_storage[3][5] ),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4698_ (.I(_0768_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4699_ (.I(_0614_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4700_ (.I(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4701_ (.A1(_0846_),
    .A2(\reg_file.reg_storage[2][5] ),
    .B(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4702_ (.A1(_0843_),
    .A2(_0844_),
    .B1(_0845_),
    .B2(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4703_ (.I(_0839_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4704_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(\reg_file.reg_storage[13][5] ),
    .I2(\reg_file.reg_storage[14][5] ),
    .I3(\reg_file.reg_storage[15][5] ),
    .S0(_0851_),
    .S1(_0841_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4705_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(\reg_file.reg_storage[9][5] ),
    .I2(\reg_file.reg_storage[10][5] ),
    .I3(\reg_file.reg_storage[11][5] ),
    .S0(_0840_),
    .S1(_0841_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4706_ (.I(_0803_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4707_ (.I0(_0842_),
    .I1(_0850_),
    .I2(_0852_),
    .I3(_0853_),
    .S0(_0854_),
    .S1(_0780_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4708_ (.A1(\pc[5] ),
    .A2(_0752_),
    .B1(_0754_),
    .B2(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4709_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4710_ (.A1(_0786_),
    .A2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4711_ (.I(_0751_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4712_ (.I(_0726_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4713_ (.I(_0740_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4714_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(\reg_file.reg_storage[5][4] ),
    .I2(\reg_file.reg_storage[6][4] ),
    .I3(\reg_file.reg_storage[7][4] ),
    .S0(_0851_),
    .S1(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4715_ (.I(_0770_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4716_ (.I(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4717_ (.I(\reg_file.reg_storage[1][4] ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4718_ (.A1(_0800_),
    .A2(\reg_file.reg_storage[3][4] ),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4719_ (.I(_0847_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4720_ (.A1(_0846_),
    .A2(\reg_file.reg_storage[2][4] ),
    .B(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4721_ (.A1(_0864_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4722_ (.I(_0839_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4723_ (.I(_0728_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4724_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(\reg_file.reg_storage[13][4] ),
    .I2(\reg_file.reg_storage[14][4] ),
    .I3(\reg_file.reg_storage[15][4] ),
    .S0(_0870_),
    .S1(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4725_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(\reg_file.reg_storage[9][4] ),
    .I2(\reg_file.reg_storage[10][4] ),
    .I3(\reg_file.reg_storage[11][4] ),
    .S0(_0870_),
    .S1(_0871_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4726_ (.I(_0605_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4727_ (.I0(_0862_),
    .I1(_0869_),
    .I2(_0872_),
    .I3(_0873_),
    .S0(_0854_),
    .S1(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4728_ (.A1(\pc[4] ),
    .A2(_0859_),
    .B1(_0860_),
    .B2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4729_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4730_ (.A1(_0811_),
    .A2(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4731_ (.A1(_0858_),
    .A2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4732_ (.I(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4733_ (.I(_0837_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4734_ (.I(_0811_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4735_ (.I(_0688_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4736_ (.A1(_0882_),
    .A2(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4737_ (.I(_0786_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4738_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(\reg_file.reg_storage[5][3] ),
    .I2(\reg_file.reg_storage[6][3] ),
    .I3(\reg_file.reg_storage[7][3] ),
    .S0(_0840_),
    .S1(_0841_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4739_ (.I(\reg_file.reg_storage[1][3] ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(_0800_),
    .A2(\reg_file.reg_storage[3][3] ),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4741_ (.A1(_0846_),
    .A2(\reg_file.reg_storage[2][3] ),
    .B(_0848_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4742_ (.A1(_0843_),
    .A2(_0887_),
    .B1(_0888_),
    .B2(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4743_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(\reg_file.reg_storage[13][3] ),
    .I2(\reg_file.reg_storage[14][3] ),
    .I3(\reg_file.reg_storage[15][3] ),
    .S0(_0851_),
    .S1(_0861_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4744_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(\reg_file.reg_storage[9][3] ),
    .I2(\reg_file.reg_storage[10][3] ),
    .I3(\reg_file.reg_storage[11][3] ),
    .S0(_0851_),
    .S1(_0861_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4745_ (.I0(_0886_),
    .I1(_0890_),
    .I2(_0891_),
    .I3(_0892_),
    .S0(_0854_),
    .S1(_0780_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4746_ (.A1(\pc[3] ),
    .A2(_0859_),
    .B1(_0860_),
    .B2(_0893_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4747_ (.I(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4748_ (.I(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4749_ (.A1(_0885_),
    .A2(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_0884_),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4751_ (.A1(_0881_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4752_ (.I(_0720_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4753_ (.I(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4754_ (.A1(_0838_),
    .A2(_0880_),
    .B(_0899_),
    .C(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4755_ (.A1(_0543_),
    .A2(_0562_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4756_ (.I(_0557_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4757_ (.I(_0545_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4758_ (.I(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4759_ (.I(_0639_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4760_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(\reg_file.reg_storage[5][3] ),
    .I2(\reg_file.reg_storage[6][3] ),
    .I3(\reg_file.reg_storage[7][3] ),
    .S0(_0906_),
    .S1(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4761_ (.A1(_0904_),
    .A2(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4762_ (.I(net112),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4763_ (.A1(_0910_),
    .A2(\reg_file.reg_storage[3][3] ),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4764_ (.I(_0703_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4765_ (.I(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4766_ (.A1(_0548_),
    .A2(\reg_file.reg_storage[2][3] ),
    .B(_0911_),
    .C(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4767_ (.I(_0704_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4768_ (.A1(_0915_),
    .A2(\reg_file.reg_storage[1][3] ),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4769_ (.A1(_0914_),
    .A2(_0916_),
    .B(_0692_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4770_ (.I(_0708_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4771_ (.A1(_0909_),
    .A2(_0917_),
    .B(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4772_ (.I(_0558_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4773_ (.I(_0905_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4774_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(\reg_file.reg_storage[13][3] ),
    .I2(\reg_file.reg_storage[14][3] ),
    .I3(\reg_file.reg_storage[15][3] ),
    .S0(_0921_),
    .S1(_0640_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4775_ (.A1(_0920_),
    .A2(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4776_ (.I(_0905_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4777_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(\reg_file.reg_storage[9][3] ),
    .I2(\reg_file.reg_storage[10][3] ),
    .I3(\reg_file.reg_storage[11][3] ),
    .S0(_0924_),
    .S1(_0699_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4778_ (.A1(net15),
    .A2(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4779_ (.A1(_0923_),
    .A2(_0926_),
    .B(_0556_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4780_ (.I(_0573_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4781_ (.A1(_0928_),
    .A2(_0638_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4782_ (.A1(net2),
    .A2(net109),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4783_ (.A1(_0929_),
    .A2(_0930_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _4784_ (.A1(_0903_),
    .A2(_0919_),
    .A3(_0927_),
    .B1(_0931_),
    .B2(_0697_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4785_ (.I(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4786_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4787_ (.A1(_0723_),
    .A2(_0834_),
    .B(_0902_),
    .C(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4788_ (.I(_0933_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4789_ (.I(_0711_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4790_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4791_ (.I(_0610_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4792_ (.I(_0726_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4793_ (.I(_0755_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4794_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4795_ (.I(_0675_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4796_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(\reg_file.reg_storage[5][13] ),
    .I2(\reg_file.reg_storage[6][13] ),
    .I3(\reg_file.reg_storage[7][13] ),
    .S0(_0942_),
    .S1(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4797_ (.I(_0771_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4798_ (.I(\reg_file.reg_storage[1][13] ),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4799_ (.A1(_0794_),
    .A2(\reg_file.reg_storage[3][13] ),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4800_ (.I(_0735_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4801_ (.I(_0948_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4802_ (.A1(_0949_),
    .A2(\reg_file.reg_storage[2][13] ),
    .B(_0761_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4803_ (.A1(_0945_),
    .A2(_0946_),
    .B1(_0947_),
    .B2(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4804_ (.I(_0678_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4805_ (.I(_0675_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4806_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(\reg_file.reg_storage[13][13] ),
    .I2(\reg_file.reg_storage[14][13] ),
    .I3(\reg_file.reg_storage[15][13] ),
    .S0(_0952_),
    .S1(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4807_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(\reg_file.reg_storage[9][13] ),
    .I2(\reg_file.reg_storage[10][13] ),
    .I3(\reg_file.reg_storage[11][13] ),
    .S0(_0952_),
    .S1(_0943_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4808_ (.I(_0803_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4809_ (.I(_0685_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4810_ (.I0(_0944_),
    .I1(_0951_),
    .I2(_0954_),
    .I3(_0955_),
    .S0(_0956_),
    .S1(_0957_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4811_ (.A1(\pc[13] ),
    .A2(_0939_),
    .B1(_0940_),
    .B2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4812_ (.I(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4813_ (.I(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4814_ (.I(_0764_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4815_ (.I(_0596_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4816_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(\reg_file.reg_storage[5][12] ),
    .I2(\reg_file.reg_storage[6][12] ),
    .I3(\reg_file.reg_storage[7][12] ),
    .S0(_0962_),
    .S1(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4817_ (.I(\reg_file.reg_storage[1][12] ),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4818_ (.I(_0739_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(_0966_),
    .A2(\reg_file.reg_storage[3][12] ),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4820_ (.I(_0736_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4821_ (.A1(_0968_),
    .A2(\reg_file.reg_storage[2][12] ),
    .B(_0867_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4822_ (.A1(_0864_),
    .A2(_0965_),
    .B1(_0967_),
    .B2(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4823_ (.I(_0764_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4824_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(\reg_file.reg_storage[13][12] ),
    .I2(\reg_file.reg_storage[14][12] ),
    .I3(\reg_file.reg_storage[15][12] ),
    .S0(_0971_),
    .S1(_0963_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4825_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(\reg_file.reg_storage[9][12] ),
    .I2(\reg_file.reg_storage[10][12] ),
    .I3(\reg_file.reg_storage[11][12] ),
    .S0(_0962_),
    .S1(_0963_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4826_ (.I0(_0964_),
    .I1(_0970_),
    .I2(_0972_),
    .I3(_0973_),
    .S0(_0956_),
    .S1(_0874_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4827_ (.A1(\pc[12] ),
    .A2(_0939_),
    .B1(_0940_),
    .B2(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4828_ (.A1(_0750_),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4829_ (.A1(_0882_),
    .A2(_0961_),
    .B(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4830_ (.I(_0587_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4831_ (.I(_0978_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4832_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(\reg_file.reg_storage[5][11] ),
    .I2(\reg_file.reg_storage[6][11] ),
    .I3(\reg_file.reg_storage[7][11] ),
    .S0(_0942_),
    .S1(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4833_ (.I(\reg_file.reg_storage[1][11] ),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4834_ (.A1(_0966_),
    .A2(\reg_file.reg_storage[3][11] ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4835_ (.A1(_0968_),
    .A2(\reg_file.reg_storage[2][11] ),
    .B(_0761_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4836_ (.A1(_0945_),
    .A2(_0981_),
    .B1(_0982_),
    .B2(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4837_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(\reg_file.reg_storage[13][11] ),
    .I2(\reg_file.reg_storage[14][11] ),
    .I3(\reg_file.reg_storage[15][11] ),
    .S0(_0942_),
    .S1(_0943_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4838_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(\reg_file.reg_storage[9][11] ),
    .I2(\reg_file.reg_storage[10][11] ),
    .I3(\reg_file.reg_storage[11][11] ),
    .S0(_0942_),
    .S1(_0943_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4839_ (.I0(_0980_),
    .I1(_0984_),
    .I2(_0985_),
    .I3(_0986_),
    .S0(_0956_),
    .S1(_0957_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4840_ (.A1(\pc[11] ),
    .A2(_0939_),
    .B1(_0940_),
    .B2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4841_ (.I(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4842_ (.A1(_0725_),
    .A2(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4843_ (.I(_0581_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4844_ (.I(_0592_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4845_ (.I(_0727_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4846_ (.I(_0675_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4847_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(\reg_file.reg_storage[5][10] ),
    .I2(\reg_file.reg_storage[6][10] ),
    .I3(\reg_file.reg_storage[7][10] ),
    .S0(_0993_),
    .S1(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4848_ (.I(_0771_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4849_ (.I(\reg_file.reg_storage[1][10] ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4850_ (.I(_0839_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4851_ (.A1(_0998_),
    .A2(\reg_file.reg_storage[3][10] ),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4852_ (.I(_0730_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4853_ (.A1(_0949_),
    .A2(\reg_file.reg_storage[2][10] ),
    .B(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4854_ (.A1(_0996_),
    .A2(_0997_),
    .B1(_0999_),
    .B2(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4855_ (.I(_0727_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4856_ (.I(_0617_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4857_ (.I(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4858_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(\reg_file.reg_storage[13][10] ),
    .I2(\reg_file.reg_storage[14][10] ),
    .I3(\reg_file.reg_storage[15][10] ),
    .S0(_1003_),
    .S1(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4859_ (.I(_0727_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4860_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(\reg_file.reg_storage[9][10] ),
    .I2(\reg_file.reg_storage[10][10] ),
    .I3(\reg_file.reg_storage[11][10] ),
    .S0(_1007_),
    .S1(_0994_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4861_ (.I(_0613_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4862_ (.I(_0685_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4863_ (.I0(_0995_),
    .I1(_1002_),
    .I2(_1006_),
    .I3(_1008_),
    .S0(_1009_),
    .S1(_1010_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4864_ (.A1(\pc[10] ),
    .A2(_0991_),
    .B1(_0992_),
    .B2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4865_ (.I(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4866_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4867_ (.A1(_0750_),
    .A2(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4868_ (.A1(_0990_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4869_ (.I(_0831_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4870_ (.I0(_0977_),
    .I1(_1016_),
    .S(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4871_ (.A1(_0938_),
    .A2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4872_ (.I(_0588_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4873_ (.I0(\reg_file.reg_storage[4][17] ),
    .I1(\reg_file.reg_storage[5][17] ),
    .I2(\reg_file.reg_storage[6][17] ),
    .I3(\reg_file.reg_storage[7][17] ),
    .S0(_1020_),
    .S1(_0978_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4874_ (.I(\reg_file.reg_storage[1][17] ),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4875_ (.A1(_0756_),
    .A2(\reg_file.reg_storage[3][17] ),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4876_ (.A1(_0948_),
    .A2(\reg_file.reg_storage[2][17] ),
    .B(_0730_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4877_ (.A1(_0771_),
    .A2(_1022_),
    .B1(_1023_),
    .B2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4878_ (.I0(\reg_file.reg_storage[12][17] ),
    .I1(\reg_file.reg_storage[13][17] ),
    .I2(\reg_file.reg_storage[14][17] ),
    .I3(\reg_file.reg_storage[15][17] ),
    .S0(_1020_),
    .S1(_0978_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4879_ (.I0(\reg_file.reg_storage[8][17] ),
    .I1(\reg_file.reg_storage[9][17] ),
    .I2(\reg_file.reg_storage[10][17] ),
    .I3(\reg_file.reg_storage[11][17] ),
    .S0(_1020_),
    .S1(_0978_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4880_ (.I0(_1021_),
    .I1(_1025_),
    .I2(_1026_),
    .I3(_1027_),
    .S0(_0604_),
    .S1(_0605_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4881_ (.A1(\pc[17] ),
    .A2(_0581_),
    .B1(_0592_),
    .B2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4882_ (.A1(_0724_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4883_ (.I(_0749_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4884_ (.I(_0993_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4885_ (.I(_0618_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4886_ (.I(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4887_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(\reg_file.reg_storage[5][16] ),
    .I2(\reg_file.reg_storage[6][16] ),
    .I3(\reg_file.reg_storage[7][16] ),
    .S0(_1032_),
    .S1(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4888_ (.I(\reg_file.reg_storage[1][16] ),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4889_ (.A1(_0817_),
    .A2(\reg_file.reg_storage[3][16] ),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4890_ (.A1(_0797_),
    .A2(\reg_file.reg_storage[2][16] ),
    .B(_0843_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4891_ (.A1(_0792_),
    .A2(_1036_),
    .B1(_1037_),
    .B2(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4892_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(\reg_file.reg_storage[13][16] ),
    .I2(\reg_file.reg_storage[14][16] ),
    .I3(\reg_file.reg_storage[15][16] ),
    .S0(_0966_),
    .S1(_1034_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4893_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(\reg_file.reg_storage[9][16] ),
    .I2(\reg_file.reg_storage[10][16] ),
    .I3(\reg_file.reg_storage[11][16] ),
    .S0(_1032_),
    .S1(_1034_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4894_ (.I0(_1035_),
    .I1(_1039_),
    .I2(_1040_),
    .I3(_1041_),
    .S0(_0805_),
    .S1(_0806_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4895_ (.A1(\pc[16] ),
    .A2(_0788_),
    .B1(_0789_),
    .B2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4896_ (.I(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4897_ (.A1(_1031_),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4898_ (.A1(_1030_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4899_ (.I(_0728_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4900_ (.I0(\reg_file.reg_storage[4][14] ),
    .I1(\reg_file.reg_storage[5][14] ),
    .I2(\reg_file.reg_storage[6][14] ),
    .I3(\reg_file.reg_storage[7][14] ),
    .S0(_0765_),
    .S1(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4901_ (.I(\reg_file.reg_storage[1][14] ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4902_ (.A1(_1032_),
    .A2(\reg_file.reg_storage[3][14] ),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4903_ (.A1(_0968_),
    .A2(\reg_file.reg_storage[2][14] ),
    .B(_0867_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4904_ (.A1(_0864_),
    .A2(_1049_),
    .B1(_1050_),
    .B2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4905_ (.I0(\reg_file.reg_storage[12][14] ),
    .I1(\reg_file.reg_storage[13][14] ),
    .I2(\reg_file.reg_storage[14][14] ),
    .I3(\reg_file.reg_storage[15][14] ),
    .S0(_0962_),
    .S1(_0963_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4906_ (.I0(\reg_file.reg_storage[8][14] ),
    .I1(\reg_file.reg_storage[9][14] ),
    .I2(\reg_file.reg_storage[10][14] ),
    .I3(\reg_file.reg_storage[11][14] ),
    .S0(_0962_),
    .S1(_1047_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4907_ (.I0(_1048_),
    .I1(_1052_),
    .I2(_1053_),
    .I3(_1054_),
    .S0(_0804_),
    .S1(_0874_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4908_ (.A1(\pc[14] ),
    .A2(_0859_),
    .B1(_0860_),
    .B2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4909_ (.I(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4910_ (.I(_1057_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4911_ (.A1(\pc[15] ),
    .A2(_0752_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4912_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(\reg_file.reg_storage[5][15] ),
    .I2(\reg_file.reg_storage[6][15] ),
    .I3(\reg_file.reg_storage[7][15] ),
    .S0(_0775_),
    .S1(_0776_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4913_ (.I(\reg_file.reg_storage[1][15] ),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(_0766_),
    .A2(\reg_file.reg_storage[3][15] ),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4915_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][15] ),
    .B(_0848_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4916_ (.A1(_0843_),
    .A2(_1061_),
    .B1(_1062_),
    .B2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4917_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(\reg_file.reg_storage[13][15] ),
    .I2(\reg_file.reg_storage[14][15] ),
    .I3(\reg_file.reg_storage[15][15] ),
    .S0(_0840_),
    .S1(_0776_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4918_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(\reg_file.reg_storage[9][15] ),
    .I2(\reg_file.reg_storage[10][15] ),
    .I3(\reg_file.reg_storage[11][15] ),
    .S0(_0775_),
    .S1(_0776_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4919_ (.I0(_1060_),
    .I1(_1064_),
    .I2(_1065_),
    .I3(_1066_),
    .S0(_0779_),
    .S1(_0780_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4920_ (.A1(_0754_),
    .A2(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4921_ (.A1(_1059_),
    .A2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4922_ (.I(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4923_ (.A1(_0725_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4924_ (.A1(_0885_),
    .A2(_1058_),
    .B(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4925_ (.I0(_1046_),
    .I1(_1072_),
    .S(_1017_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4926_ (.A1(_0901_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4927_ (.A1(_0936_),
    .A2(_1019_),
    .A3(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4928_ (.A1(_0543_),
    .A2(_0562_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4929_ (.I(_1076_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4930_ (.I(_1077_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4931_ (.I(_0639_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4932_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(\reg_file.reg_storage[5][4] ),
    .I2(\reg_file.reg_storage[6][4] ),
    .I3(\reg_file.reg_storage[7][4] ),
    .S0(_0921_),
    .S1(_1079_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4933_ (.I(_0644_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4934_ (.I0(\reg_file.reg_storage[2][4] ),
    .I1(\reg_file.reg_storage[3][4] ),
    .S(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4935_ (.I0(\reg_file.reg_storage[1][4] ),
    .I1(_1082_),
    .S(_1079_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4936_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(\reg_file.reg_storage[13][4] ),
    .I2(\reg_file.reg_storage[14][4] ),
    .I3(\reg_file.reg_storage[15][4] ),
    .S0(_0906_),
    .S1(_0907_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4937_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(\reg_file.reg_storage[9][4] ),
    .I2(\reg_file.reg_storage[10][4] ),
    .I3(\reg_file.reg_storage[11][4] ),
    .S0(_0921_),
    .S1(_1079_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4938_ (.I(_0573_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4939_ (.I0(_1080_),
    .I1(_1083_),
    .I2(_1084_),
    .I3(_1085_),
    .S0(_0707_),
    .S1(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4940_ (.A1(net3),
    .A2(_0693_),
    .B1(net111),
    .B2(net17),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4941_ (.I(_1088_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4942_ (.A1(_0698_),
    .A2(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4943_ (.A1(_1078_),
    .A2(net99),
    .B(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4944_ (.I(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4945_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4946_ (.A1(_1075_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4947_ (.I(_0617_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4948_ (.I0(\reg_file.reg_storage[4][25] ),
    .I1(\reg_file.reg_storage[5][25] ),
    .I2(\reg_file.reg_storage[6][25] ),
    .I3(\reg_file.reg_storage[7][25] ),
    .S0(_0673_),
    .S1(_1095_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4949_ (.I(\reg_file.reg_storage[1][25] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4950_ (.I(_0630_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4951_ (.I(_1098_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4952_ (.A1(_1099_),
    .A2(\reg_file.reg_storage[3][25] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4953_ (.A1(_0736_),
    .A2(\reg_file.reg_storage[2][25] ),
    .B(_0615_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4954_ (.A1(_0863_),
    .A2(_1097_),
    .B1(_1100_),
    .B2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4955_ (.I0(\reg_file.reg_storage[12][25] ),
    .I1(\reg_file.reg_storage[13][25] ),
    .I2(\reg_file.reg_storage[14][25] ),
    .I3(\reg_file.reg_storage[15][25] ),
    .S0(_1098_),
    .S1(_0596_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4956_ (.I0(\reg_file.reg_storage[8][25] ),
    .I1(\reg_file.reg_storage[9][25] ),
    .I2(\reg_file.reg_storage[10][25] ),
    .I3(\reg_file.reg_storage[11][25] ),
    .S0(_0673_),
    .S1(_1095_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4957_ (.I0(_1096_),
    .I1(_1102_),
    .I2(_1103_),
    .I3(_1104_),
    .S0(_0613_),
    .S1(_0611_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4958_ (.A1(\pc[25] ),
    .A2(_0610_),
    .B1(_0726_),
    .B2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4959_ (.I(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4960_ (.I(_0749_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4961_ (.I0(\reg_file.reg_storage[4][24] ),
    .I1(\reg_file.reg_storage[5][24] ),
    .I2(\reg_file.reg_storage[6][24] ),
    .I3(\reg_file.reg_storage[7][24] ),
    .S0(_0993_),
    .S1(_0953_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4962_ (.I(\reg_file.reg_storage[1][24] ),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4963_ (.A1(_0998_),
    .A2(\reg_file.reg_storage[3][24] ),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4964_ (.A1(_0949_),
    .A2(\reg_file.reg_storage[2][24] ),
    .B(_1000_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4965_ (.A1(_0996_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4966_ (.I0(\reg_file.reg_storage[12][24] ),
    .I1(\reg_file.reg_storage[13][24] ),
    .I2(\reg_file.reg_storage[14][24] ),
    .I3(\reg_file.reg_storage[15][24] ),
    .S0(_1007_),
    .S1(_0994_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4967_ (.I0(\reg_file.reg_storage[8][24] ),
    .I1(\reg_file.reg_storage[9][24] ),
    .I2(\reg_file.reg_storage[10][24] ),
    .I3(\reg_file.reg_storage[11][24] ),
    .S0(_1007_),
    .S1(_0994_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4968_ (.I0(_1109_),
    .I1(_1113_),
    .I2(_1114_),
    .I3(_1115_),
    .S0(_1009_),
    .S1(_0957_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4969_ (.A1(\pc[24] ),
    .A2(_0991_),
    .B1(_0992_),
    .B2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4970_ (.I(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4971_ (.A1(_1108_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4972_ (.A1(_1031_),
    .A2(_1107_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4973_ (.A1(\pc[23] ),
    .A2(_0670_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4974_ (.I(_0629_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4975_ (.I0(\reg_file.reg_storage[12][23] ),
    .I1(\reg_file.reg_storage[13][23] ),
    .I2(\reg_file.reg_storage[14][23] ),
    .I3(\reg_file.reg_storage[15][23] ),
    .S0(_0952_),
    .S1(_0953_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4976_ (.I0(\reg_file.reg_storage[8][23] ),
    .I1(\reg_file.reg_storage[9][23] ),
    .I2(\reg_file.reg_storage[10][23] ),
    .I3(\reg_file.reg_storage[11][23] ),
    .S0(_0952_),
    .S1(_0953_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4977_ (.I0(_1123_),
    .I1(_1124_),
    .S(_0804_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4978_ (.A1(_0757_),
    .A2(\reg_file.reg_storage[3][23] ),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4979_ (.A1(_0797_),
    .A2(\reg_file.reg_storage[2][23] ),
    .B(_1126_),
    .C(_0945_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4980_ (.A1(_0790_),
    .A2(\reg_file.reg_storage[1][23] ),
    .B(_0804_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4981_ (.I0(\reg_file.reg_storage[4][23] ),
    .I1(\reg_file.reg_storage[5][23] ),
    .S(_1007_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4982_ (.A1(_0765_),
    .A2(\reg_file.reg_storage[7][23] ),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4983_ (.I(_0948_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4984_ (.A1(_1131_),
    .A2(\reg_file.reg_storage[6][23] ),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4985_ (.A1(_0871_),
    .A2(_1130_),
    .A3(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4986_ (.A1(_1034_),
    .A2(_1129_),
    .B(_1133_),
    .C(net9),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4987_ (.A1(_1127_),
    .A2(_1128_),
    .B(_1134_),
    .C(_1122_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4988_ (.A1(_1122_),
    .A2(_1125_),
    .B(_1135_),
    .C(_0753_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4989_ (.A1(_1121_),
    .A2(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4990_ (.A1(_0724_),
    .A2(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4991_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(\reg_file.reg_storage[5][22] ),
    .I2(\reg_file.reg_storage[6][22] ),
    .I3(\reg_file.reg_storage[7][22] ),
    .S0(_0941_),
    .S1(_1033_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4992_ (.I(\reg_file.reg_storage[1][22] ),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4993_ (.A1(_0993_),
    .A2(\reg_file.reg_storage[3][22] ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4994_ (.A1(_0768_),
    .A2(\reg_file.reg_storage[2][22] ),
    .B(_0847_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4995_ (.A1(_1000_),
    .A2(_1140_),
    .B1(_1141_),
    .B2(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4996_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(\reg_file.reg_storage[13][22] ),
    .I2(\reg_file.reg_storage[14][22] ),
    .I3(\reg_file.reg_storage[15][22] ),
    .S0(_0941_),
    .S1(_0758_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4997_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(\reg_file.reg_storage[9][22] ),
    .I2(\reg_file.reg_storage[10][22] ),
    .I3(\reg_file.reg_storage[11][22] ),
    .S0(_0941_),
    .S1(_0758_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4998_ (.I0(_1139_),
    .I1(_1143_),
    .I2(_1144_),
    .I3(_1145_),
    .S0(_0803_),
    .S1(_0686_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4999_ (.A1(\pc[22] ),
    .A2(_0751_),
    .B1(_0753_),
    .B2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5000_ (.I(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5001_ (.A1(_1108_),
    .A2(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5002_ (.A1(_1138_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5003_ (.I(_0830_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5004_ (.I(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5005_ (.I0(_1120_),
    .I1(_1150_),
    .S(_1152_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5006_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(\reg_file.reg_storage[5][21] ),
    .I2(\reg_file.reg_storage[6][21] ),
    .I3(\reg_file.reg_storage[7][21] ),
    .S0(_1020_),
    .S1(_1004_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5007_ (.I(\reg_file.reg_storage[1][21] ),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5008_ (.A1(_0678_),
    .A2(\reg_file.reg_storage[3][21] ),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5009_ (.A1(_0948_),
    .A2(\reg_file.reg_storage[2][21] ),
    .B(_0770_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5010_ (.A1(_0847_),
    .A2(_1155_),
    .B1(_1156_),
    .B2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5011_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(\reg_file.reg_storage[13][21] ),
    .I2(\reg_file.reg_storage[14][21] ),
    .I3(\reg_file.reg_storage[15][21] ),
    .S0(_0755_),
    .S1(_0618_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5012_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(\reg_file.reg_storage[9][21] ),
    .I2(\reg_file.reg_storage[10][21] ),
    .I3(\reg_file.reg_storage[11][21] ),
    .S0(_0755_),
    .S1(_1004_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5013_ (.I0(_1154_),
    .I1(_1158_),
    .I2(_1159_),
    .I3(_1160_),
    .S0(_0612_),
    .S1(_0685_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5014_ (.A1(\pc[21] ),
    .A2(_0609_),
    .B1(_0671_),
    .B2(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5015_ (.A1(_0724_),
    .A2(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5016_ (.A1(\pc[20] ),
    .A2(_0991_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5017_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(\reg_file.reg_storage[5][20] ),
    .I2(\reg_file.reg_storage[6][20] ),
    .I3(\reg_file.reg_storage[7][20] ),
    .S0(_1003_),
    .S1(_1005_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5018_ (.I(\reg_file.reg_storage[1][20] ),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5019_ (.A1(_0998_),
    .A2(\reg_file.reg_storage[3][20] ),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5020_ (.A1(_0949_),
    .A2(\reg_file.reg_storage[2][20] ),
    .B(_1000_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5021_ (.A1(_0996_),
    .A2(_1166_),
    .B1(_1167_),
    .B2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5022_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(\reg_file.reg_storage[13][20] ),
    .I2(\reg_file.reg_storage[14][20] ),
    .I3(\reg_file.reg_storage[15][20] ),
    .S0(_1003_),
    .S1(_1005_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5023_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(\reg_file.reg_storage[9][20] ),
    .I2(\reg_file.reg_storage[10][20] ),
    .I3(\reg_file.reg_storage[11][20] ),
    .S0(_1003_),
    .S1(_1005_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5024_ (.I0(_1165_),
    .I1(_1169_),
    .I2(_1170_),
    .I3(_1171_),
    .S0(_1009_),
    .S1(_1010_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5025_ (.A1(_0992_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5026_ (.A1(_1164_),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5027_ (.I(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5028_ (.I(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5029_ (.A1(_1108_),
    .A2(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5030_ (.A1(_1163_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5031_ (.I(_0578_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5032_ (.I(_0739_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5033_ (.I(_1004_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5034_ (.I0(\reg_file.reg_storage[4][19] ),
    .I1(\reg_file.reg_storage[5][19] ),
    .I2(\reg_file.reg_storage[6][19] ),
    .I3(\reg_file.reg_storage[7][19] ),
    .S0(_1180_),
    .S1(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5035_ (.I(\reg_file.reg_storage[1][19] ),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5036_ (.A1(_0998_),
    .A2(\reg_file.reg_storage[3][19] ),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5037_ (.A1(_1131_),
    .A2(\reg_file.reg_storage[2][19] ),
    .B(_0731_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5038_ (.A1(_0996_),
    .A2(_1183_),
    .B1(_1184_),
    .B2(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5039_ (.I0(\reg_file.reg_storage[12][19] ),
    .I1(\reg_file.reg_storage[13][19] ),
    .I2(\reg_file.reg_storage[14][19] ),
    .I3(\reg_file.reg_storage[15][19] ),
    .S0(_1180_),
    .S1(_1181_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5040_ (.I0(\reg_file.reg_storage[8][19] ),
    .I1(\reg_file.reg_storage[9][19] ),
    .I2(\reg_file.reg_storage[10][19] ),
    .I3(\reg_file.reg_storage[11][19] ),
    .S0(_1180_),
    .S1(_1181_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5041_ (.I0(_1182_),
    .I1(_1186_),
    .I2(_1187_),
    .I3(_1188_),
    .S0(_1009_),
    .S1(_1010_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5042_ (.A1(\pc[19] ),
    .A2(_0991_),
    .B1(_0992_),
    .B2(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5043_ (.I(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5044_ (.A1(_1179_),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5045_ (.I0(\reg_file.reg_storage[4][18] ),
    .I1(\reg_file.reg_storage[5][18] ),
    .I2(\reg_file.reg_storage[6][18] ),
    .I3(\reg_file.reg_storage[7][18] ),
    .S0(_0673_),
    .S1(_1095_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5046_ (.I(\reg_file.reg_storage[1][18] ),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5047_ (.A1(_0756_),
    .A2(\reg_file.reg_storage[3][18] ),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5048_ (.A1(_0736_),
    .A2(\reg_file.reg_storage[2][18] ),
    .B(_0615_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5049_ (.A1(_0863_),
    .A2(_1194_),
    .B1(_1195_),
    .B2(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5050_ (.I0(\reg_file.reg_storage[12][18] ),
    .I1(\reg_file.reg_storage[13][18] ),
    .I2(\reg_file.reg_storage[14][18] ),
    .I3(\reg_file.reg_storage[15][18] ),
    .S0(_1098_),
    .S1(_0596_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5051_ (.I0(\reg_file.reg_storage[8][18] ),
    .I1(\reg_file.reg_storage[9][18] ),
    .I2(\reg_file.reg_storage[10][18] ),
    .I3(\reg_file.reg_storage[11][18] ),
    .S0(_1098_),
    .S1(_1095_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5052_ (.I0(_1193_),
    .I1(_1197_),
    .I2(_1198_),
    .I3(_1199_),
    .S0(_0604_),
    .S1(_0605_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5053_ (.A1(\pc[18] ),
    .A2(_0581_),
    .B1(_0592_),
    .B2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5054_ (.A1(_1031_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5055_ (.A1(_1192_),
    .A2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5056_ (.I0(_1178_),
    .I1(_1203_),
    .S(_1152_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5057_ (.I(_0937_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5058_ (.I0(_1153_),
    .I1(_1204_),
    .S(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5059_ (.I(_0933_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5060_ (.I(_1151_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5061_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(\reg_file.reg_storage[5][29] ),
    .I2(\reg_file.reg_storage[6][29] ),
    .I3(\reg_file.reg_storage[7][29] ),
    .S0(_0971_),
    .S1(_0979_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5062_ (.I(\reg_file.reg_storage[1][29] ),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5063_ (.A1(_0966_),
    .A2(\reg_file.reg_storage[3][29] ),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5064_ (.A1(_0968_),
    .A2(\reg_file.reg_storage[2][29] ),
    .B(_0761_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5065_ (.A1(_0945_),
    .A2(_1210_),
    .B1(_1211_),
    .B2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5066_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(\reg_file.reg_storage[13][29] ),
    .I2(\reg_file.reg_storage[14][29] ),
    .I3(\reg_file.reg_storage[15][29] ),
    .S0(_0971_),
    .S1(_0979_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5067_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(\reg_file.reg_storage[9][29] ),
    .I2(\reg_file.reg_storage[10][29] ),
    .I3(\reg_file.reg_storage[11][29] ),
    .S0(_0971_),
    .S1(_0979_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5068_ (.I0(_1209_),
    .I1(_1213_),
    .I2(_1214_),
    .I3(_1215_),
    .S0(_0956_),
    .S1(_0957_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5069_ (.A1(\pc[29] ),
    .A2(_0939_),
    .B1(_0940_),
    .B2(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5070_ (.I(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5071_ (.A1(_1031_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5072_ (.A1(\pc[28] ),
    .A2(_0788_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5073_ (.I0(\reg_file.reg_storage[12][28] ),
    .I1(\reg_file.reg_storage[13][28] ),
    .I2(\reg_file.reg_storage[14][28] ),
    .I3(\reg_file.reg_storage[15][28] ),
    .S0(_0794_),
    .S1(_0814_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5074_ (.I0(\reg_file.reg_storage[8][28] ),
    .I1(\reg_file.reg_storage[9][28] ),
    .I2(\reg_file.reg_storage[10][28] ),
    .I3(\reg_file.reg_storage[11][28] ),
    .S0(_0794_),
    .S1(_0814_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5075_ (.I0(_1221_),
    .I1(_1222_),
    .S(_0779_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5076_ (.I0(\reg_file.reg_storage[4][28] ),
    .I1(\reg_file.reg_storage[5][28] ),
    .I2(\reg_file.reg_storage[6][28] ),
    .I3(\reg_file.reg_storage[7][28] ),
    .S0(_0813_),
    .S1(_0814_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5077_ (.A1(_0805_),
    .A2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5078_ (.I(_1047_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5079_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][28] ),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5080_ (.A1(_0817_),
    .A2(\reg_file.reg_storage[3][28] ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5081_ (.A1(_1226_),
    .A2(_1227_),
    .A3(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5082_ (.I(\reg_file.reg_storage[1][28] ),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5083_ (.A1(_0762_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5084_ (.A1(_1229_),
    .A2(_1231_),
    .B(net9),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5085_ (.A1(_1225_),
    .A2(_1232_),
    .B(_1122_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _5086_ (.A1(_1122_),
    .A2(_1223_),
    .B(_1233_),
    .C(_0754_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5087_ (.A1(_1220_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5088_ (.A1(_1179_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5089_ (.A1(_1219_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5090_ (.I0(\reg_file.reg_storage[4][27] ),
    .I1(\reg_file.reg_storage[5][27] ),
    .I2(\reg_file.reg_storage[6][27] ),
    .I3(\reg_file.reg_storage[7][27] ),
    .S0(_1099_),
    .S1(_0680_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5091_ (.I(\reg_file.reg_storage[1][27] ),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5092_ (.A1(_0775_),
    .A2(\reg_file.reg_storage[3][27] ),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5093_ (.A1(_1131_),
    .A2(\reg_file.reg_storage[2][27] ),
    .B(_0863_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5094_ (.A1(_0848_),
    .A2(_1239_),
    .B1(_1240_),
    .B2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5095_ (.I0(\reg_file.reg_storage[12][27] ),
    .I1(\reg_file.reg_storage[13][27] ),
    .I2(\reg_file.reg_storage[14][27] ),
    .I3(\reg_file.reg_storage[15][27] ),
    .S0(_1099_),
    .S1(_1033_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5096_ (.I0(\reg_file.reg_storage[8][27] ),
    .I1(\reg_file.reg_storage[9][27] ),
    .I2(\reg_file.reg_storage[10][27] ),
    .I3(\reg_file.reg_storage[11][27] ),
    .S0(_1099_),
    .S1(_1033_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5097_ (.I0(_1238_),
    .I1(_1242_),
    .I2(_1243_),
    .I3(_1244_),
    .S0(_0684_),
    .S1(_0686_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5098_ (.A1(\pc[27] ),
    .A2(_0670_),
    .B1(_0672_),
    .B2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5099_ (.I(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5100_ (.I0(\reg_file.reg_storage[4][26] ),
    .I1(\reg_file.reg_storage[5][26] ),
    .I2(\reg_file.reg_storage[6][26] ),
    .I3(\reg_file.reg_storage[7][26] ),
    .S0(_1180_),
    .S1(_1181_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5101_ (.I(\reg_file.reg_storage[1][26] ),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5102_ (.A1(_0813_),
    .A2(\reg_file.reg_storage[3][26] ),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5103_ (.A1(_1131_),
    .A2(\reg_file.reg_storage[2][26] ),
    .B(_0731_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5104_ (.A1(_0772_),
    .A2(_1249_),
    .B1(_1250_),
    .B2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5105_ (.I0(\reg_file.reg_storage[12][26] ),
    .I1(\reg_file.reg_storage[13][26] ),
    .I2(\reg_file.reg_storage[14][26] ),
    .I3(\reg_file.reg_storage[15][26] ),
    .S0(_0733_),
    .S1(_0676_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5106_ (.I0(\reg_file.reg_storage[8][26] ),
    .I1(\reg_file.reg_storage[9][26] ),
    .I2(\reg_file.reg_storage[10][26] ),
    .I3(\reg_file.reg_storage[11][26] ),
    .S0(_0733_),
    .S1(_0676_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5107_ (.I0(_1248_),
    .I1(_1252_),
    .I2(_1253_),
    .I3(_1254_),
    .S0(_0684_),
    .S1(_1010_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5108_ (.A1(\pc[26] ),
    .A2(_0670_),
    .B1(_0672_),
    .B2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5109_ (.A1(_1108_),
    .A2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5110_ (.A1(_0811_),
    .A2(_1247_),
    .B(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5111_ (.A1(_1152_),
    .A2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5112_ (.A1(_1208_),
    .A2(_1237_),
    .B(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5113_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(\reg_file.reg_storage[5][30] ),
    .I2(\reg_file.reg_storage[6][30] ),
    .I3(\reg_file.reg_storage[7][30] ),
    .S0(_0870_),
    .S1(_0861_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5114_ (.I(\reg_file.reg_storage[1][30] ),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5115_ (.A1(_1032_),
    .A2(\reg_file.reg_storage[3][30] ),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5116_ (.A1(_0846_),
    .A2(\reg_file.reg_storage[2][30] ),
    .B(_0867_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5117_ (.A1(_0864_),
    .A2(_1262_),
    .B1(_1263_),
    .B2(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5118_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(\reg_file.reg_storage[13][30] ),
    .I2(\reg_file.reg_storage[14][30] ),
    .I3(\reg_file.reg_storage[15][30] ),
    .S0(_0765_),
    .S1(_1047_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5119_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(\reg_file.reg_storage[9][30] ),
    .I2(\reg_file.reg_storage[10][30] ),
    .I3(\reg_file.reg_storage[11][30] ),
    .S0(_0870_),
    .S1(_0871_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5120_ (.I0(_1261_),
    .I1(_1265_),
    .I2(_1266_),
    .I3(_1267_),
    .S0(_0854_),
    .S1(_0874_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5121_ (.A1(\pc[30] ),
    .A2(_0859_),
    .B1(_0860_),
    .B2(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5122_ (.I(_1269_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5123_ (.A1(_1179_),
    .A2(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5124_ (.I0(\reg_file.reg_storage[4][31] ),
    .I1(\reg_file.reg_storage[5][31] ),
    .I2(\reg_file.reg_storage[6][31] ),
    .I3(\reg_file.reg_storage[7][31] ),
    .S0(_0795_),
    .S1(_1226_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5125_ (.I(\reg_file.reg_storage[1][31] ),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_0795_),
    .A2(\reg_file.reg_storage[3][31] ),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5127_ (.A1(_0797_),
    .A2(\reg_file.reg_storage[2][31] ),
    .B(_0792_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5128_ (.A1(_0792_),
    .A2(_1273_),
    .B1(_1274_),
    .B2(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5129_ (.I0(\reg_file.reg_storage[12][31] ),
    .I1(\reg_file.reg_storage[13][31] ),
    .I2(\reg_file.reg_storage[14][31] ),
    .I3(\reg_file.reg_storage[15][31] ),
    .S0(_0817_),
    .S1(_1226_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5130_ (.I0(\reg_file.reg_storage[8][31] ),
    .I1(\reg_file.reg_storage[9][31] ),
    .I2(\reg_file.reg_storage[10][31] ),
    .I3(\reg_file.reg_storage[11][31] ),
    .S0(_0795_),
    .S1(_1226_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5131_ (.I0(_1272_),
    .I1(_1276_),
    .I2(_1277_),
    .I3(_1278_),
    .S0(_0805_),
    .S1(_0806_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5132_ (.A1(\pc[31] ),
    .A2(_0788_),
    .B1(_0789_),
    .B2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5133_ (.A1(_1179_),
    .A2(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5134_ (.A1(_0837_),
    .A2(_1271_),
    .A3(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5135_ (.A1(_0900_),
    .A2(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5136_ (.A1(_0722_),
    .A2(_1260_),
    .B(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(_1207_),
    .A2(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5138_ (.A1(_0936_),
    .A2(_1206_),
    .B(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5139_ (.I(_0532_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5140_ (.A1(_0536_),
    .A2(_0525_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5141_ (.A1(_1287_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5142_ (.A1(_0935_),
    .A2(_1094_),
    .B1(_1286_),
    .B2(_1093_),
    .C(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5143_ (.I(_0536_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5144_ (.I(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5145_ (.I(_0669_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5146_ (.A1(_1293_),
    .A2(_0626_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5147_ (.A1(_0672_),
    .A2(_0687_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5148_ (.A1(_1294_),
    .A2(_1295_),
    .B1(_0696_),
    .B2(_0710_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(_1292_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5150_ (.I(net24),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5151_ (.A1(_1298_),
    .A2(_1287_),
    .A3(_0537_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5152_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5153_ (.A1(_0688_),
    .A2(_0717_),
    .A3(net115),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5154_ (.A1(_1297_),
    .A2(_1300_),
    .A3(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5155_ (.I(_0933_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5156_ (.I(_1092_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5157_ (.A1(_0531_),
    .A2(_0507_),
    .A3(_1288_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5158_ (.A1(_1304_),
    .A2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5159_ (.A1(_1303_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5160_ (.I(_0937_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5161_ (.I(_1208_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5162_ (.A1(_0636_),
    .A2(_0885_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5163_ (.A1(_0884_),
    .A2(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5164_ (.A1(_0555_),
    .A2(_0575_),
    .A3(_0607_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5165_ (.I(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5166_ (.A1(_0833_),
    .A2(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5167_ (.A1(_1309_),
    .A2(_1311_),
    .B(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5168_ (.A1(_1308_),
    .A2(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5169_ (.A1(_1296_),
    .A2(_1301_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5170_ (.A1(_1298_),
    .A2(_1287_),
    .A3(_0526_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5171_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5172_ (.A1(_1307_),
    .A2(_1316_),
    .B1(_1317_),
    .B2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5173_ (.A1(_0716_),
    .A2(_1290_),
    .A3(_1302_),
    .A4(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5174_ (.A1(_0540_),
    .A2(_0715_),
    .B(_1321_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5175_ (.I(_1322_),
    .ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5176_ (.A1(_0528_),
    .A2(_0534_),
    .A3(_0538_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5177_ (.I(_1323_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5178_ (.I(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5179_ (.A1(_0883_),
    .A2(_0713_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5180_ (.A1(_0668_),
    .A2(_0714_),
    .B(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5181_ (.I(_0691_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5182_ (.I(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5183_ (.A1(_0929_),
    .A2(_0930_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5184_ (.I(_0928_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5185_ (.I(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5186_ (.I(_1332_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5187_ (.A1(_0909_),
    .A2(_0917_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5188_ (.I(_1331_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5189_ (.A1(_1335_),
    .A2(_0923_),
    .A3(_0926_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5190_ (.A1(_1333_),
    .A2(_1334_),
    .B(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5191_ (.I(_1077_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5192_ (.A1(_1329_),
    .A2(_1330_),
    .B1(_1337_),
    .B2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5193_ (.A1(_0828_),
    .A2(_0748_),
    .A3(_0711_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5194_ (.A1(_0662_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5195_ (.A1(_1339_),
    .A2(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5196_ (.A1(_0895_),
    .A2(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5197_ (.A1(_0895_),
    .A2(_1342_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5198_ (.I(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5199_ (.A1(_1343_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5200_ (.A1(_1327_),
    .A2(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5201_ (.I(_1304_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5202_ (.I(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5203_ (.I(_1207_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5204_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5205_ (.I(_1152_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5206_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5207_ (.I(_0885_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5208_ (.I(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5209_ (.I(_1106_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5210_ (.I(_0786_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5211_ (.I(_1357_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5212_ (.I(_1256_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5213_ (.I(_1359_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5214_ (.A1(_1358_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5215_ (.A1(_1355_),
    .A2(_1356_),
    .B(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5216_ (.A1(_1121_),
    .A2(_1136_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5217_ (.I(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5218_ (.I(_1357_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5219_ (.A1(_1365_),
    .A2(_1118_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5220_ (.A1(_1358_),
    .A2(_1364_),
    .B(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5221_ (.A1(_0833_),
    .A2(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5222_ (.A1(_1353_),
    .A2(_1362_),
    .B(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5223_ (.A1(_1365_),
    .A2(_1148_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5224_ (.I(_0750_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5225_ (.I(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5226_ (.I(_1162_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5227_ (.A1(_1372_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5228_ (.A1(_1370_),
    .A2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5229_ (.I(_1357_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5230_ (.A1(_1376_),
    .A2(_1176_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5231_ (.I(_0882_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5232_ (.A1(_1378_),
    .A2(_1191_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5233_ (.A1(_1377_),
    .A2(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5234_ (.I(_1017_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5235_ (.I0(_1375_),
    .I1(_1380_),
    .S(_1381_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5236_ (.I0(_1369_),
    .I1(_1382_),
    .S(_1308_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5237_ (.I(_0934_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5238_ (.I(_0900_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5239_ (.I(_0836_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5240_ (.I(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5241_ (.I(_1270_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5242_ (.A1(_1358_),
    .A2(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5243_ (.A1(_1355_),
    .A2(_1217_),
    .B(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5244_ (.A1(_1220_),
    .A2(_1234_),
    .B(_1372_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5245_ (.I(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5246_ (.I(_1247_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5247_ (.A1(_1372_),
    .A2(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5248_ (.A1(_1392_),
    .A2(_1394_),
    .B(_1386_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5249_ (.A1(_1387_),
    .A2(_1390_),
    .B(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5250_ (.I(_0721_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5251_ (.I(_1280_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5252_ (.A1(_1358_),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5253_ (.A1(_1397_),
    .A2(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5254_ (.I(_0837_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5255_ (.I(_1401_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5256_ (.A1(_1385_),
    .A2(_1396_),
    .B1(_1400_),
    .B2(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5257_ (.A1(_1384_),
    .A2(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5258_ (.A1(_1351_),
    .A2(_1383_),
    .B(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5259_ (.I(_1339_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5260_ (.I(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5261_ (.I(_1407_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5262_ (.I(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5263_ (.A1(_1357_),
    .A2(_0975_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5264_ (.I(_1371_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5265_ (.A1(_1411_),
    .A2(_0989_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(_1410_),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5267_ (.I(_1354_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5268_ (.I(_0961_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5269_ (.I(_0725_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5270_ (.I(_1056_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5271_ (.A1(_1416_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5272_ (.A1(_1414_),
    .A2(_1415_),
    .B(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5273_ (.I0(_1413_),
    .I1(_1419_),
    .S(_0838_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_1416_),
    .A2(_1201_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5275_ (.A1(_1371_),
    .A2(_1029_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5276_ (.A1(_1421_),
    .A2(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5277_ (.A1(_1416_),
    .A2(_1044_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(_1378_),
    .A2(_1070_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5279_ (.A1(_1424_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5280_ (.I0(_1423_),
    .I1(_1426_),
    .S(_1381_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5281_ (.I0(_1420_),
    .I1(_1427_),
    .S(_1385_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5282_ (.I(_1408_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5283_ (.I(_0938_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5284_ (.A1(_1411_),
    .A2(_0746_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5285_ (.A1(_1376_),
    .A2(_1014_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5286_ (.A1(_1431_),
    .A2(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5287_ (.A1(_1372_),
    .A2(_0809_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5288_ (.A1(_1376_),
    .A2(_0783_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5289_ (.A1(_1434_),
    .A2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5290_ (.I0(_1433_),
    .I1(_1436_),
    .S(_1353_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5291_ (.I(_1386_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5292_ (.A1(_1378_),
    .A2(_0896_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5293_ (.I(_0877_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5294_ (.A1(_1354_),
    .A2(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5295_ (.A1(_1439_),
    .A2(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(_1371_),
    .A2(_0857_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5297_ (.A1(_1376_),
    .A2(_0825_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5298_ (.A1(_1443_),
    .A2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_0838_),
    .A2(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5300_ (.I(_1205_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5301_ (.A1(_1438_),
    .A2(_1442_),
    .B(_1446_),
    .C(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5302_ (.A1(_1430_),
    .A2(_1437_),
    .B(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5303_ (.A1(_1429_),
    .A2(_1449_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5304_ (.I(_1304_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5305_ (.A1(_1409_),
    .A2(_1428_),
    .B(_1450_),
    .C(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5306_ (.A1(_1349_),
    .A2(_1405_),
    .B(_1452_),
    .C(_1289_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5307_ (.I(_1384_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5308_ (.I(_0896_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5309_ (.I(_1300_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5310_ (.I(_1291_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5311_ (.A1(_1409_),
    .A2(_0896_),
    .B(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5312_ (.A1(_1454_),
    .A2(_1455_),
    .B(_1456_),
    .C(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5313_ (.I(_1307_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5314_ (.I(_0722_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5315_ (.I(_0608_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5316_ (.A1(_0666_),
    .A2(_1365_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5317_ (.A1(_1462_),
    .A2(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5318_ (.A1(_1416_),
    .A2(_0883_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(_1439_),
    .A2(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5320_ (.I(_1017_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5321_ (.I0(_1464_),
    .I1(_1466_),
    .S(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5322_ (.A1(_1461_),
    .A2(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5323_ (.A1(_1339_),
    .A2(_0894_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5324_ (.I(_1319_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5325_ (.A1(_1460_),
    .A2(_1469_),
    .B1(_1470_),
    .B2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5326_ (.A1(_1453_),
    .A2(_1459_),
    .A3(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5327_ (.A1(_1325_),
    .A2(_1347_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5328_ (.I(_1474_),
    .ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5329_ (.A1(_1327_),
    .A2(_1344_),
    .B(_1343_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _5330_ (.A1(_0653_),
    .A2(_0576_),
    .A3(_0719_),
    .A4(_0932_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5331_ (.I(_1476_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5332_ (.A1(_0659_),
    .A2(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5333_ (.A1(_1091_),
    .A2(_1478_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5334_ (.A1(_0877_),
    .A2(_1479_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5335_ (.I(_0716_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5336_ (.A1(_1475_),
    .A2(_1480_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5337_ (.A1(_1481_),
    .A2(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5338_ (.A1(_1475_),
    .A2(_1480_),
    .B(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5339_ (.I(_1451_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5340_ (.I(_0936_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5341_ (.I0(_1150_),
    .I1(_1178_),
    .S(_0829_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5342_ (.I0(_1258_),
    .I1(_1120_),
    .S(_0829_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5343_ (.I0(_1487_),
    .I1(_1488_),
    .S(_0901_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5344_ (.A1(_1271_),
    .A2(_1281_),
    .B(_0835_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5345_ (.A1(_0835_),
    .A2(_1237_),
    .B(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5346_ (.A1(_1397_),
    .A2(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(_1350_),
    .A2(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5348_ (.A1(_1486_),
    .A2(_1489_),
    .B(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5349_ (.I(_1429_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5350_ (.I0(_1046_),
    .I1(_1203_),
    .S(_0835_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5351_ (.I0(_1072_),
    .I1(_0977_),
    .S(_0830_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5352_ (.I(_1205_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5353_ (.I0(_1496_),
    .I1(_1497_),
    .S(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5354_ (.I(_1461_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5355_ (.I0(_1016_),
    .I1(_0785_),
    .S(_1151_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5356_ (.A1(_1500_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5357_ (.I(_0711_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5358_ (.I(_1503_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5359_ (.I(_1504_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5360_ (.A1(_0836_),
    .A2(_0827_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5361_ (.A1(_0836_),
    .A2(_0880_),
    .B(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5362_ (.A1(_1505_),
    .A2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5363_ (.A1(_1409_),
    .A2(_1502_),
    .A3(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5364_ (.I(_1348_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5365_ (.A1(_1495_),
    .A2(_1499_),
    .B(_1509_),
    .C(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5366_ (.I(_1289_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5367_ (.A1(_1485_),
    .A2(_1494_),
    .B(_1511_),
    .C(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5368_ (.I(_1299_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5369_ (.I(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5370_ (.I(_1515_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5371_ (.I(_1348_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5372_ (.I(_1457_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5373_ (.A1(_1440_),
    .A2(_1517_),
    .B(_1518_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5374_ (.A1(_1440_),
    .A2(_1485_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5375_ (.A1(_1516_),
    .A2(_1519_),
    .A3(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5376_ (.I(_0722_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5377_ (.I(_1311_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5378_ (.A1(_0878_),
    .A2(_0897_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5379_ (.A1(_1309_),
    .A2(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5380_ (.A1(_1309_),
    .A2(_1523_),
    .B(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5381_ (.A1(_0831_),
    .A2(_1313_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5382_ (.A1(_1385_),
    .A2(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5383_ (.A1(_1522_),
    .A2(_1526_),
    .B(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5384_ (.A1(_0876_),
    .A2(_1091_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5385_ (.I(_1319_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5386_ (.I(_1531_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5387_ (.A1(_1460_),
    .A2(_1529_),
    .B1(_1530_),
    .B2(_1532_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5388_ (.A1(_1484_),
    .A2(_1513_),
    .A3(_1521_),
    .A4(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5389_ (.I(_1534_),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5390_ (.I(_0856_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5391_ (.I(_0637_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5392_ (.A1(_0491_),
    .A2(_0502_),
    .A3(_0500_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5393_ (.I(_1537_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5394_ (.A1(net18),
    .A2(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5395_ (.I(_0645_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5396_ (.I(_0570_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5397_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(\reg_file.reg_storage[5][5] ),
    .I2(\reg_file.reg_storage[6][5] ),
    .I3(\reg_file.reg_storage[7][5] ),
    .S0(_1540_),
    .S1(_1541_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5398_ (.I(_0644_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5399_ (.I0(\reg_file.reg_storage[2][5] ),
    .I1(\reg_file.reg_storage[3][5] ),
    .S(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5400_ (.I0(\reg_file.reg_storage[1][5] ),
    .I1(_1544_),
    .S(_1541_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5401_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(\reg_file.reg_storage[13][5] ),
    .I2(\reg_file.reg_storage[14][5] ),
    .I3(\reg_file.reg_storage[15][5] ),
    .S0(_1540_),
    .S1(_1541_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5402_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(\reg_file.reg_storage[9][5] ),
    .I2(\reg_file.reg_storage[10][5] ),
    .I3(\reg_file.reg_storage[11][5] ),
    .S0(_1540_),
    .S1(_1541_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5403_ (.I0(_1542_),
    .I1(_1545_),
    .I2(_1546_),
    .I3(_1547_),
    .S0(_0904_),
    .S1(_1086_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5404_ (.I(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5405_ (.I(_0903_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5406_ (.A1(_1536_),
    .A2(_1539_),
    .B1(_1549_),
    .B2(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5407_ (.I(_1551_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5408_ (.A1(_0653_),
    .A2(_0576_),
    .A3(_0719_),
    .A4(_0932_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5409_ (.A1(_0527_),
    .A2(_0506_),
    .A3(_0526_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5410_ (.A1(_1091_),
    .A2(net97),
    .B(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5411_ (.A1(_1552_),
    .A2(_1555_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5412_ (.A1(_1535_),
    .A2(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5413_ (.A1(_1440_),
    .A2(_1479_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5414_ (.A1(_1558_),
    .A2(_1482_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5415_ (.A1(_1557_),
    .A2(_1559_),
    .B(_1481_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5416_ (.A1(_1557_),
    .A2(_1559_),
    .B(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5417_ (.I(_1093_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5418_ (.I(_1562_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5419_ (.I(_1208_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5420_ (.I0(_1399_),
    .I1(_1390_),
    .S(_1564_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5421_ (.A1(_1498_),
    .A2(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5422_ (.A1(_1392_),
    .A2(_1394_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5423_ (.I0(_1567_),
    .I1(_1362_),
    .S(_1564_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5424_ (.I0(_1367_),
    .I1(_1375_),
    .S(_1564_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5425_ (.A1(_1308_),
    .A2(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5426_ (.A1(_1498_),
    .A2(_1568_),
    .B(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5427_ (.I(_1408_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5428_ (.I0(_1566_),
    .I1(_1571_),
    .S(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5429_ (.I(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5430_ (.I(_0934_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5431_ (.I(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5432_ (.I(_1386_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5433_ (.I0(_1445_),
    .I1(_1436_),
    .S(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5434_ (.I0(_1433_),
    .I1(_1413_),
    .S(_0881_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5435_ (.I0(_1578_),
    .I1(_1579_),
    .S(_1522_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5436_ (.I0(_1423_),
    .I1(_1380_),
    .S(_0881_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5437_ (.A1(_1500_),
    .A2(_1581_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5438_ (.I(_0938_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5439_ (.I0(_1419_),
    .I1(_1426_),
    .S(_0881_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5440_ (.A1(_1583_),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5441_ (.A1(_1351_),
    .A2(_1582_),
    .A3(_1585_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5442_ (.A1(_1576_),
    .A2(_1580_),
    .B(_1586_),
    .C(_1349_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5443_ (.A1(_1563_),
    .A2(_1574_),
    .B(_1587_),
    .C(_1512_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5444_ (.A1(_1401_),
    .A2(_1464_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5445_ (.A1(_1441_),
    .A2(_1443_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5446_ (.I0(_1466_),
    .I1(_1590_),
    .S(_0832_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5447_ (.A1(_0938_),
    .A2(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5448_ (.A1(_1447_),
    .A2(_1589_),
    .B(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5449_ (.I(_1593_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5450_ (.I(_1552_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5451_ (.A1(_1535_),
    .A2(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5452_ (.I(_1531_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(_1535_),
    .A2(_1595_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5454_ (.I(_1514_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5455_ (.A1(_1535_),
    .A2(_1595_),
    .B(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5456_ (.A1(_1518_),
    .A2(_1598_),
    .B(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5457_ (.A1(_1460_),
    .A2(_1594_),
    .B1(_1596_),
    .B2(_1597_),
    .C(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5458_ (.A1(_1561_),
    .A2(_1588_),
    .A3(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5459_ (.I(_1603_),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5460_ (.A1(_1430_),
    .A2(_1073_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5461_ (.A1(_1500_),
    .A2(_1204_),
    .B(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5462_ (.I(_0723_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5463_ (.A1(_1505_),
    .A2(_0834_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5464_ (.I(_1207_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5465_ (.I(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5466_ (.A1(_1606_),
    .A2(_1018_),
    .B(_1607_),
    .C(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5467_ (.I(_1087_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5468_ (.A1(_1536_),
    .A2(_1088_),
    .B1(_1611_),
    .B2(_1550_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_1612_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5470_ (.I(_1613_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5471_ (.I(_1614_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5472_ (.I(_1615_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5473_ (.A1(_1454_),
    .A2(_1605_),
    .B(_1610_),
    .C(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5474_ (.I(_1504_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5475_ (.I0(_1260_),
    .I1(_1153_),
    .S(_1618_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5476_ (.I(_1350_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5477_ (.A1(_1618_),
    .A2(_1282_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5478_ (.A1(_1620_),
    .A2(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5479_ (.A1(_1576_),
    .A2(_1619_),
    .B(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5480_ (.I(_1289_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5481_ (.A1(_1563_),
    .A2(_1623_),
    .B(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5482_ (.I(_0824_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5483_ (.A1(net19),
    .A2(_1538_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5484_ (.I(_0644_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5485_ (.I(_0565_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5486_ (.I0(\reg_file.reg_storage[4][6] ),
    .I1(\reg_file.reg_storage[5][6] ),
    .I2(\reg_file.reg_storage[6][6] ),
    .I3(\reg_file.reg_storage[7][6] ),
    .S0(_1628_),
    .S1(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5487_ (.I0(\reg_file.reg_storage[2][6] ),
    .I1(\reg_file.reg_storage[3][6] ),
    .S(_1081_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5488_ (.I0(\reg_file.reg_storage[1][6] ),
    .I1(_1631_),
    .S(_1629_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5489_ (.I(_0905_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5490_ (.I0(\reg_file.reg_storage[12][6] ),
    .I1(\reg_file.reg_storage[13][6] ),
    .I2(\reg_file.reg_storage[14][6] ),
    .I3(\reg_file.reg_storage[15][6] ),
    .S0(_1633_),
    .S1(_0640_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5491_ (.I0(\reg_file.reg_storage[8][6] ),
    .I1(\reg_file.reg_storage[9][6] ),
    .I2(\reg_file.reg_storage[10][6] ),
    .I3(\reg_file.reg_storage[11][6] ),
    .S0(_1633_),
    .S1(_1629_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5492_ (.I0(_1630_),
    .I1(_1632_),
    .I2(_1634_),
    .I3(_1635_),
    .S0(_0904_),
    .S1(_1086_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5493_ (.I(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5494_ (.A1(_0697_),
    .A2(_1627_),
    .B1(_1637_),
    .B2(_1550_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5495_ (.I(_1638_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5496_ (.I(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5497_ (.A1(_1613_),
    .A2(_1552_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5498_ (.A1(_1477_),
    .A2(_1641_),
    .B(_0656_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5499_ (.A1(_1640_),
    .A2(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5500_ (.A1(_1626_),
    .A2(_1643_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5501_ (.I(_1557_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5502_ (.A1(_0857_),
    .A2(_1556_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5503_ (.A1(_0877_),
    .A2(_1479_),
    .B1(_1556_),
    .B2(_0856_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5504_ (.A1(_1646_),
    .A2(_1647_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5505_ (.A1(_1482_),
    .A2(_1645_),
    .B(_1648_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5506_ (.A1(_1644_),
    .A2(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5507_ (.I(_0539_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5508_ (.A1(_1644_),
    .A2(_1649_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5509_ (.A1(_1651_),
    .A2(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5510_ (.A1(_1092_),
    .A2(_1305_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5511_ (.A1(_1407_),
    .A2(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(_0858_),
    .A2(_0826_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5513_ (.I0(_1524_),
    .I1(_1656_),
    .S(_1353_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5514_ (.A1(_1430_),
    .A2(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5515_ (.A1(_1618_),
    .A2(_1315_),
    .B(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5516_ (.A1(_0824_),
    .A2(_1639_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5517_ (.I(_0523_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5518_ (.A1(_1298_),
    .A2(_1287_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5519_ (.A1(_1661_),
    .A2(_0537_),
    .A3(_1662_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5520_ (.I(_1663_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5521_ (.A1(_0825_),
    .A2(_1640_),
    .B(_1292_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5522_ (.A1(_1626_),
    .A2(_1639_),
    .B(_1665_),
    .C(_1300_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5523_ (.A1(_1655_),
    .A2(_1659_),
    .B1(_1660_),
    .B2(_1664_),
    .C(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5524_ (.A1(_1650_),
    .A2(_1653_),
    .B(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5525_ (.A1(_1617_),
    .A2(_1625_),
    .B(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5526_ (.I(_1669_),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5527_ (.I(_1554_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5528_ (.A1(net20),
    .A2(_1537_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5529_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(\reg_file.reg_storage[5][7] ),
    .I2(\reg_file.reg_storage[6][7] ),
    .I3(\reg_file.reg_storage[7][7] ),
    .S0(_0906_),
    .S1(_1079_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5530_ (.I0(\reg_file.reg_storage[2][7] ),
    .I1(\reg_file.reg_storage[3][7] ),
    .S(_1081_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5531_ (.I0(\reg_file.reg_storage[1][7] ),
    .I1(_1673_),
    .S(_0907_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5532_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(\reg_file.reg_storage[13][7] ),
    .I2(\reg_file.reg_storage[14][7] ),
    .I3(\reg_file.reg_storage[15][7] ),
    .S0(_0924_),
    .S1(_0699_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5533_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(\reg_file.reg_storage[9][7] ),
    .I2(\reg_file.reg_storage[10][7] ),
    .I3(\reg_file.reg_storage[11][7] ),
    .S0(_0924_),
    .S1(_0907_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5534_ (.I0(_1672_),
    .I1(_1674_),
    .I2(_1675_),
    .I3(_1676_),
    .S0(_0707_),
    .S1(_1086_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5535_ (.I(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5536_ (.A1(_0697_),
    .A2(_1671_),
    .B1(_1678_),
    .B2(_1550_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5537_ (.I(_1679_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5538_ (.A1(_1612_),
    .A2(_1551_),
    .A3(_1638_),
    .A4(_1679_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5539_ (.A1(net100),
    .A2(_1681_),
    .B(_1554_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5540_ (.A1(_1477_),
    .A2(_1639_),
    .A3(_1641_),
    .B(_1679_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5541_ (.A1(_1670_),
    .A2(_1680_),
    .B1(_1682_),
    .B2(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5542_ (.A1(_0808_),
    .A2(_1684_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5543_ (.A1(_0825_),
    .A2(_1643_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5544_ (.A1(_1686_),
    .A2(_1652_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5545_ (.A1(_1685_),
    .A2(_1687_),
    .B(_1651_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5546_ (.A1(_1685_),
    .A2(_1687_),
    .B(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5547_ (.I(_1205_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5548_ (.I0(_1396_),
    .I1(_1369_),
    .S(_1690_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5549_ (.A1(_1398_),
    .A2(_1340_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5550_ (.A1(_1350_),
    .A2(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5551_ (.A1(_1486_),
    .A2(_1691_),
    .B(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5552_ (.I(_1407_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5553_ (.I(_1695_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5554_ (.I0(_1427_),
    .I1(_1382_),
    .S(_1461_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5555_ (.A1(_1500_),
    .A2(_1420_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5556_ (.A1(_1583_),
    .A2(_1437_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5557_ (.A1(_1409_),
    .A2(_1698_),
    .A3(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5558_ (.A1(_1696_),
    .A2(_1697_),
    .B(_1700_),
    .C(_1510_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5559_ (.A1(_1485_),
    .A2(_1694_),
    .B(_1701_),
    .C(_1512_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5560_ (.I(_0808_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5561_ (.I(_1680_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5562_ (.I(_1291_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5563_ (.I(_1705_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5564_ (.A1(_0809_),
    .A2(_1704_),
    .B(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5565_ (.A1(_1703_),
    .A2(_1680_),
    .B(_1707_),
    .C(_1516_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5566_ (.A1(_1444_),
    .A2(_1434_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5567_ (.I0(_1590_),
    .I1(_1709_),
    .S(_1467_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5568_ (.I0(_1468_),
    .I1(_1710_),
    .S(_1690_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5569_ (.I(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5570_ (.A1(_0808_),
    .A2(_1704_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5571_ (.A1(_1460_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1532_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5572_ (.A1(_1689_),
    .A2(_1702_),
    .A3(_1708_),
    .A4(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5573_ (.I(_1715_),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5574_ (.A1(_1644_),
    .A2(_1685_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5575_ (.A1(_1475_),
    .A2(_1480_),
    .A3(_1645_),
    .A4(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5576_ (.A1(_1703_),
    .A2(_1684_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5577_ (.A1(_1703_),
    .A2(_1684_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5578_ (.A1(_1686_),
    .A2(_1718_),
    .B1(_1716_),
    .B2(_1648_),
    .C(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5579_ (.A1(_1717_),
    .A2(_1720_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5580_ (.A1(net21),
    .A2(_1538_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5581_ (.I(_1543_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5582_ (.I(_0703_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5583_ (.I(_1724_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5584_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(\reg_file.reg_storage[5][8] ),
    .I2(\reg_file.reg_storage[6][8] ),
    .I3(\reg_file.reg_storage[7][8] ),
    .S0(_1723_),
    .S1(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5585_ (.I0(\reg_file.reg_storage[2][8] ),
    .I1(\reg_file.reg_storage[3][8] ),
    .S(_0906_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5586_ (.I(_0559_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5587_ (.I0(\reg_file.reg_storage[1][8] ),
    .I1(_1727_),
    .S(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5588_ (.I(_1543_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5589_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(\reg_file.reg_storage[13][8] ),
    .I2(\reg_file.reg_storage[14][8] ),
    .I3(\reg_file.reg_storage[15][8] ),
    .S0(_1730_),
    .S1(_1728_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5590_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(\reg_file.reg_storage[9][8] ),
    .I2(\reg_file.reg_storage[10][8] ),
    .I3(\reg_file.reg_storage[11][8] ),
    .S0(_1730_),
    .S1(_1728_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5591_ (.I0(_1726_),
    .I1(_1729_),
    .I2(_1731_),
    .I3(_1732_),
    .S0(_0920_),
    .S1(_0928_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5592_ (.I(_1733_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5593_ (.I(_0903_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5594_ (.A1(_1536_),
    .A2(_1722_),
    .B1(_1734_),
    .B2(_1735_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5595_ (.I(_1736_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5596_ (.A1(_1682_),
    .A2(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5597_ (.A1(_0782_),
    .A2(_1738_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5598_ (.A1(_1721_),
    .A2(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5599_ (.A1(_1721_),
    .A2(_1739_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5600_ (.A1(_1325_),
    .A2(_1740_),
    .A3(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5601_ (.I(_1614_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5602_ (.A1(_1695_),
    .A2(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5603_ (.I(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5604_ (.I0(_1488_),
    .I1(_1491_),
    .S(_0720_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5605_ (.I0(_1501_),
    .I1(_1497_),
    .S(_0721_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5606_ (.I0(_1496_),
    .I1(_1487_),
    .S(_0720_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5607_ (.I0(_1747_),
    .I1(_1748_),
    .S(_1575_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5608_ (.I(_1615_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5609_ (.A1(_1745_),
    .A2(_1746_),
    .B1(_1749_),
    .B2(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5610_ (.A1(_0784_),
    .A2(_0810_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5611_ (.I0(_1656_),
    .I1(_1752_),
    .S(_1564_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5612_ (.I0(_1526_),
    .I1(_1753_),
    .S(_1504_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5613_ (.A1(_0937_),
    .A2(_1527_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5614_ (.I0(_1754_),
    .I1(_1755_),
    .S(_1575_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5615_ (.I(_1737_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5616_ (.A1(_0783_),
    .A2(_1757_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5617_ (.I(_0783_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5618_ (.A1(_1759_),
    .A2(_1757_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5619_ (.A1(_1457_),
    .A2(_1760_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5620_ (.I(_1514_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5621_ (.A1(_1759_),
    .A2(_1757_),
    .B(_1761_),
    .C(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5622_ (.A1(_1306_),
    .A2(_1756_),
    .B1(_1758_),
    .B2(_1664_),
    .C(_1763_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5623_ (.A1(_1624_),
    .A2(_1751_),
    .B(_1764_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5624_ (.A1(_1742_),
    .A2(_1765_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5625_ (.I(_1654_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5626_ (.A1(_1431_),
    .A2(_1435_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5627_ (.I(_1208_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5628_ (.I0(_1709_),
    .I1(_1767_),
    .S(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5629_ (.I0(_1591_),
    .I1(_1769_),
    .S(_1504_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5630_ (.I(_1207_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5631_ (.I(_1771_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5632_ (.I(_0838_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5633_ (.A1(_1773_),
    .A2(_1522_),
    .A3(_1464_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5634_ (.A1(_1772_),
    .A2(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5635_ (.A1(_1454_),
    .A2(_1770_),
    .B(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5636_ (.I(_0746_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5637_ (.I(_0637_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5638_ (.A1(net22),
    .A2(_1538_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5639_ (.I(_1724_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5640_ (.I0(\reg_file.reg_storage[4][9] ),
    .I1(\reg_file.reg_storage[5][9] ),
    .I2(\reg_file.reg_storage[6][9] ),
    .I3(\reg_file.reg_storage[7][9] ),
    .S0(_1723_),
    .S1(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5641_ (.I0(\reg_file.reg_storage[2][9] ),
    .I1(\reg_file.reg_storage[3][9] ),
    .S(_0921_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5642_ (.I0(\reg_file.reg_storage[1][9] ),
    .I1(_1782_),
    .S(_1725_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5643_ (.I0(\reg_file.reg_storage[12][9] ),
    .I1(\reg_file.reg_storage[13][9] ),
    .I2(\reg_file.reg_storage[14][9] ),
    .I3(\reg_file.reg_storage[15][9] ),
    .S0(_1723_),
    .S1(_1725_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5644_ (.I0(\reg_file.reg_storage[8][9] ),
    .I1(\reg_file.reg_storage[9][9] ),
    .I2(\reg_file.reg_storage[10][9] ),
    .I3(\reg_file.reg_storage[11][9] ),
    .S0(_1723_),
    .S1(_1725_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5645_ (.I0(_1781_),
    .I1(_1783_),
    .I2(_1784_),
    .I3(_1785_),
    .S0(_0920_),
    .S1(_0918_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5646_ (.I(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5647_ (.A1(_1778_),
    .A2(_1779_),
    .B1(_1787_),
    .B2(_1735_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5648_ (.I(_1788_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5649_ (.I(_1789_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5650_ (.I(_1661_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5651_ (.A1(_1777_),
    .A2(_1790_),
    .B(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5652_ (.A1(_1777_),
    .A2(_1790_),
    .B(_1515_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5653_ (.A1(_0744_),
    .A2(_1789_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5654_ (.A1(_1792_),
    .A2(_1793_),
    .B1(_1794_),
    .B2(_1664_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5655_ (.I(_0661_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5656_ (.A1(_1682_),
    .A2(_1737_),
    .B(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5657_ (.A1(_0745_),
    .A2(_1789_),
    .A3(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5658_ (.A1(_1759_),
    .A2(_1738_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5659_ (.A1(_1799_),
    .A2(_1740_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5660_ (.A1(_1798_),
    .A2(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5661_ (.A1(_0936_),
    .A2(_1304_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5662_ (.I(_1503_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5663_ (.I0(_1565_),
    .I1(_1568_),
    .S(_1803_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5664_ (.I(_1303_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5665_ (.I0(_1581_),
    .I1(_1569_),
    .S(_1461_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5666_ (.A1(_1805_),
    .A2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5667_ (.I(_1408_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5668_ (.I0(_1579_),
    .I1(_1584_),
    .S(_1397_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5669_ (.A1(_1808_),
    .A2(_1809_),
    .B(_1743_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5670_ (.A1(_1802_),
    .A2(_1804_),
    .B1(_1807_),
    .B2(_1810_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5671_ (.I(_0538_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5672_ (.A1(_1481_),
    .A2(_1801_),
    .B1(_1811_),
    .B2(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5673_ (.A1(_1766_),
    .A2(_1776_),
    .B(_1795_),
    .C(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5674_ (.I(_1814_),
    .ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5675_ (.A1(_1739_),
    .A2(_1798_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5676_ (.A1(_1790_),
    .A2(_1797_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5677_ (.A1(_0746_),
    .A2(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5678_ (.A1(_0745_),
    .A2(_1816_),
    .B(_1799_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5679_ (.A1(_1817_),
    .A2(_1818_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5680_ (.A1(_1721_),
    .A2(_1815_),
    .B(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5681_ (.I(_1537_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5682_ (.A1(net24),
    .A2(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5683_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(\reg_file.reg_storage[5][10] ),
    .I2(\reg_file.reg_storage[6][10] ),
    .I3(\reg_file.reg_storage[7][10] ),
    .S0(_1730_),
    .S1(_1728_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5684_ (.I0(\reg_file.reg_storage[2][10] ),
    .I1(\reg_file.reg_storage[3][10] ),
    .S(_0924_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5685_ (.I(_0703_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5686_ (.I0(\reg_file.reg_storage[1][10] ),
    .I1(_1824_),
    .S(_1825_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5687_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(\reg_file.reg_storage[13][10] ),
    .I2(\reg_file.reg_storage[14][10] ),
    .I3(\reg_file.reg_storage[15][10] ),
    .S0(_0910_),
    .S1(_1825_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5688_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(\reg_file.reg_storage[9][10] ),
    .I2(\reg_file.reg_storage[10][10] ),
    .I3(\reg_file.reg_storage[11][10] ),
    .S0(_1730_),
    .S1(_1825_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5689_ (.I0(_1823_),
    .I1(_1826_),
    .I2(_1827_),
    .I3(_1828_),
    .S0(_0920_),
    .S1(_0928_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5690_ (.I(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5691_ (.A1(_1536_),
    .A2(_1822_),
    .B1(_1830_),
    .B2(_1735_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5692_ (.I(_1831_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5693_ (.I(_1832_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _5694_ (.A1(_1613_),
    .A2(_1552_),
    .A3(_1638_),
    .A4(_1679_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5695_ (.A1(_1737_),
    .A2(_1789_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5696_ (.I(_0661_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5697_ (.A1(_1476_),
    .A2(_1834_),
    .A3(_1835_),
    .B(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5698_ (.A1(_1833_),
    .A2(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5699_ (.A1(_1013_),
    .A2(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5700_ (.A1(_1820_),
    .A2(_1839_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5701_ (.I(_1324_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5702_ (.A1(_1820_),
    .A2(_1839_),
    .B(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5703_ (.A1(_1840_),
    .A2(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5704_ (.I(_1695_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5705_ (.A1(_1015_),
    .A2(_0747_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5706_ (.A1(_1387_),
    .A2(_1752_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5707_ (.A1(_1438_),
    .A2(_1845_),
    .B(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5708_ (.I(_1503_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5709_ (.I0(_1657_),
    .I1(_1847_),
    .S(_1848_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5710_ (.A1(_1808_),
    .A2(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5711_ (.A1(_1844_),
    .A2(_1316_),
    .B(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5712_ (.I(_1802_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5713_ (.I(_1303_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5714_ (.A1(_1019_),
    .A2(_1074_),
    .B(_1608_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5715_ (.A1(_1853_),
    .A2(_1206_),
    .B(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5716_ (.I(_1093_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5717_ (.A1(_1284_),
    .A2(_1852_),
    .B1(_1855_),
    .B2(_1856_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5718_ (.I(_1812_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5719_ (.I(_1014_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5720_ (.A1(_1859_),
    .A2(_1831_),
    .B(_1661_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5721_ (.A1(_1014_),
    .A2(_1833_),
    .B(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5722_ (.A1(_1012_),
    .A2(_1833_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5723_ (.A1(_1515_),
    .A2(_1861_),
    .B1(_1862_),
    .B2(_1471_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5724_ (.A1(_1306_),
    .A2(_1851_),
    .B1(_1857_),
    .B2(_1858_),
    .C(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5725_ (.A1(_1843_),
    .A2(_1864_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_1865_),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5727_ (.I(_1651_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5728_ (.I(_0988_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5729_ (.I(_0553_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5730_ (.I(_1081_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5731_ (.I(_1869_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5732_ (.I(_1870_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5733_ (.I(_0552_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5734_ (.A1(_0693_),
    .A2(_1872_),
    .A3(_1868_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5735_ (.I(net25),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _5736_ (.A1(net30),
    .A2(_0693_),
    .B1(_1868_),
    .B2(_1871_),
    .C1(_1873_),
    .C2(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5737_ (.I(_1543_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5738_ (.I(_0570_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5739_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(\reg_file.reg_storage[5][11] ),
    .I2(\reg_file.reg_storage[6][11] ),
    .I3(\reg_file.reg_storage[7][11] ),
    .S0(_1876_),
    .S1(_1877_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5740_ (.I0(\reg_file.reg_storage[2][11] ),
    .I1(\reg_file.reg_storage[3][11] ),
    .S(_1633_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5741_ (.I0(\reg_file.reg_storage[1][11] ),
    .I1(_1879_),
    .S(_1780_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5742_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(\reg_file.reg_storage[13][11] ),
    .I2(\reg_file.reg_storage[14][11] ),
    .I3(\reg_file.reg_storage[15][11] ),
    .S0(_1876_),
    .S1(_1780_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5743_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(\reg_file.reg_storage[9][11] ),
    .I2(\reg_file.reg_storage[10][11] ),
    .I3(\reg_file.reg_storage[11][11] ),
    .S0(_1876_),
    .S1(_1780_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5744_ (.I0(_1878_),
    .I1(_1880_),
    .I2(_1881_),
    .I3(_1882_),
    .S0(_0692_),
    .S1(_0918_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5745_ (.I(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5746_ (.A1(_1778_),
    .A2(_1875_),
    .B1(_1884_),
    .B2(_1735_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5747_ (.I(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5748_ (.I(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5749_ (.A1(_1477_),
    .A2(_1834_),
    .A3(_1831_),
    .A4(_1835_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5750_ (.A1(_1670_),
    .A2(_1888_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5751_ (.A1(_1867_),
    .A2(_1887_),
    .A3(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5752_ (.A1(_1013_),
    .A2(_1838_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5753_ (.A1(_1891_),
    .A2(_1840_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5754_ (.A1(_1890_),
    .A2(_1892_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5755_ (.A1(_1432_),
    .A2(_1412_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5756_ (.I0(_1767_),
    .I1(_1894_),
    .S(_0833_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5757_ (.I0(_1710_),
    .I1(_1895_),
    .S(_1848_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5758_ (.A1(_1608_),
    .A2(_1469_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5759_ (.A1(_1384_),
    .A2(_1896_),
    .B(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5760_ (.A1(_0989_),
    .A2(_1887_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5761_ (.I(_1319_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5762_ (.I(_1900_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5763_ (.I(_1292_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5764_ (.I(_1867_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5765_ (.A1(_1903_),
    .A2(_1886_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5766_ (.I(_1299_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5767_ (.A1(_1903_),
    .A2(_1886_),
    .B(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5768_ (.A1(_1902_),
    .A2(_1904_),
    .B(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5769_ (.A1(_1766_),
    .A2(_1898_),
    .B1(_1899_),
    .B2(_1901_),
    .C(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5770_ (.I0(_1428_),
    .I1(_1383_),
    .S(_1575_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5771_ (.A1(_1403_),
    .A2(_1852_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5772_ (.A1(_1616_),
    .A2(_1909_),
    .B(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5773_ (.A1(_1624_),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5774_ (.A1(_1866_),
    .A2(_1893_),
    .B(_1908_),
    .C(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5775_ (.I(_1913_),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5776_ (.I(_1802_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5777_ (.A1(_1495_),
    .A2(_1499_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5778_ (.A1(_1454_),
    .A2(_1489_),
    .B(_1750_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5779_ (.A1(_1492_),
    .A2(_1914_),
    .B1(_1915_),
    .B2(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5780_ (.A1(_0976_),
    .A2(_0990_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5781_ (.A1(_1467_),
    .A2(_1845_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5782_ (.A1(_1438_),
    .A2(_1918_),
    .B(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5783_ (.I0(_1753_),
    .I1(_1920_),
    .S(_1803_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5784_ (.A1(_1351_),
    .A2(_1529_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5785_ (.A1(_1609_),
    .A2(_1921_),
    .B(_1922_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5786_ (.I(_0975_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5787_ (.A1(_1872_),
    .A2(_1868_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5788_ (.A1(_0551_),
    .A2(_0553_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5789_ (.A1(net25),
    .A2(_1926_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5790_ (.A1(net4),
    .A2(_1925_),
    .B(_1927_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5791_ (.I(_1076_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5792_ (.I(_1628_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5793_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(\reg_file.reg_storage[5][12] ),
    .I2(\reg_file.reg_storage[6][12] ),
    .I3(\reg_file.reg_storage[7][12] ),
    .S0(_1930_),
    .S1(_0915_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5794_ (.I(_0913_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5795_ (.I(_1876_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5796_ (.A1(_1933_),
    .A2(\reg_file.reg_storage[3][12] ),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5797_ (.I(_0547_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5798_ (.I(_0912_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5799_ (.A1(_1935_),
    .A2(\reg_file.reg_storage[2][12] ),
    .B(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5800_ (.A1(_1932_),
    .A2(_0965_),
    .B1(_1934_),
    .B2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5801_ (.I(_1633_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5802_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(\reg_file.reg_storage[13][12] ),
    .I2(\reg_file.reg_storage[14][12] ),
    .I3(\reg_file.reg_storage[15][12] ),
    .S0(_1939_),
    .S1(_1877_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5803_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(\reg_file.reg_storage[9][12] ),
    .I2(\reg_file.reg_storage[10][12] ),
    .I3(\reg_file.reg_storage[11][12] ),
    .S0(_1939_),
    .S1(_0915_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5804_ (.I(_0707_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5805_ (.I(_0708_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5806_ (.I0(_1931_),
    .I1(_1938_),
    .I2(_1940_),
    .I3(_1941_),
    .S0(_1942_),
    .S1(_1943_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(_1929_),
    .A2(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5808_ (.A1(_1778_),
    .A2(_1928_),
    .B(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5809_ (.I(_1946_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5810_ (.I(_1947_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5811_ (.A1(_1924_),
    .A2(_1948_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5812_ (.I(_1924_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5813_ (.A1(_1950_),
    .A2(_1948_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5814_ (.A1(_1950_),
    .A2(_1948_),
    .B(_1905_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5815_ (.A1(_1902_),
    .A2(_1951_),
    .B(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5816_ (.A1(_1654_),
    .A2(_1923_),
    .B1(_1949_),
    .B2(_1471_),
    .C(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5817_ (.A1(_1736_),
    .A2(_1788_),
    .A3(_1885_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5818_ (.A1(net100),
    .A2(_1681_),
    .A3(_1832_),
    .A4(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5819_ (.I(_1956_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5820_ (.A1(_0662_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5821_ (.A1(_1947_),
    .A2(_1958_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5822_ (.A1(_1950_),
    .A2(_1959_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5823_ (.A1(_1839_),
    .A2(_1890_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5824_ (.A1(_1815_),
    .A2(_1961_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5825_ (.A1(_1817_),
    .A2(_1818_),
    .A3(_1839_),
    .A4(_1890_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5826_ (.A1(_1887_),
    .A2(_1889_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5827_ (.A1(_1903_),
    .A2(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5828_ (.A1(_1903_),
    .A2(_1964_),
    .B(_1891_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5829_ (.A1(_1965_),
    .A2(_1966_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5830_ (.A1(_1721_),
    .A2(_1962_),
    .B(_1963_),
    .C(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5831_ (.A1(_1960_),
    .A2(_1968_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5832_ (.A1(_1651_),
    .A2(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5833_ (.A1(_1960_),
    .A2(_1968_),
    .B(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5834_ (.A1(_1858_),
    .A2(_1917_),
    .B(_1954_),
    .C(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5835_ (.I(_1972_),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5836_ (.A1(net5),
    .A2(_1925_),
    .B(_1927_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _5837_ (.I(_1540_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5838_ (.I(_1724_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5839_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(\reg_file.reg_storage[5][13] ),
    .I2(\reg_file.reg_storage[6][13] ),
    .I3(\reg_file.reg_storage[7][13] ),
    .S0(_1974_),
    .S1(_1975_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5840_ (.I(_1869_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5841_ (.A1(_1977_),
    .A2(\reg_file.reg_storage[3][13] ),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5842_ (.A1(_1935_),
    .A2(\reg_file.reg_storage[2][13] ),
    .B(_1936_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5843_ (.A1(_1932_),
    .A2(_0946_),
    .B1(_1978_),
    .B2(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5844_ (.I(_1724_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5845_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(\reg_file.reg_storage[13][13] ),
    .I2(\reg_file.reg_storage[14][13] ),
    .I3(\reg_file.reg_storage[15][13] ),
    .S0(_1930_),
    .S1(_1981_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5846_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(\reg_file.reg_storage[9][13] ),
    .I2(\reg_file.reg_storage[10][13] ),
    .I3(\reg_file.reg_storage[11][13] ),
    .S0(_1930_),
    .S1(_1981_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5847_ (.I0(_1976_),
    .I1(_1980_),
    .I2(_1982_),
    .I3(_1983_),
    .S0(_1942_),
    .S1(_1943_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5848_ (.A1(_1929_),
    .A2(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5849_ (.A1(_1778_),
    .A2(_1973_),
    .B(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5850_ (.I(_1986_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5851_ (.I(_1987_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5852_ (.A1(_1415_),
    .A2(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5853_ (.A1(_1518_),
    .A2(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5854_ (.A1(_1415_),
    .A2(_1988_),
    .B(_1990_),
    .C(_1516_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5855_ (.A1(_1354_),
    .A2(_1415_),
    .B(_1410_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5856_ (.I0(_1894_),
    .I1(_1992_),
    .S(_1768_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5857_ (.I0(_1769_),
    .I1(_1993_),
    .S(_1803_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5858_ (.A1(_1486_),
    .A2(_1594_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5859_ (.A1(_1805_),
    .A2(_1994_),
    .B(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5860_ (.A1(_0959_),
    .A2(_1988_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5861_ (.I(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5862_ (.A1(_1766_),
    .A2(_1996_),
    .B1(_1998_),
    .B2(_1532_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5863_ (.A1(_1950_),
    .A2(_1959_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5864_ (.A1(_1947_),
    .A2(net110),
    .B(_1836_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5865_ (.A1(_1987_),
    .A2(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5866_ (.A1(_0959_),
    .A2(_2002_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5867_ (.A1(_2000_),
    .A2(_1969_),
    .B(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5868_ (.A1(_2000_),
    .A2(_1969_),
    .A3(_2003_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5869_ (.A1(_1481_),
    .A2(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5870_ (.I(_1743_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5871_ (.A1(_1582_),
    .A2(_1585_),
    .B(_1351_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5872_ (.I(_1303_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5873_ (.A1(_2009_),
    .A2(_1571_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5874_ (.A1(_2007_),
    .A2(_2008_),
    .A3(_2010_),
    .B1(_1566_),
    .B2(_1745_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5875_ (.A1(_2004_),
    .A2(_2006_),
    .B1(_2011_),
    .B2(_1624_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5876_ (.A1(_1991_),
    .A2(_1999_),
    .A3(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5877_ (.I(_2013_),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5878_ (.A1(_1696_),
    .A2(_1605_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5879_ (.A1(_1495_),
    .A2(_1619_),
    .B(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5880_ (.A1(_1621_),
    .A2(_1914_),
    .B1(_2015_),
    .B2(_1485_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5881_ (.I(_0901_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5882_ (.I(_1381_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5883_ (.A1(_1365_),
    .A2(_1058_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5884_ (.A1(_1414_),
    .A2(_0960_),
    .B(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5885_ (.A1(_1401_),
    .A2(_2020_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5886_ (.A1(_2018_),
    .A2(_1918_),
    .B(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5887_ (.A1(_2017_),
    .A2(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5888_ (.A1(_1430_),
    .A2(_1847_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5889_ (.A1(_2023_),
    .A2(_2024_),
    .B(_1429_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5890_ (.A1(_1844_),
    .A2(_1659_),
    .B(_2025_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5891_ (.A1(_0482_),
    .A2(_1925_),
    .B(_1927_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5892_ (.I0(\reg_file.reg_storage[4][14] ),
    .I1(\reg_file.reg_storage[5][14] ),
    .I2(\reg_file.reg_storage[6][14] ),
    .I3(\reg_file.reg_storage[7][14] ),
    .S0(_1974_),
    .S1(_1975_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(_1977_),
    .A2(\reg_file.reg_storage[3][14] ),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5894_ (.A1(_1935_),
    .A2(\reg_file.reg_storage[2][14] ),
    .B(_1936_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5895_ (.A1(_1932_),
    .A2(_1049_),
    .B1(_2029_),
    .B2(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5896_ (.I0(\reg_file.reg_storage[12][14] ),
    .I1(\reg_file.reg_storage[13][14] ),
    .I2(\reg_file.reg_storage[14][14] ),
    .I3(\reg_file.reg_storage[15][14] ),
    .S0(_1930_),
    .S1(_1981_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5897_ (.I0(\reg_file.reg_storage[8][14] ),
    .I1(\reg_file.reg_storage[9][14] ),
    .I2(\reg_file.reg_storage[10][14] ),
    .I3(\reg_file.reg_storage[11][14] ),
    .S0(_1974_),
    .S1(_1981_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5898_ (.I0(_2028_),
    .I1(_2031_),
    .I2(_2032_),
    .I3(_2033_),
    .S0(_1942_),
    .S1(_1943_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5899_ (.A1(_1929_),
    .A2(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5900_ (.A1(_0698_),
    .A2(_2027_),
    .B(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5901_ (.I(_2036_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5902_ (.I(_2037_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5903_ (.A1(_1057_),
    .A2(_2038_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5904_ (.A1(_1058_),
    .A2(_2038_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5905_ (.A1(_1058_),
    .A2(_2038_),
    .B(_1905_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5906_ (.A1(_1902_),
    .A2(_2040_),
    .B(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5907_ (.A1(_1766_),
    .A2(_2026_),
    .B1(_2039_),
    .B2(_1901_),
    .C(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5908_ (.I(_1324_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5909_ (.A1(_0960_),
    .A2(_2002_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5910_ (.A1(_0960_),
    .A2(_2002_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5911_ (.A1(_2000_),
    .A2(_2045_),
    .B(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5912_ (.A1(_1960_),
    .A2(_1968_),
    .A3(_2003_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5913_ (.A1(_2047_),
    .A2(_2048_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5914_ (.A1(_1946_),
    .A2(_1987_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5915_ (.A1(_1957_),
    .A2(_2050_),
    .B(_1836_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5916_ (.A1(_2037_),
    .A2(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5917_ (.A1(_1417_),
    .A2(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5918_ (.A1(_1417_),
    .A2(_2052_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5919_ (.A1(_2053_),
    .A2(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5920_ (.A1(_2049_),
    .A2(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5921_ (.A1(_2049_),
    .A2(_2055_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5922_ (.A1(_2044_),
    .A2(_2056_),
    .A3(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5923_ (.A1(_1858_),
    .A2(_2016_),
    .B(_2043_),
    .C(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5924_ (.I(_2059_),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5925_ (.A1(_1418_),
    .A2(_1425_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5926_ (.I0(_1992_),
    .I1(_2060_),
    .S(_0832_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5927_ (.I0(_1895_),
    .I1(_2061_),
    .S(_1447_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5928_ (.A1(_1429_),
    .A2(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5929_ (.A1(_1808_),
    .A2(_1712_),
    .B(_2063_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5930_ (.I(_1069_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5931_ (.I(_1926_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5932_ (.A1(net25),
    .A2(_0552_),
    .A3(_1868_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5933_ (.I(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5934_ (.A1(_0735_),
    .A2(_2066_),
    .B(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5935_ (.A1(_0690_),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5936_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(\reg_file.reg_storage[5][15] ),
    .I2(\reg_file.reg_storage[6][15] ),
    .I3(\reg_file.reg_storage[7][15] ),
    .S0(_1939_),
    .S1(_0915_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5937_ (.I(_0913_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5938_ (.A1(_1933_),
    .A2(\reg_file.reg_storage[3][15] ),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5939_ (.A1(_1935_),
    .A2(\reg_file.reg_storage[2][15] ),
    .B(_1936_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5940_ (.A1(_2072_),
    .A2(_1061_),
    .B1(_2073_),
    .B2(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5941_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(\reg_file.reg_storage[13][15] ),
    .I2(\reg_file.reg_storage[14][15] ),
    .I3(\reg_file.reg_storage[15][15] ),
    .S0(_1869_),
    .S1(_1877_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5942_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(\reg_file.reg_storage[9][15] ),
    .I2(\reg_file.reg_storage[10][15] ),
    .I3(\reg_file.reg_storage[11][15] ),
    .S0(_1939_),
    .S1(_1877_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5943_ (.I0(_2071_),
    .I1(_2075_),
    .I2(_2076_),
    .I3(_2077_),
    .S0(_1942_),
    .S1(_0918_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5944_ (.A1(_1076_),
    .A2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5945_ (.A1(_2070_),
    .A2(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5946_ (.I(_2080_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5947_ (.A1(_2065_),
    .A2(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5948_ (.A1(_2065_),
    .A2(_2081_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5949_ (.A1(_1706_),
    .A2(_2082_),
    .B(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5950_ (.A1(_1069_),
    .A2(_2081_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5951_ (.I(_1900_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5952_ (.A1(_1516_),
    .A2(_2084_),
    .B1(_2085_),
    .B2(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5953_ (.A1(_1957_),
    .A2(_2037_),
    .A3(_2050_),
    .B(_1796_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5954_ (.A1(_2080_),
    .A2(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5955_ (.A1(_1069_),
    .A2(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5956_ (.A1(_2053_),
    .A2(_2057_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5957_ (.A1(_2090_),
    .A2(_2091_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5958_ (.I0(_1697_),
    .I1(_1691_),
    .S(_1608_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5959_ (.A1(_1398_),
    .A2(_1340_),
    .A3(_1744_),
    .B1(_2093_),
    .B2(_1750_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5960_ (.A1(_2044_),
    .A2(_2092_),
    .B1(_2094_),
    .B2(_1512_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5961_ (.A1(_1306_),
    .A2(_2064_),
    .B(_2087_),
    .C(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5962_ (.I(_2096_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5963_ (.I(_0690_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5964_ (.A1(_0770_),
    .A2(_2066_),
    .B(_2068_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5965_ (.A1(_2097_),
    .A2(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5966_ (.I(_1076_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5967_ (.I(_0910_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5968_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(\reg_file.reg_storage[5][16] ),
    .I2(\reg_file.reg_storage[6][16] ),
    .I3(\reg_file.reg_storage[7][16] ),
    .S0(_2101_),
    .S1(_0641_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5969_ (.I(_0913_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5970_ (.A1(_1870_),
    .A2(\reg_file.reg_storage[3][16] ),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5971_ (.I(_0548_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5972_ (.I(_0912_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5973_ (.A1(_2105_),
    .A2(\reg_file.reg_storage[2][16] ),
    .B(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5974_ (.A1(_2103_),
    .A2(_1036_),
    .B1(_2104_),
    .B2(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5975_ (.I(_0910_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5976_ (.I(_0640_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5977_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(\reg_file.reg_storage[13][16] ),
    .I2(\reg_file.reg_storage[14][16] ),
    .I3(\reg_file.reg_storage[15][16] ),
    .S0(_2109_),
    .S1(_2110_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5978_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(\reg_file.reg_storage[9][16] ),
    .I2(\reg_file.reg_storage[10][16] ),
    .I3(\reg_file.reg_storage[11][16] ),
    .S0(_2101_),
    .S1(_2110_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5979_ (.I(_0904_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5980_ (.I(_0708_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5981_ (.I0(_2102_),
    .I1(_2108_),
    .I2(_2111_),
    .I3(_2112_),
    .S0(_2113_),
    .S1(_2114_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5982_ (.A1(_2100_),
    .A2(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5983_ (.A1(_2099_),
    .A2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5984_ (.I(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5985_ (.A1(net101),
    .A2(_1681_),
    .A3(_1833_),
    .A4(_1955_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5986_ (.A1(_1947_),
    .A2(_1987_),
    .A3(_2037_),
    .A4(_2080_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5987_ (.A1(_2119_),
    .A2(_2120_),
    .B(_1670_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5988_ (.A1(_2118_),
    .A2(_2121_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5989_ (.A1(_1044_),
    .A2(_2122_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5990_ (.I(_2123_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5991_ (.A1(_1056_),
    .A2(_2052_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5992_ (.A1(_1960_),
    .A2(_2003_),
    .A3(_2125_),
    .A4(_2090_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5993_ (.A1(_1963_),
    .A2(_1967_),
    .B(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5994_ (.A1(_1717_),
    .A2(_1720_),
    .B(_1962_),
    .C(_2126_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5995_ (.A1(_1070_),
    .A2(_2089_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5996_ (.A1(_2065_),
    .A2(_2089_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5997_ (.A1(_2053_),
    .A2(_2130_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5998_ (.A1(_2065_),
    .A2(_2089_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5999_ (.A1(_2047_),
    .A2(_2055_),
    .A3(_2129_),
    .B1(_2131_),
    .B2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _6000_ (.A1(_2127_),
    .A2(_2128_),
    .A3(_2133_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6001_ (.A1(_2124_),
    .A2(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6002_ (.A1(_2124_),
    .A2(_2134_),
    .B(_2044_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6003_ (.I(_1305_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6004_ (.I(_2137_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6005_ (.I(_2138_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6006_ (.A1(_1045_),
    .A2(_1071_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6007_ (.A1(_1381_),
    .A2(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6008_ (.A1(_1309_),
    .A2(_2020_),
    .B(_2141_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6009_ (.I0(_1920_),
    .I1(_2142_),
    .S(_1848_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6010_ (.I0(_1754_),
    .I1(_2143_),
    .S(_1572_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6011_ (.A1(_1755_),
    .A2(_1745_),
    .B1(_2144_),
    .B2(_1750_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6012_ (.A1(_2139_),
    .A2(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6013_ (.A1(_1812_),
    .A2(_1614_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6014_ (.I(_2147_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6015_ (.I(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6016_ (.I(_1746_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6017_ (.A1(_1406_),
    .A2(_1748_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6018_ (.A1(_1406_),
    .A2(_2150_),
    .B(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6019_ (.I(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6020_ (.I(_1043_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6021_ (.I(_2118_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6022_ (.A1(_2154_),
    .A2(_2155_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6023_ (.I(_1705_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6024_ (.A1(_2154_),
    .A2(_2155_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6025_ (.I(_1514_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6026_ (.A1(_2154_),
    .A2(_2155_),
    .B(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6027_ (.A1(_2157_),
    .A2(_2158_),
    .B(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6028_ (.A1(_2149_),
    .A2(_2153_),
    .B1(_2156_),
    .B2(_2086_),
    .C(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6029_ (.A1(_2135_),
    .A2(_2136_),
    .B(_2146_),
    .C(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6030_ (.I(_2163_),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6031_ (.A1(_1044_),
    .A2(_2122_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6032_ (.A1(_2164_),
    .A2(_2135_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6033_ (.I(_1029_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6034_ (.I(_1926_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6035_ (.I(_2067_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6036_ (.A1(_0603_),
    .A2(_2167_),
    .B(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6037_ (.A1(_2097_),
    .A2(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6038_ (.I0(\reg_file.reg_storage[4][17] ),
    .I1(\reg_file.reg_storage[5][17] ),
    .I2(\reg_file.reg_storage[6][17] ),
    .I3(\reg_file.reg_storage[7][17] ),
    .S0(_2101_),
    .S1(_0641_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6039_ (.A1(_1870_),
    .A2(\reg_file.reg_storage[3][17] ),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6040_ (.A1(_2105_),
    .A2(\reg_file.reg_storage[2][17] ),
    .B(_2072_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6041_ (.A1(_2103_),
    .A2(_1022_),
    .B1(_2172_),
    .B2(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6042_ (.I0(\reg_file.reg_storage[12][17] ),
    .I1(\reg_file.reg_storage[13][17] ),
    .I2(\reg_file.reg_storage[14][17] ),
    .I3(\reg_file.reg_storage[15][17] ),
    .S0(_2109_),
    .S1(_2110_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6043_ (.I0(\reg_file.reg_storage[8][17] ),
    .I1(\reg_file.reg_storage[9][17] ),
    .I2(\reg_file.reg_storage[10][17] ),
    .I3(\reg_file.reg_storage[11][17] ),
    .S0(_2101_),
    .S1(_0641_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6044_ (.I0(_2171_),
    .I1(_2174_),
    .I2(_2175_),
    .I3(_2176_),
    .S0(_2113_),
    .S1(_2114_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6045_ (.A1(_2100_),
    .A2(_2177_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6046_ (.A1(_2170_),
    .A2(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6047_ (.I(_2179_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6048_ (.I(_2180_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6049_ (.I(_0659_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6050_ (.A1(_2155_),
    .A2(_2121_),
    .B(_2182_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6051_ (.A1(_2166_),
    .A2(_2181_),
    .A3(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6052_ (.A1(_2165_),
    .A2(_2184_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(_1914_),
    .A2(_1774_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6054_ (.A1(_1422_),
    .A2(_1424_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6055_ (.I0(_2060_),
    .I1(_2187_),
    .S(_1768_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6056_ (.I0(_1993_),
    .I1(_2188_),
    .S(_1803_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6057_ (.I(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6058_ (.A1(_1853_),
    .A2(_1770_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6059_ (.A1(_1609_),
    .A2(_2190_),
    .B(_2191_),
    .C(_1856_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6060_ (.A1(_2186_),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6061_ (.A1(_2139_),
    .A2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6062_ (.A1(_1805_),
    .A2(_1804_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6063_ (.A1(_1620_),
    .A2(_1806_),
    .B(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6064_ (.A1(_2166_),
    .A2(_2180_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6065_ (.I(_2166_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6066_ (.A1(_2198_),
    .A2(_2181_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6067_ (.A1(_2198_),
    .A2(_2181_),
    .B(_2159_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6068_ (.A1(_2157_),
    .A2(_2199_),
    .B(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6069_ (.A1(_2148_),
    .A2(_2196_),
    .B1(_2197_),
    .B2(_1901_),
    .C(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6070_ (.A1(_1866_),
    .A2(_2185_),
    .B(_2194_),
    .C(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6071_ (.I(_2203_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6072_ (.A1(_2181_),
    .A2(_2183_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6073_ (.A1(_2198_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6074_ (.A1(_2198_),
    .A2(_2204_),
    .B(_2164_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6075_ (.A1(_2205_),
    .A2(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6076_ (.A1(_2124_),
    .A2(_2134_),
    .A3(_2184_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6077_ (.I(_1201_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6078_ (.A1(_0629_),
    .A2(_2066_),
    .B(_2068_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6079_ (.A1(_2097_),
    .A2(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6080_ (.I(_1628_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6081_ (.I(_0704_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6082_ (.I0(\reg_file.reg_storage[4][18] ),
    .I1(\reg_file.reg_storage[5][18] ),
    .I2(\reg_file.reg_storage[6][18] ),
    .I3(\reg_file.reg_storage[7][18] ),
    .S0(_2212_),
    .S1(_2213_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6083_ (.A1(_1977_),
    .A2(\reg_file.reg_storage[3][18] ),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6084_ (.A1(_2105_),
    .A2(\reg_file.reg_storage[2][18] ),
    .B(_2106_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6085_ (.A1(_1932_),
    .A2(_1194_),
    .B1(_2215_),
    .B2(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6086_ (.I0(\reg_file.reg_storage[12][18] ),
    .I1(\reg_file.reg_storage[13][18] ),
    .I2(\reg_file.reg_storage[14][18] ),
    .I3(\reg_file.reg_storage[15][18] ),
    .S0(_1974_),
    .S1(_1975_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6087_ (.I0(\reg_file.reg_storage[8][18] ),
    .I1(\reg_file.reg_storage[9][18] ),
    .I2(\reg_file.reg_storage[10][18] ),
    .I3(\reg_file.reg_storage[11][18] ),
    .S0(_2212_),
    .S1(_1975_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6088_ (.I0(_2214_),
    .I1(_2217_),
    .I2(_2218_),
    .I3(_2219_),
    .S0(_2113_),
    .S1(_1943_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6089_ (.A1(_1929_),
    .A2(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6090_ (.A1(_2211_),
    .A2(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _6091_ (.A1(_1946_),
    .A2(_1986_),
    .A3(_2036_),
    .A4(_2080_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6092_ (.A1(_2118_),
    .A2(_2180_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6093_ (.A1(_1956_),
    .A2(_2223_),
    .A3(_2224_),
    .B(_0656_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6094_ (.A1(_2222_),
    .A2(_2225_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6095_ (.A1(_2209_),
    .A2(_2226_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6096_ (.I(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6097_ (.A1(_2207_),
    .A2(_2208_),
    .A3(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6098_ (.A1(_2207_),
    .A2(_2208_),
    .B(_2228_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6099_ (.A1(_1325_),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6100_ (.I(_2137_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6101_ (.A1(_1316_),
    .A2(_1852_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6102_ (.A1(_1030_),
    .A2(_1202_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6103_ (.I0(_2140_),
    .I1(_2234_),
    .S(_1352_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6104_ (.A1(_0723_),
    .A2(_2235_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6105_ (.A1(_1583_),
    .A2(_2022_),
    .B(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6106_ (.A1(_1853_),
    .A2(_1849_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6107_ (.A1(_1772_),
    .A2(_2237_),
    .B(_2238_),
    .C(_1562_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6108_ (.A1(_2233_),
    .A2(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6109_ (.A1(_2232_),
    .A2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6110_ (.I(_2222_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6111_ (.A1(_2209_),
    .A2(_2242_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6112_ (.I(_2209_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6113_ (.A1(_2244_),
    .A2(_2242_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6114_ (.A1(_2244_),
    .A2(_2242_),
    .B(_1905_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6115_ (.A1(_2157_),
    .A2(_2245_),
    .B(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6116_ (.A1(_1286_),
    .A2(_2148_),
    .B1(_2243_),
    .B2(_1901_),
    .C(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6117_ (.A1(_2229_),
    .A2(_2231_),
    .B(_2241_),
    .C(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6118_ (.I(_2249_),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6119_ (.I(net11),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6120_ (.A1(_2250_),
    .A2(_2066_),
    .B(_2068_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6121_ (.A1(_2097_),
    .A2(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6122_ (.I0(\reg_file.reg_storage[4][19] ),
    .I1(\reg_file.reg_storage[5][19] ),
    .I2(\reg_file.reg_storage[6][19] ),
    .I3(\reg_file.reg_storage[7][19] ),
    .S0(_2109_),
    .S1(_2213_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6123_ (.A1(_1870_),
    .A2(\reg_file.reg_storage[3][19] ),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6124_ (.A1(_2105_),
    .A2(\reg_file.reg_storage[2][19] ),
    .B(_2106_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6125_ (.A1(_2103_),
    .A2(_1183_),
    .B1(_2254_),
    .B2(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6126_ (.I0(\reg_file.reg_storage[12][19] ),
    .I1(\reg_file.reg_storage[13][19] ),
    .I2(\reg_file.reg_storage[14][19] ),
    .I3(\reg_file.reg_storage[15][19] ),
    .S0(_2212_),
    .S1(_2213_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6127_ (.I0(\reg_file.reg_storage[8][19] ),
    .I1(\reg_file.reg_storage[9][19] ),
    .I2(\reg_file.reg_storage[10][19] ),
    .I3(\reg_file.reg_storage[11][19] ),
    .S0(_2109_),
    .S1(_2213_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6128_ (.I0(_2253_),
    .I1(_2256_),
    .I2(_2257_),
    .I3(_2258_),
    .S0(_2113_),
    .S1(_2114_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6129_ (.A1(_2100_),
    .A2(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6130_ (.A1(_2252_),
    .A2(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6131_ (.I(_2242_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6132_ (.A1(_1670_),
    .A2(_2262_),
    .B(_2225_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6133_ (.A1(_1190_),
    .A2(_2261_),
    .A3(_2263_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6134_ (.I(_2264_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6135_ (.A1(_2244_),
    .A2(_2226_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6136_ (.A1(_2266_),
    .A2(_2230_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6137_ (.A1(_2265_),
    .A2(_2267_),
    .B(_0540_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6138_ (.A1(_2265_),
    .A2(_2267_),
    .B(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6139_ (.A1(_1469_),
    .A2(_1914_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_1421_),
    .A2(_1379_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6141_ (.I0(_2187_),
    .I1(_2271_),
    .S(_0832_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6142_ (.I0(_2061_),
    .I1(_2272_),
    .S(_1503_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6143_ (.I(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6144_ (.A1(_2009_),
    .A2(_1896_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6145_ (.A1(_1609_),
    .A2(_2274_),
    .B(_2275_),
    .C(_1856_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6146_ (.A1(_2270_),
    .A2(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6147_ (.A1(_2139_),
    .A2(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6148_ (.I(_1190_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6149_ (.I(_2261_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6150_ (.I(_2280_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6151_ (.A1(_1191_),
    .A2(_2281_),
    .B(_1706_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6152_ (.A1(_2279_),
    .A2(_2280_),
    .B(_2282_),
    .C(_1456_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6153_ (.A1(_2279_),
    .A2(_2280_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6154_ (.A1(_1405_),
    .A2(_2149_),
    .B1(_2284_),
    .B2(_1532_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6155_ (.A1(_2269_),
    .A2(_2278_),
    .A3(_2283_),
    .A4(_2285_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6156_ (.I(_2286_),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6157_ (.I(_0548_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6158_ (.I(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6159_ (.I(_1872_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6160_ (.A1(net25),
    .A2(_1872_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6161_ (.A1(_2288_),
    .A2(_2289_),
    .B(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6162_ (.A1(_0691_),
    .A2(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6163_ (.I(_1825_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6164_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(\reg_file.reg_storage[5][20] ),
    .I2(\reg_file.reg_storage[6][20] ),
    .I3(\reg_file.reg_storage[7][20] ),
    .S0(_1933_),
    .S1(_2293_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6165_ (.I(_2106_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6166_ (.I(_2212_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6167_ (.A1(_2296_),
    .A2(\reg_file.reg_storage[3][20] ),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6168_ (.A1(_2287_),
    .A2(\reg_file.reg_storage[2][20] ),
    .B(_2072_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6169_ (.A1(_2295_),
    .A2(_1166_),
    .B1(_2297_),
    .B2(_2298_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6170_ (.I(_1869_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6171_ (.I(_1629_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6172_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(\reg_file.reg_storage[13][20] ),
    .I2(\reg_file.reg_storage[14][20] ),
    .I3(\reg_file.reg_storage[15][20] ),
    .S0(_2300_),
    .S1(_2301_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6173_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(\reg_file.reg_storage[9][20] ),
    .I2(\reg_file.reg_storage[10][20] ),
    .I3(\reg_file.reg_storage[11][20] ),
    .S0(_2300_),
    .S1(_2301_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6174_ (.I(_0692_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6175_ (.I0(_2294_),
    .I1(_2299_),
    .I2(_2302_),
    .I3(_2303_),
    .S0(_2304_),
    .S1(_1331_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6176_ (.A1(_1077_),
    .A2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6177_ (.A1(_2292_),
    .A2(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6178_ (.I(_2307_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _6179_ (.A1(_2117_),
    .A2(_2179_),
    .A3(_2222_),
    .A4(_2261_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6180_ (.A1(_1957_),
    .A2(_2223_),
    .A3(_2309_),
    .B(_1796_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6181_ (.A1(_2308_),
    .A2(_2310_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6182_ (.A1(_1176_),
    .A2(_2311_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6183_ (.A1(_2124_),
    .A2(_2184_),
    .A3(_2228_),
    .A4(_2265_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6184_ (.A1(_2227_),
    .A2(_2264_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6185_ (.A1(_2281_),
    .A2(_2263_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6186_ (.A1(_2244_),
    .A2(_2226_),
    .B1(_2315_),
    .B2(_2279_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6187_ (.A1(_2279_),
    .A2(_2315_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _6188_ (.A1(_2205_),
    .A2(_2206_),
    .A3(_2314_),
    .B1(_2316_),
    .B2(_2317_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6189_ (.A1(_2134_),
    .A2(_2313_),
    .B(_2318_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6190_ (.A1(_2312_),
    .A2(_2319_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6191_ (.A1(_2312_),
    .A2(_2319_),
    .B(_0540_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6192_ (.A1(_0723_),
    .A2(_2142_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6193_ (.A1(_1177_),
    .A2(_1192_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6194_ (.I0(_2234_),
    .I1(_2323_),
    .S(_1467_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6195_ (.A1(_1308_),
    .A2(_2324_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6196_ (.A1(_2322_),
    .A2(_2325_),
    .B(_1771_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6197_ (.A1(_1805_),
    .A2(_1921_),
    .B(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6198_ (.A1(_1529_),
    .A2(_1852_),
    .B1(_2327_),
    .B2(_1562_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6199_ (.I(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6200_ (.I(_2137_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6201_ (.A1(_1175_),
    .A2(_2308_),
    .B(_1791_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6202_ (.A1(_1175_),
    .A2(_2308_),
    .B(_1599_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6203_ (.A1(_1174_),
    .A2(_2308_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6204_ (.A1(_1494_),
    .A2(_2148_),
    .B1(_2333_),
    .B2(_1900_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6205_ (.A1(_2331_),
    .A2(_2332_),
    .B(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6206_ (.A1(_2320_),
    .A2(_2321_),
    .B1(_2329_),
    .B2(_2330_),
    .C(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6207_ (.I(_2336_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6208_ (.I(_1162_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6209_ (.I(_2103_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6210_ (.A1(_2338_),
    .A2(_2289_),
    .B(_2290_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6211_ (.A1(_0691_),
    .A2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6212_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(\reg_file.reg_storage[5][21] ),
    .I2(\reg_file.reg_storage[6][21] ),
    .I3(\reg_file.reg_storage[7][21] ),
    .S0(_1933_),
    .S1(_2293_),
    .Z(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6213_ (.A1(_2296_),
    .A2(\reg_file.reg_storage[3][21] ),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6214_ (.A1(_2287_),
    .A2(\reg_file.reg_storage[2][21] ),
    .B(_2072_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6215_ (.A1(_2295_),
    .A2(_1155_),
    .B1(_2342_),
    .B2(_2343_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6216_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(\reg_file.reg_storage[13][21] ),
    .I2(\reg_file.reg_storage[14][21] ),
    .I3(\reg_file.reg_storage[15][21] ),
    .S0(_2300_),
    .S1(_2301_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6217_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(\reg_file.reg_storage[9][21] ),
    .I2(\reg_file.reg_storage[10][21] ),
    .I3(\reg_file.reg_storage[11][21] ),
    .S0(_2300_),
    .S1(_2301_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6218_ (.I0(_2341_),
    .I1(_2344_),
    .I2(_2345_),
    .I3(_2346_),
    .S0(_2304_),
    .S1(_2114_),
    .Z(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6219_ (.A1(_2100_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6220_ (.A1(_2340_),
    .A2(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6221_ (.I(_2349_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6222_ (.I(_1554_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6223_ (.I(_2307_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6224_ (.A1(_2351_),
    .A2(_2352_),
    .B(_2310_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6225_ (.A1(_2337_),
    .A2(_2350_),
    .A3(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6226_ (.A1(_1175_),
    .A2(_2311_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6227_ (.A1(_2355_),
    .A2(_2320_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6228_ (.A1(_2354_),
    .A2(_2356_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6229_ (.A1(_1374_),
    .A2(_1377_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6230_ (.I0(_2271_),
    .I1(_2358_),
    .S(_1768_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6231_ (.I0(_2188_),
    .I1(_2359_),
    .S(_1447_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6232_ (.I0(_1994_),
    .I1(_2360_),
    .S(_1695_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6233_ (.A1(_1593_),
    .A2(_1744_),
    .B1(_2361_),
    .B2(_2007_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6234_ (.I(_2350_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6235_ (.A1(_1373_),
    .A2(_2363_),
    .B(_1705_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6236_ (.A1(_2337_),
    .A2(_2350_),
    .B(_2364_),
    .C(_1762_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6237_ (.A1(_2337_),
    .A2(_2349_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6238_ (.A1(_1531_),
    .A2(_2366_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6239_ (.A1(_2365_),
    .A2(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6240_ (.A1(_1574_),
    .A2(_2149_),
    .B1(_2362_),
    .B2(_2138_),
    .C(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6241_ (.A1(_1866_),
    .A2(_2357_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6242_ (.I(_2370_),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6243_ (.A1(_2350_),
    .A2(_2353_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6244_ (.A1(_1373_),
    .A2(_2371_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6245_ (.A1(_1373_),
    .A2(_2371_),
    .B(_2355_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6246_ (.A1(_2372_),
    .A2(_2373_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6247_ (.A1(_2312_),
    .A2(_2354_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6248_ (.A1(_2319_),
    .A2(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6249_ (.I(_2304_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6250_ (.I(_2290_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6251_ (.A1(_2377_),
    .A2(_2289_),
    .B(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6252_ (.A1(_1328_),
    .A2(_2379_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6253_ (.I(_2296_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6254_ (.I(_2293_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6255_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(\reg_file.reg_storage[5][22] ),
    .I2(\reg_file.reg_storage[6][22] ),
    .I3(\reg_file.reg_storage[7][22] ),
    .S0(_2381_),
    .S1(_2382_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6256_ (.I(_2295_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6257_ (.I(_1628_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_2385_),
    .A2(\reg_file.reg_storage[3][22] ),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6259_ (.A1(_2288_),
    .A2(\reg_file.reg_storage[2][22] ),
    .B(_2338_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6260_ (.A1(_2384_),
    .A2(_1140_),
    .B1(_2386_),
    .B2(_2387_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6261_ (.I(_2293_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6262_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(\reg_file.reg_storage[13][22] ),
    .I2(\reg_file.reg_storage[14][22] ),
    .I3(\reg_file.reg_storage[15][22] ),
    .S0(_1871_),
    .S1(_2389_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6263_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(\reg_file.reg_storage[9][22] ),
    .I2(\reg_file.reg_storage[10][22] ),
    .I3(\reg_file.reg_storage[11][22] ),
    .S0(_1871_),
    .S1(_2389_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6264_ (.I(_2304_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6265_ (.I0(_2383_),
    .I1(_2388_),
    .I2(_2390_),
    .I3(_2391_),
    .S0(_2392_),
    .S1(_1332_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6266_ (.A1(_1078_),
    .A2(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6267_ (.A1(_2380_),
    .A2(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6268_ (.A1(_2307_),
    .A2(_2349_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _6269_ (.A1(_1956_),
    .A2(_2223_),
    .A3(_2309_),
    .A4(_2396_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6270_ (.A1(_0662_),
    .A2(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6271_ (.A1(_2395_),
    .A2(_2398_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6272_ (.A1(_2399_),
    .A2(_1148_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6273_ (.I(_2400_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6274_ (.A1(_2374_),
    .A2(_2376_),
    .A3(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6275_ (.I(_0716_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6276_ (.A1(_2374_),
    .A2(_2376_),
    .B(_2401_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6277_ (.A1(_2403_),
    .A2(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6278_ (.A1(_2402_),
    .A2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6279_ (.A1(_1149_),
    .A2(_1163_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6280_ (.I0(_2323_),
    .I1(_2407_),
    .S(_1352_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6281_ (.I0(_2235_),
    .I1(_2408_),
    .S(_1690_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6282_ (.A1(_1808_),
    .A2(_2409_),
    .B(_1615_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6283_ (.A1(_1696_),
    .A2(_2023_),
    .A3(_2024_),
    .B(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6284_ (.A1(_1659_),
    .A2(_1745_),
    .B(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6285_ (.A1(_2139_),
    .A2(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6286_ (.I(_1147_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6287_ (.A1(_2414_),
    .A2(_2395_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6288_ (.I(_2414_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6289_ (.I(_2395_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6290_ (.A1(_2416_),
    .A2(_2417_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6291_ (.A1(_2416_),
    .A2(_2417_),
    .B(_1762_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6292_ (.A1(_1518_),
    .A2(_2418_),
    .B(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6293_ (.A1(_1623_),
    .A2(_2149_),
    .B1(_2415_),
    .B2(_1597_),
    .C(_2420_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6294_ (.A1(_2406_),
    .A2(_2413_),
    .A3(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6295_ (.I(_2422_),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6296_ (.A1(_0556_),
    .A2(_2289_),
    .B(_2378_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6297_ (.A1(_1329_),
    .A2(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6298_ (.I(_1977_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6299_ (.I(_2425_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6300_ (.I(_2110_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6301_ (.I(_2427_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6302_ (.I0(\reg_file.reg_storage[4][23] ),
    .I1(\reg_file.reg_storage[5][23] ),
    .I2(\reg_file.reg_storage[6][23] ),
    .I3(\reg_file.reg_storage[7][23] ),
    .S0(_2426_),
    .S1(_2428_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6303_ (.I(\reg_file.reg_storage[1][23] ),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6304_ (.I(_2381_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6305_ (.A1(_2431_),
    .A2(\reg_file.reg_storage[3][23] ),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6306_ (.I(_2287_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6307_ (.I(_2295_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6308_ (.A1(_2433_),
    .A2(\reg_file.reg_storage[2][23] ),
    .B(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6309_ (.A1(_2384_),
    .A2(_2430_),
    .B1(_2432_),
    .B2(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6310_ (.I0(\reg_file.reg_storage[12][23] ),
    .I1(\reg_file.reg_storage[13][23] ),
    .I2(\reg_file.reg_storage[14][23] ),
    .I3(\reg_file.reg_storage[15][23] ),
    .S0(_2381_),
    .S1(_2382_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6311_ (.I0(\reg_file.reg_storage[8][23] ),
    .I1(\reg_file.reg_storage[9][23] ),
    .I2(\reg_file.reg_storage[10][23] ),
    .I3(\reg_file.reg_storage[11][23] ),
    .S0(_2381_),
    .S1(_2382_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6312_ (.I0(_2429_),
    .I1(_2436_),
    .I2(_2437_),
    .I3(_2438_),
    .S0(_2392_),
    .S1(_1332_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_1078_),
    .A2(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6314_ (.A1(_2424_),
    .A2(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6315_ (.I(_2441_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6316_ (.A1(_2417_),
    .A2(_2397_),
    .B(_0659_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6317_ (.A1(_2442_),
    .A2(_2443_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6318_ (.A1(_1137_),
    .A2(_2444_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6319_ (.A1(_2416_),
    .A2(_2399_),
    .B(_2404_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6320_ (.A1(_2445_),
    .A2(_2446_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6321_ (.A1(_1414_),
    .A2(_1364_),
    .B(_1370_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6322_ (.I0(_2358_),
    .I1(_2448_),
    .S(_1352_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6323_ (.I0(_2272_),
    .I1(_2449_),
    .S(_1690_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6324_ (.I0(_2062_),
    .I1(_2450_),
    .S(_1572_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _6325_ (.A1(_1711_),
    .A2(_1744_),
    .B1(_2451_),
    .B2(_2007_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6326_ (.A1(_1364_),
    .A2(_2442_),
    .B(_1791_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6327_ (.A1(_1364_),
    .A2(_2442_),
    .B(_1599_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6328_ (.A1(_1363_),
    .A2(_2441_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6329_ (.A1(_1694_),
    .A2(_2147_),
    .B1(_2455_),
    .B2(_1900_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6330_ (.A1(_2453_),
    .A2(_2454_),
    .B(_2456_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6331_ (.A1(_1841_),
    .A2(_2447_),
    .B1(_2452_),
    .B2(_2330_),
    .C(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _6332_ (.I(_2458_),
    .ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6333_ (.A1(net17),
    .A2(_1821_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6334_ (.A1(_2378_),
    .A2(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6335_ (.A1(_1328_),
    .A2(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6336_ (.I0(\reg_file.reg_storage[4][24] ),
    .I1(\reg_file.reg_storage[5][24] ),
    .I2(\reg_file.reg_storage[6][24] ),
    .I3(\reg_file.reg_storage[7][24] ),
    .S0(_1871_),
    .S1(_2389_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6337_ (.I(_2425_),
    .Z(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6338_ (.A1(_2463_),
    .A2(\reg_file.reg_storage[3][24] ),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6339_ (.A1(_2288_),
    .A2(\reg_file.reg_storage[2][24] ),
    .B(_2338_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6340_ (.A1(_2434_),
    .A2(_1110_),
    .B1(_2464_),
    .B2(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6341_ (.I0(\reg_file.reg_storage[12][24] ),
    .I1(\reg_file.reg_storage[13][24] ),
    .I2(\reg_file.reg_storage[14][24] ),
    .I3(\reg_file.reg_storage[15][24] ),
    .S0(_2425_),
    .S1(_2427_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6342_ (.I0(\reg_file.reg_storage[8][24] ),
    .I1(\reg_file.reg_storage[9][24] ),
    .I2(\reg_file.reg_storage[10][24] ),
    .I3(\reg_file.reg_storage[11][24] ),
    .S0(_2425_),
    .S1(_2389_),
    .Z(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6343_ (.I0(_2462_),
    .I1(_2466_),
    .I2(_2467_),
    .I3(_2468_),
    .S0(_2392_),
    .S1(_1331_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6344_ (.A1(_1077_),
    .A2(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6345_ (.A1(_2461_),
    .A2(_2470_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6346_ (.I(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _6347_ (.A1(_2395_),
    .A2(_2397_),
    .A3(_2441_),
    .B(_1836_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6348_ (.A1(_2472_),
    .A2(_2473_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6349_ (.A1(_1118_),
    .A2(_2474_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6350_ (.A1(_2123_),
    .A2(_2184_),
    .A3(_2228_),
    .A4(_2265_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6351_ (.A1(_2476_),
    .A2(_2375_),
    .A3(_2401_),
    .A4(_2445_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _6352_ (.A1(_2127_),
    .A2(_2128_),
    .A3(net103),
    .B(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6353_ (.A1(_2372_),
    .A2(_2373_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6354_ (.A1(_2401_),
    .A2(_2445_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6355_ (.A1(_2375_),
    .A2(_2400_),
    .A3(_2445_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6356_ (.A1(_1363_),
    .A2(_2444_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6357_ (.A1(_2416_),
    .A2(_2399_),
    .B1(_2444_),
    .B2(_1363_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6358_ (.A1(_2482_),
    .A2(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6359_ (.A1(_2479_),
    .A2(_2480_),
    .B1(_2481_),
    .B2(_2318_),
    .C(_2484_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6360_ (.A1(_2478_),
    .A2(_2485_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6361_ (.A1(_2475_),
    .A2(_2486_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6362_ (.A1(_2475_),
    .A2(_2486_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6363_ (.A1(_2487_),
    .A2(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6364_ (.A1(_1606_),
    .A2(_2324_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6365_ (.A1(_1119_),
    .A2(_1138_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6366_ (.I0(_2407_),
    .I1(_2491_),
    .S(_2018_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6367_ (.A1(_1505_),
    .A2(_2492_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6368_ (.A1(_1844_),
    .A2(_2490_),
    .A3(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6369_ (.A1(_1495_),
    .A2(_2143_),
    .B(_2494_),
    .C(_1349_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6370_ (.A1(_1616_),
    .A2(_1756_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6371_ (.A1(_2232_),
    .A2(_2495_),
    .A3(_2496_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6372_ (.A1(_1812_),
    .A2(_0934_),
    .A3(_1743_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6373_ (.I(_2498_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6374_ (.I(_1117_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6375_ (.A1(_2500_),
    .A2(_2472_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6376_ (.I(_2472_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6377_ (.A1(_1118_),
    .A2(_2502_),
    .B(_1705_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6378_ (.A1(_2500_),
    .A2(_2472_),
    .B(_2503_),
    .C(_2159_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6379_ (.A1(_0540_),
    .A2(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6380_ (.A1(_2150_),
    .A2(_2499_),
    .B1(_2501_),
    .B2(_2086_),
    .C(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6381_ (.A1(_1325_),
    .A2(_2489_),
    .B1(_2497_),
    .B2(_2506_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6382_ (.A1(_2500_),
    .A2(_2474_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6383_ (.I(_2290_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6384_ (.I(_1821_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6385_ (.A1(net18),
    .A2(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6386_ (.A1(_2508_),
    .A2(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6387_ (.A1(_1329_),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6388_ (.I(_2427_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6389_ (.I0(\reg_file.reg_storage[4][25] ),
    .I1(\reg_file.reg_storage[5][25] ),
    .I2(\reg_file.reg_storage[6][25] ),
    .I3(\reg_file.reg_storage[7][25] ),
    .S0(_2426_),
    .S1(_2513_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6390_ (.I(_2296_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6391_ (.A1(_2515_),
    .A2(\reg_file.reg_storage[3][25] ),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6392_ (.A1(_2433_),
    .A2(\reg_file.reg_storage[2][25] ),
    .B(_2434_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6393_ (.A1(_2384_),
    .A2(_1097_),
    .B1(_2516_),
    .B2(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6394_ (.I0(\reg_file.reg_storage[12][25] ),
    .I1(\reg_file.reg_storage[13][25] ),
    .I2(\reg_file.reg_storage[14][25] ),
    .I3(\reg_file.reg_storage[15][25] ),
    .S0(_2426_),
    .S1(_2428_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6395_ (.I0(\reg_file.reg_storage[8][25] ),
    .I1(\reg_file.reg_storage[9][25] ),
    .I2(\reg_file.reg_storage[10][25] ),
    .I3(\reg_file.reg_storage[11][25] ),
    .S0(_2426_),
    .S1(_2428_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6396_ (.I0(_2514_),
    .I1(_2518_),
    .I2(_2519_),
    .I3(_2520_),
    .S0(_2392_),
    .S1(_1332_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6397_ (.A1(_1338_),
    .A2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6398_ (.A1(_2512_),
    .A2(_2522_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6399_ (.A1(_2502_),
    .A2(_2473_),
    .B(_2351_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6400_ (.A1(_1107_),
    .A2(_2523_),
    .A3(_2524_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6401_ (.A1(_2507_),
    .A2(_2488_),
    .A3(_2525_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6402_ (.A1(_2507_),
    .A2(_2488_),
    .B(_2525_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6403_ (.A1(_2403_),
    .A2(_2526_),
    .A3(_2527_),
    .Z(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6404_ (.I(_1107_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6405_ (.A1(_1414_),
    .A2(_2529_),
    .B(_1366_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6406_ (.I0(_2448_),
    .I1(_2530_),
    .S(_2018_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6407_ (.I0(_2359_),
    .I1(_2531_),
    .S(_1618_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6408_ (.A1(_1620_),
    .A2(_2190_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6409_ (.A1(_1576_),
    .A2(_2532_),
    .B(_2533_),
    .C(_1510_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6410_ (.A1(_1563_),
    .A2(_1776_),
    .B(_2534_),
    .C(_2232_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6411_ (.A1(_1107_),
    .A2(_2523_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6412_ (.I(_2523_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6413_ (.A1(_2529_),
    .A2(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6414_ (.A1(_2529_),
    .A2(_2537_),
    .B(_1762_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6415_ (.A1(_1706_),
    .A2(_2538_),
    .B(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6416_ (.A1(_1804_),
    .A2(_2499_),
    .B1(_2536_),
    .B2(_1597_),
    .C(_2540_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6417_ (.A1(_2528_),
    .A2(_2535_),
    .A3(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6418_ (.I(_2542_),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6419_ (.A1(_2475_),
    .A2(_2525_),
    .Z(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6420_ (.A1(_2537_),
    .A2(_2524_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6421_ (.A1(_1356_),
    .A2(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6422_ (.A1(_1356_),
    .A2(_2544_),
    .B(_2507_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6423_ (.A1(_2545_),
    .A2(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6424_ (.A1(_2486_),
    .A2(_2543_),
    .B(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6425_ (.A1(net19),
    .A2(_2509_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6426_ (.A1(_2508_),
    .A2(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6427_ (.A1(_1329_),
    .A2(_2550_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6428_ (.I0(\reg_file.reg_storage[4][26] ),
    .I1(\reg_file.reg_storage[5][26] ),
    .I2(\reg_file.reg_storage[6][26] ),
    .I3(\reg_file.reg_storage[7][26] ),
    .S0(_2385_),
    .S1(_2513_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6429_ (.I(_2338_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6430_ (.A1(_2515_),
    .A2(\reg_file.reg_storage[3][26] ),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6431_ (.A1(_2433_),
    .A2(\reg_file.reg_storage[2][26] ),
    .B(_2434_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6432_ (.A1(_2553_),
    .A2(_1249_),
    .B1(_2554_),
    .B2(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6433_ (.I0(\reg_file.reg_storage[12][26] ),
    .I1(\reg_file.reg_storage[13][26] ),
    .I2(\reg_file.reg_storage[14][26] ),
    .I3(\reg_file.reg_storage[15][26] ),
    .S0(_2463_),
    .S1(_2513_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6434_ (.I0(\reg_file.reg_storage[8][26] ),
    .I1(\reg_file.reg_storage[9][26] ),
    .I2(\reg_file.reg_storage[10][26] ),
    .I3(\reg_file.reg_storage[11][26] ),
    .S0(_2463_),
    .S1(_2513_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6435_ (.I0(_2552_),
    .I1(_2556_),
    .I2(_2557_),
    .I3(_2558_),
    .S0(_2377_),
    .S1(_1335_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6436_ (.A1(_1338_),
    .A2(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6437_ (.A1(_2551_),
    .A2(_2560_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6438_ (.I(_2561_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6439_ (.A1(_2471_),
    .A2(_2523_),
    .B(_1796_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6440_ (.A1(_2473_),
    .A2(_2563_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6441_ (.A1(_2562_),
    .A2(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6442_ (.A1(_1256_),
    .A2(_2565_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6443_ (.I(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6444_ (.A1(_2548_),
    .A2(_2567_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6445_ (.A1(_2548_),
    .A2(_2567_),
    .B(_2044_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6446_ (.A1(_1616_),
    .A2(_1851_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6447_ (.A1(_1411_),
    .A2(_2529_),
    .B(_1257_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6448_ (.I0(_2491_),
    .I1(_2571_),
    .S(_1353_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6449_ (.I0(_2408_),
    .I1(_2572_),
    .S(_1583_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6450_ (.A1(_1620_),
    .A2(_2237_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6451_ (.A1(_1576_),
    .A2(_2573_),
    .B(_2574_),
    .C(_1349_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6452_ (.A1(_2232_),
    .A2(_2570_),
    .A3(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6453_ (.I(_2498_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6454_ (.I(_2561_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6455_ (.A1(_1359_),
    .A2(_2578_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6456_ (.A1(_1360_),
    .A2(_2578_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6457_ (.A1(_1360_),
    .A2(_2578_),
    .B(_2159_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6458_ (.A1(_2157_),
    .A2(_2580_),
    .B(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6459_ (.A1(_1284_),
    .A2(_2577_),
    .B1(_2579_),
    .B2(_2086_),
    .C(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6460_ (.A1(_2568_),
    .A2(_2569_),
    .B(_2576_),
    .C(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6461_ (.I(_2584_),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6462_ (.I(_1328_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6463_ (.I(_2378_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6464_ (.I(_1821_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6465_ (.A1(net20),
    .A2(_2587_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6466_ (.A1(_2586_),
    .A2(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6467_ (.A1(_2585_),
    .A2(_2589_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6468_ (.I(_1078_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6469_ (.I(_2385_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6470_ (.I(_2382_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6471_ (.I0(\reg_file.reg_storage[4][27] ),
    .I1(\reg_file.reg_storage[5][27] ),
    .I2(\reg_file.reg_storage[6][27] ),
    .I3(\reg_file.reg_storage[7][27] ),
    .S0(_2592_),
    .S1(_2593_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6472_ (.I(_2384_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6473_ (.I(_2515_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6474_ (.A1(_2596_),
    .A2(\reg_file.reg_storage[3][27] ),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6475_ (.I(_2288_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6476_ (.A1(_2598_),
    .A2(\reg_file.reg_storage[2][27] ),
    .B(_2553_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6477_ (.A1(_2595_),
    .A2(_1239_),
    .B1(_2597_),
    .B2(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6478_ (.I0(\reg_file.reg_storage[12][27] ),
    .I1(\reg_file.reg_storage[13][27] ),
    .I2(\reg_file.reg_storage[14][27] ),
    .I3(\reg_file.reg_storage[15][27] ),
    .S0(_2515_),
    .S1(_2593_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6479_ (.I0(\reg_file.reg_storage[8][27] ),
    .I1(\reg_file.reg_storage[9][27] ),
    .I2(\reg_file.reg_storage[10][27] ),
    .I3(\reg_file.reg_storage[11][27] ),
    .S0(_2592_),
    .S1(_2593_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6480_ (.I(_2377_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6481_ (.I0(_2594_),
    .I1(_2600_),
    .I2(_2601_),
    .I3(_2602_),
    .S0(_2603_),
    .S1(_1335_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6482_ (.A1(_2591_),
    .A2(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6483_ (.A1(_2590_),
    .A2(_2605_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6484_ (.A1(_2351_),
    .A2(_2562_),
    .B(_2563_),
    .C(_2473_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6485_ (.A1(_2606_),
    .A2(_2607_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6486_ (.A1(_1246_),
    .A2(_2608_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6487_ (.A1(_1360_),
    .A2(_2565_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6488_ (.A1(_2610_),
    .A2(_2568_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6489_ (.A1(_2609_),
    .A2(_2611_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6490_ (.A1(_2609_),
    .A2(_2611_),
    .B(_2403_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6491_ (.I(_2606_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6492_ (.A1(_1393_),
    .A2(_2614_),
    .B(_1791_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6493_ (.A1(_1393_),
    .A2(_2614_),
    .B(_1456_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6494_ (.A1(_1247_),
    .A2(_2606_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6495_ (.A1(_1403_),
    .A2(_2577_),
    .B1(_2617_),
    .B2(_1531_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6496_ (.A1(_1394_),
    .A2(_1361_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6497_ (.A1(_1387_),
    .A2(_2530_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6498_ (.A1(_1438_),
    .A2(_2619_),
    .B(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6499_ (.I0(_2449_),
    .I1(_2621_),
    .S(_1848_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6500_ (.A1(_1771_),
    .A2(_2274_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6501_ (.A1(_1384_),
    .A2(_2622_),
    .B(_2623_),
    .C(_1348_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6502_ (.A1(_1856_),
    .A2(_1898_),
    .B(_2624_),
    .C(_2137_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6503_ (.A1(_2615_),
    .A2(_2616_),
    .B(_2618_),
    .C(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6504_ (.A1(_2612_),
    .A2(_2613_),
    .B(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6505_ (.I(_2627_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6506_ (.A1(_1355_),
    .A2(_1246_),
    .B(_1236_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6507_ (.A1(_1402_),
    .A2(_2571_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6508_ (.A1(_1773_),
    .A2(_2628_),
    .B(_2629_),
    .C(_1498_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6509_ (.A1(_1505_),
    .A2(_2492_),
    .B(_2630_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6510_ (.A1(_1696_),
    .A2(_2631_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6511_ (.A1(_1772_),
    .A2(_2322_),
    .A3(_2325_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6512_ (.A1(_1517_),
    .A2(_2632_),
    .A3(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6513_ (.A1(_1563_),
    .A2(_1923_),
    .B(_2634_),
    .C(_2330_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6514_ (.A1(net21),
    .A2(_2509_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6515_ (.A1(_2508_),
    .A2(_2636_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6516_ (.A1(_2585_),
    .A2(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6517_ (.I(_2385_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6518_ (.I(_2428_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6519_ (.I0(\reg_file.reg_storage[4][28] ),
    .I1(\reg_file.reg_storage[5][28] ),
    .I2(\reg_file.reg_storage[6][28] ),
    .I3(\reg_file.reg_storage[7][28] ),
    .S0(_2639_),
    .S1(_2640_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6520_ (.I(_2553_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6521_ (.I(_2463_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6522_ (.A1(_2643_),
    .A2(\reg_file.reg_storage[3][28] ),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6523_ (.A1(_2598_),
    .A2(\reg_file.reg_storage[2][28] ),
    .B(_2595_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6524_ (.A1(_2642_),
    .A2(_1230_),
    .B1(_2644_),
    .B2(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6525_ (.I0(\reg_file.reg_storage[12][28] ),
    .I1(\reg_file.reg_storage[13][28] ),
    .I2(\reg_file.reg_storage[14][28] ),
    .I3(\reg_file.reg_storage[15][28] ),
    .S0(_2592_),
    .S1(_2593_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6526_ (.I0(\reg_file.reg_storage[8][28] ),
    .I1(\reg_file.reg_storage[9][28] ),
    .I2(\reg_file.reg_storage[10][28] ),
    .I3(\reg_file.reg_storage[11][28] ),
    .S0(_2592_),
    .S1(_2640_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6527_ (.I0(_2641_),
    .I1(_2646_),
    .I2(_2647_),
    .I3(_2648_),
    .S0(_2603_),
    .S1(_1333_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6528_ (.A1(_2591_),
    .A2(_2649_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6529_ (.A1(_2638_),
    .A2(_2650_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6530_ (.A1(_1235_),
    .A2(_2651_),
    .Z(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6531_ (.I(_1235_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6532_ (.I(_2651_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6533_ (.A1(_2653_),
    .A2(_2654_),
    .B(_1661_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6534_ (.A1(_2653_),
    .A2(_2654_),
    .B(_1599_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6535_ (.A1(_2655_),
    .A2(_2656_),
    .B(_0716_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6536_ (.A1(_1492_),
    .A2(_2499_),
    .B1(_2652_),
    .B2(_1597_),
    .C(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6537_ (.A1(_1247_),
    .A2(_2608_),
    .B(_2610_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6538_ (.A1(_1393_),
    .A2(_2608_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6539_ (.A1(_2547_),
    .A2(_2566_),
    .A3(_2609_),
    .B1(_2659_),
    .B2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6540_ (.A1(_2543_),
    .A2(_2566_),
    .A3(_2609_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6541_ (.A1(_2478_),
    .A2(_2485_),
    .B(_2662_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6542_ (.A1(_2182_),
    .A2(_2614_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6543_ (.A1(_2607_),
    .A2(_2664_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6544_ (.A1(_2654_),
    .A2(_2665_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6545_ (.A1(_2653_),
    .A2(_2666_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6546_ (.A1(_2661_),
    .A2(_2663_),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6547_ (.A1(_2667_),
    .A2(_2661_),
    .A3(_2663_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6548_ (.A1(_2668_),
    .A2(_2669_),
    .B(_2403_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6549_ (.A1(_2635_),
    .A2(_2658_),
    .B(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6550_ (.I(_2671_),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6551_ (.I(_1218_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6552_ (.A1(_1411_),
    .A2(_2672_),
    .B(_1391_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6553_ (.A1(_1577_),
    .A2(_2673_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6554_ (.A1(_1402_),
    .A2(_2619_),
    .B(_2674_),
    .C(_2017_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6555_ (.A1(_1606_),
    .A2(_2531_),
    .B(_2675_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6556_ (.A1(_1853_),
    .A2(_2360_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6557_ (.A1(_1772_),
    .A2(_2676_),
    .B(_2677_),
    .C(_1562_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6558_ (.A1(_2007_),
    .A2(_1996_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6559_ (.A1(_2678_),
    .A2(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6560_ (.I(_2577_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6561_ (.A1(net22),
    .A2(_2509_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6562_ (.A1(_2508_),
    .A2(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6563_ (.A1(_2585_),
    .A2(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6564_ (.I(_2427_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6565_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(\reg_file.reg_storage[5][29] ),
    .I2(\reg_file.reg_storage[6][29] ),
    .I3(\reg_file.reg_storage[7][29] ),
    .S0(_2431_),
    .S1(_2685_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6566_ (.A1(_2639_),
    .A2(\reg_file.reg_storage[3][29] ),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6567_ (.A1(_2433_),
    .A2(\reg_file.reg_storage[2][29] ),
    .B(_2553_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6568_ (.A1(_2595_),
    .A2(_1210_),
    .B1(_2687_),
    .B2(_2688_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6569_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(\reg_file.reg_storage[13][29] ),
    .I2(\reg_file.reg_storage[14][29] ),
    .I3(\reg_file.reg_storage[15][29] ),
    .S0(_2431_),
    .S1(_2685_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6570_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(\reg_file.reg_storage[9][29] ),
    .I2(\reg_file.reg_storage[10][29] ),
    .I3(\reg_file.reg_storage[11][29] ),
    .S0(_2431_),
    .S1(_2685_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6571_ (.I0(_2686_),
    .I1(_2689_),
    .I2(_2690_),
    .I3(_2691_),
    .S0(_2377_),
    .S1(_1335_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6572_ (.A1(_1338_),
    .A2(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6573_ (.A1(_2684_),
    .A2(_2693_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6574_ (.A1(_1217_),
    .A2(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6575_ (.I(_2694_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6576_ (.A1(_1217_),
    .A2(_2696_),
    .B(_1292_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6577_ (.A1(_2672_),
    .A2(_2694_),
    .B(_2697_),
    .C(_1300_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6578_ (.A1(_1566_),
    .A2(_2681_),
    .B1(_2695_),
    .B2(_1663_),
    .C(_2698_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6579_ (.A1(_2653_),
    .A2(_2666_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6580_ (.A1(_2700_),
    .A2(_2668_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6581_ (.A1(_2182_),
    .A2(_2651_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6582_ (.A1(_2607_),
    .A2(_2664_),
    .A3(_2702_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6583_ (.A1(_2696_),
    .A2(_2703_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6584_ (.A1(_2672_),
    .A2(_2704_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6585_ (.A1(_2672_),
    .A2(_2704_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6586_ (.A1(_2705_),
    .A2(_2706_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6587_ (.A1(_2701_),
    .A2(_2707_),
    .B(_1324_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6588_ (.A1(_2701_),
    .A2(_2707_),
    .B(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6589_ (.A1(_2330_),
    .A2(_2680_),
    .B(_2699_),
    .C(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6590_ (.I(_2710_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6591_ (.I(_2700_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6592_ (.I(_2706_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6593_ (.A1(_2711_),
    .A2(_2705_),
    .B(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6594_ (.A1(_2661_),
    .A2(_2663_),
    .B(_2707_),
    .C(_2667_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6595_ (.A1(_1298_),
    .A2(_2587_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6596_ (.A1(_2586_),
    .A2(_2715_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6597_ (.I(_2685_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6598_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(\reg_file.reg_storage[5][30] ),
    .I2(\reg_file.reg_storage[6][30] ),
    .I3(\reg_file.reg_storage[7][30] ),
    .S0(_2596_),
    .S1(_2717_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_2643_),
    .A2(\reg_file.reg_storage[3][30] ),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6600_ (.A1(_2598_),
    .A2(\reg_file.reg_storage[2][30] ),
    .B(_2595_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6601_ (.A1(_2642_),
    .A2(_1262_),
    .B1(_2719_),
    .B2(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6602_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(\reg_file.reg_storage[13][30] ),
    .I2(\reg_file.reg_storage[14][30] ),
    .I3(\reg_file.reg_storage[15][30] ),
    .S0(_2639_),
    .S1(_2640_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6603_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(\reg_file.reg_storage[9][30] ),
    .I2(\reg_file.reg_storage[10][30] ),
    .I3(\reg_file.reg_storage[11][30] ),
    .S0(_2639_),
    .S1(_2640_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6604_ (.I0(_2718_),
    .I1(_2721_),
    .I2(_2722_),
    .I3(_2723_),
    .S0(_2603_),
    .S1(_1333_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6605_ (.A1(_2591_),
    .A2(_2724_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6606_ (.A1(_0698_),
    .A2(_2716_),
    .B(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6607_ (.I(_2726_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6608_ (.A1(_2182_),
    .A2(_2694_),
    .B(_2703_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6609_ (.A1(_2727_),
    .A2(_2728_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6610_ (.A1(_1269_),
    .A2(_2729_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6611_ (.A1(_2713_),
    .A2(_2714_),
    .A3(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6612_ (.A1(_2713_),
    .A2(_2714_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6613_ (.I(_2730_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6614_ (.A1(_2733_),
    .A2(_2732_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6615_ (.A1(_1841_),
    .A2(_2731_),
    .A3(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6616_ (.A1(_1387_),
    .A2(_1219_),
    .A3(_1271_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6617_ (.A1(_1577_),
    .A2(_2628_),
    .B(_2736_),
    .C(_1397_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6618_ (.A1(_2017_),
    .A2(_2572_),
    .B(_2737_),
    .C(_1771_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6619_ (.A1(_1572_),
    .A2(_2409_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6620_ (.A1(_1615_),
    .A2(_2738_),
    .A3(_2739_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6621_ (.A1(_1517_),
    .A2(_2026_),
    .B(_2740_),
    .C(_2138_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6622_ (.I(_2727_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6623_ (.A1(_1269_),
    .A2(_2742_),
    .B(_1902_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6624_ (.A1(_1388_),
    .A2(_2727_),
    .B(_2743_),
    .C(_1456_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6625_ (.A1(_1270_),
    .A2(_2726_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6626_ (.A1(_1621_),
    .A2(_2577_),
    .B1(_2745_),
    .B2(_1471_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6627_ (.A1(_2735_),
    .A2(_2741_),
    .A3(_2744_),
    .A4(_2746_),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6628_ (.I(_2747_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6629_ (.A1(_1388_),
    .A2(_2729_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6630_ (.A1(_2734_),
    .A2(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6631_ (.A1(_1874_),
    .A2(_2585_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6632_ (.I0(\reg_file.reg_storage[4][31] ),
    .I1(\reg_file.reg_storage[5][31] ),
    .I2(\reg_file.reg_storage[6][31] ),
    .I3(\reg_file.reg_storage[7][31] ),
    .S0(_2643_),
    .S1(_2717_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6633_ (.A1(_2643_),
    .A2(\reg_file.reg_storage[3][31] ),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6634_ (.A1(_2598_),
    .A2(\reg_file.reg_storage[2][31] ),
    .B(_2642_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6635_ (.A1(_2642_),
    .A2(_1273_),
    .B1(_2752_),
    .B2(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6636_ (.I0(\reg_file.reg_storage[12][31] ),
    .I1(\reg_file.reg_storage[13][31] ),
    .I2(\reg_file.reg_storage[14][31] ),
    .I3(\reg_file.reg_storage[15][31] ),
    .S0(_2596_),
    .S1(_2717_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6637_ (.I0(\reg_file.reg_storage[8][31] ),
    .I1(\reg_file.reg_storage[9][31] ),
    .I2(\reg_file.reg_storage[10][31] ),
    .I3(\reg_file.reg_storage[11][31] ),
    .S0(_2596_),
    .S1(_2717_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6638_ (.I0(_2751_),
    .I1(_2754_),
    .I2(_2755_),
    .I3(_2756_),
    .S0(_2603_),
    .S1(_1333_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6639_ (.A1(_2591_),
    .A2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6640_ (.A1(_2750_),
    .A2(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6641_ (.A1(_1280_),
    .A2(_2759_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6642_ (.A1(_2742_),
    .A2(_2728_),
    .B(_2351_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6643_ (.A1(_2749_),
    .A2(_2760_),
    .A3(_2761_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6644_ (.A1(_1355_),
    .A2(_1388_),
    .B(_1399_),
    .C(_1401_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6645_ (.A1(_1577_),
    .A2(_2673_),
    .B(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6646_ (.A1(_1385_),
    .A2(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6647_ (.A1(_1522_),
    .A2(_2621_),
    .B(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6648_ (.A1(_1486_),
    .A2(_2450_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6649_ (.A1(_2009_),
    .A2(_2766_),
    .B(_2767_),
    .C(_1451_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6650_ (.A1(_1510_),
    .A2(_2064_),
    .B(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6651_ (.A1(_0523_),
    .A2(_2760_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6652_ (.A1(_2750_),
    .A2(_2758_),
    .B(_0537_),
    .C(_1398_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6653_ (.A1(_2770_),
    .A2(_2771_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _6654_ (.A1(_2138_),
    .A2(_2769_),
    .B1(_2772_),
    .B2(_1662_),
    .C1(_1692_),
    .C2(_2499_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6655_ (.A1(_1866_),
    .A2(_2762_),
    .B(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6656_ (.I(_2774_),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6657_ (.A1(_0531_),
    .A2(_0507_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6658_ (.A1(_2333_),
    .A2(_2366_),
    .A3(_2415_),
    .A4(_2455_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6659_ (.A1(_2156_),
    .A2(_2197_),
    .A3(_2243_),
    .A4(_2284_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6660_ (.A1(_2501_),
    .A2(_2536_),
    .A3(_2579_),
    .A4(_2617_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6661_ (.I(_2652_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6662_ (.A1(_2779_),
    .A2(_2695_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6663_ (.A1(_2745_),
    .A2(_2760_),
    .A3(_2780_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6664_ (.A1(_2776_),
    .A2(_2777_),
    .A3(_2778_),
    .A4(_2781_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _6665_ (.A1(_1949_),
    .A2(_1998_),
    .A3(_2039_),
    .A4(_2085_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6666_ (.A1(_1758_),
    .A2(_1794_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6667_ (.A1(_1862_),
    .A2(_1899_),
    .A3(_2783_),
    .A4(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6668_ (.A1(_0666_),
    .A2(_0830_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6669_ (.I(_1660_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6670_ (.A1(_1462_),
    .A2(_1313_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6671_ (.A1(_2787_),
    .A2(_1713_),
    .A3(_2788_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6672_ (.A1(_1317_),
    .A2(_1470_),
    .A3(_1530_),
    .A4(_1596_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6673_ (.A1(_2785_),
    .A2(_2786_),
    .A3(_2789_),
    .A4(_2790_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6674_ (.A1(_2782_),
    .A2(_2791_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6675_ (.I(_1530_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6676_ (.A1(_0829_),
    .A2(_1313_),
    .B(_0665_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6677_ (.A1(_0828_),
    .A2(_1312_),
    .B1(_1296_),
    .B2(_1301_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6678_ (.A1(_0883_),
    .A2(_0719_),
    .B1(_2794_),
    .B2(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6679_ (.A1(net105),
    .A2(_0895_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6680_ (.A1(_1470_),
    .A2(_2796_),
    .B(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6681_ (.A1(_0876_),
    .A2(_1613_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6682_ (.A1(_2793_),
    .A2(_2798_),
    .B(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6683_ (.A1(_0857_),
    .A2(_1595_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6684_ (.A1(_1596_),
    .A2(_2800_),
    .B(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6685_ (.A1(_1626_),
    .A2(_1640_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6686_ (.A1(_1660_),
    .A2(_2802_),
    .B(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6687_ (.A1(_0809_),
    .A2(_1680_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6688_ (.A1(_1713_),
    .A2(_2804_),
    .B(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6689_ (.A1(_0745_),
    .A2(_1790_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6690_ (.A1(_0782_),
    .A2(_1757_),
    .A3(_1794_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6691_ (.A1(_2807_),
    .A2(_2808_),
    .B(_1862_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6692_ (.A1(_1013_),
    .A2(_1831_),
    .B(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6693_ (.A1(_1899_),
    .A2(_2810_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6694_ (.A1(_0989_),
    .A2(_1886_),
    .B(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6695_ (.A1(_0959_),
    .A2(_1988_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6696_ (.A1(_0975_),
    .A2(_1948_),
    .A3(_1997_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6697_ (.A1(_2813_),
    .A2(_2814_),
    .B(_2039_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6698_ (.A1(_1417_),
    .A2(_2038_),
    .B(_2815_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6699_ (.A1(_1070_),
    .A2(_2081_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6700_ (.A1(_2783_),
    .A2(_2812_),
    .B1(_2816_),
    .B2(_2085_),
    .C(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6701_ (.A1(_2785_),
    .A2(_2806_),
    .B(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6702_ (.I(_2778_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6703_ (.I(_2243_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6704_ (.A1(_1043_),
    .A2(_2118_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6705_ (.A1(_1029_),
    .A2(_2180_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6706_ (.A1(_2197_),
    .A2(_2822_),
    .B(_2823_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6707_ (.A1(_2209_),
    .A2(_2262_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6708_ (.A1(_2821_),
    .A2(_2824_),
    .B(_2825_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6709_ (.A1(_1191_),
    .A2(_2280_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6710_ (.A1(_2284_),
    .A2(_2826_),
    .B(_2827_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6711_ (.A1(_1148_),
    .A2(_2417_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6712_ (.I(_2415_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6713_ (.A1(_1174_),
    .A2(_2352_),
    .A3(_2366_),
    .B1(_2363_),
    .B2(_2337_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6714_ (.A1(_2830_),
    .A2(_2831_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6715_ (.A1(_2829_),
    .A2(_2832_),
    .B(_2455_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6716_ (.A1(_1137_),
    .A2(_2442_),
    .B1(_2776_),
    .B2(_2828_),
    .C(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6717_ (.A1(_1356_),
    .A2(_2537_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6718_ (.A1(_2500_),
    .A2(_2502_),
    .A3(_2536_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6719_ (.A1(_2835_),
    .A2(_2836_),
    .B(_2579_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6720_ (.A1(_1256_),
    .A2(_2578_),
    .B(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6721_ (.A1(_1246_),
    .A2(_2614_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6722_ (.A1(_2820_),
    .A2(_2834_),
    .B1(_2838_),
    .B2(_2617_),
    .C(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6723_ (.A1(_1269_),
    .A2(_2727_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6724_ (.I(_2745_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6725_ (.A1(_2654_),
    .A2(_2695_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6726_ (.A1(_1218_),
    .A2(_2696_),
    .B1(_2843_),
    .B2(_1235_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6727_ (.A1(_2842_),
    .A2(_2844_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6728_ (.A1(_2841_),
    .A2(_2845_),
    .B(_2760_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6729_ (.A1(_1280_),
    .A2(_2759_),
    .B1(_2781_),
    .B2(_2840_),
    .C(_2846_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6730_ (.A1(_2782_),
    .A2(_2819_),
    .B(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6731_ (.A1(_2770_),
    .A2(_2848_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6732_ (.A1(_0533_),
    .A2(_2775_),
    .A3(_2792_),
    .A4(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6733_ (.A1(_0882_),
    .A2(_0607_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6734_ (.A1(_1151_),
    .A2(_1310_),
    .A3(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6735_ (.A1(_0831_),
    .A2(_0898_),
    .B(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6736_ (.A1(_0721_),
    .A2(_1507_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6737_ (.A1(_0900_),
    .A2(_2853_),
    .B(_2854_),
    .C(_1406_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6738_ (.A1(_1407_),
    .A2(_1747_),
    .B(_2855_),
    .C(_1092_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6739_ (.A1(_1614_),
    .A2(_2152_),
    .B(_0538_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6740_ (.A1(_0534_),
    .A2(_2792_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6741_ (.A1(_1378_),
    .A2(_0607_),
    .B(_1291_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6742_ (.A1(_1299_),
    .A2(_2851_),
    .A3(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6743_ (.A1(_1318_),
    .A2(_2788_),
    .B(_1323_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6744_ (.A1(_1655_),
    .A2(_1755_),
    .B(_2860_),
    .C(_2861_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6745_ (.A1(_2856_),
    .A2(_2857_),
    .B(_2858_),
    .C(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6746_ (.A1(_0539_),
    .A2(_2788_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6747_ (.A1(_2850_),
    .A2(_2863_),
    .B(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6748_ (.I(_2865_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6749_ (.A1(_1402_),
    .A2(_1463_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6750_ (.A1(_1773_),
    .A2(_1442_),
    .B1(_1465_),
    .B2(_2866_),
    .C(_2017_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6751_ (.A1(_1606_),
    .A2(_1578_),
    .B(_2867_),
    .C(_2009_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6752_ (.A1(_1844_),
    .A2(_1809_),
    .B(_1451_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6753_ (.A1(_1517_),
    .A2(_2196_),
    .B1(_2868_),
    .B2(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6754_ (.A1(_1858_),
    .A2(_2870_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6755_ (.A1(_1307_),
    .A2(_1774_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6756_ (.A1(_0636_),
    .A2(_2018_),
    .B(_1457_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6757_ (.A1(_0666_),
    .A2(_1773_),
    .B(_1515_),
    .C(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6758_ (.A1(_1664_),
    .A2(_2786_),
    .B(_2872_),
    .C(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6759_ (.A1(_1462_),
    .A2(_0658_),
    .B(_1841_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6760_ (.A1(_1462_),
    .A2(_0658_),
    .B(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6761_ (.A1(_2871_),
    .A2(_2875_),
    .A3(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6762_ (.I(_2878_),
    .ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6763_ (.I(_0669_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6764_ (.A1(net12),
    .A2(net1),
    .A3(_0511_),
    .A4(_0512_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6765_ (.A1(_0491_),
    .A2(_0511_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6766_ (.A1(_0535_),
    .A2(net65),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6767_ (.A1(_0489_),
    .A2(_2881_),
    .B1(_2882_),
    .B2(_0530_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6768_ (.A1(net12),
    .A2(net1),
    .A3(_2883_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6769_ (.A1(_2880_),
    .A2(_2884_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6770_ (.I(_2885_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6771_ (.I(_2886_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6772_ (.A1(net12),
    .A2(net1),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6773_ (.A1(_0582_),
    .A2(_0492_),
    .A3(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6774_ (.I(_2889_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6775_ (.I(_2890_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6776_ (.A1(net12),
    .A2(net1),
    .A3(_2883_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6777_ (.I(_2892_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6778_ (.I(_2893_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6779_ (.I(_0695_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6780_ (.I(\pc[0] ),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6781_ (.A1(_2896_),
    .A2(_0554_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6782_ (.A1(_0664_),
    .A2(_0642_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6783_ (.A1(_0664_),
    .A2(_0642_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6784_ (.A1(_2897_),
    .A2(_2898_),
    .B(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6785_ (.A1(_1293_),
    .A2(_2895_),
    .A3(_2900_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6786_ (.A1(net87),
    .A2(_2891_),
    .B1(_2894_),
    .B2(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6787_ (.A1(_2879_),
    .A2(_2887_),
    .B(_2902_),
    .ZN(\pc_next[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6788_ (.I(\pc[3] ),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6789_ (.A1(_1293_),
    .A2(_2903_),
    .Z(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6790_ (.I(_2892_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6791_ (.I(_2905_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6792_ (.I(_1330_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6793_ (.A1(_0669_),
    .A2(_2895_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6794_ (.A1(_2879_),
    .A2(_2895_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6795_ (.A1(_2908_),
    .A2(_2900_),
    .B(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6796_ (.A1(_2903_),
    .A2(_2907_),
    .A3(_2910_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6797_ (.A1(net90),
    .A2(_2891_),
    .B1(_2906_),
    .B2(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6798_ (.A1(_2887_),
    .A2(_2904_),
    .B(_2912_),
    .ZN(\pc_next[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6799_ (.A1(\pc[2] ),
    .A2(\pc[3] ),
    .A3(\pc[4] ),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6800_ (.I(\pc[4] ),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6801_ (.A1(_2879_),
    .A2(_2903_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6802_ (.A1(_2914_),
    .A2(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6803_ (.A1(_2913_),
    .A2(_2916_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6804_ (.I(_2890_),
    .Z(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6805_ (.A1(_2914_),
    .A2(_1089_),
    .Z(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6806_ (.A1(_2914_),
    .A2(_1089_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6807_ (.A1(_2919_),
    .A2(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6808_ (.A1(\pc[3] ),
    .A2(_2907_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6809_ (.A1(_2903_),
    .A2(_2907_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6810_ (.A1(_2922_),
    .A2(_2910_),
    .B(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6811_ (.A1(_2921_),
    .A2(_2924_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6812_ (.A1(net91),
    .A2(_2918_),
    .B1(_2906_),
    .B2(_2925_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6813_ (.A1(_2887_),
    .A2(_2917_),
    .B(_2926_),
    .ZN(\pc_next[4] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6814_ (.I(_2885_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6815_ (.I(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6816_ (.I(\pc[5] ),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6817_ (.A1(_2929_),
    .A2(_2913_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6818_ (.A1(_2929_),
    .A2(_1539_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6819_ (.A1(_2921_),
    .A2(_2924_),
    .B(_2919_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6820_ (.I(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6821_ (.A1(_2931_),
    .A2(_2933_),
    .Z(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6822_ (.A1(net92),
    .A2(_2918_),
    .B1(_2906_),
    .B2(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6823_ (.A1(_2928_),
    .A2(_2930_),
    .B(_2935_),
    .ZN(\pc_next[5] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6824_ (.I(\pc[5] ),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6825_ (.A1(_2936_),
    .A2(_2913_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6826_ (.A1(_0812_),
    .A2(_2937_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6827_ (.I(_2587_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6828_ (.A1(_2929_),
    .A2(net18),
    .A3(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6829_ (.A1(net18),
    .A2(_2587_),
    .B(_2929_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6830_ (.A1(_2940_),
    .A2(_2933_),
    .B(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6831_ (.A1(\pc[6] ),
    .A2(_1627_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6832_ (.A1(_2942_),
    .A2(_2943_),
    .Z(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6833_ (.A1(net93),
    .A2(_2918_),
    .B1(_2906_),
    .B2(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6834_ (.A1(_2928_),
    .A2(_2938_),
    .B(_2945_),
    .ZN(\pc_next[6] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6835_ (.A1(_0787_),
    .A2(\pc[6] ),
    .A3(_2937_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6836_ (.A1(_0812_),
    .A2(_2937_),
    .B(_0787_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6837_ (.A1(_2946_),
    .A2(_2947_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6838_ (.I(_2905_),
    .Z(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6839_ (.I(\pc[7] ),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6840_ (.A1(_2950_),
    .A2(_1671_),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6841_ (.A1(_0812_),
    .A2(net19),
    .A3(_2939_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6842_ (.A1(_2942_),
    .A2(_2943_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6843_ (.A1(_2952_),
    .A2(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6844_ (.A1(_2951_),
    .A2(_2954_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6845_ (.A1(net94),
    .A2(_2918_),
    .B1(_2949_),
    .B2(_2955_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6846_ (.A1(_2928_),
    .A2(_2948_),
    .B(_2956_),
    .ZN(\pc_next[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6847_ (.I(\pc[8] ),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6848_ (.A1(_2957_),
    .A2(_2946_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6849_ (.I(_2890_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6850_ (.A1(_2957_),
    .A2(_1722_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6851_ (.A1(_2943_),
    .A2(_2951_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6852_ (.A1(_2931_),
    .A2(_2961_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6853_ (.I(_1671_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6854_ (.A1(_2919_),
    .A2(_2940_),
    .B(_2941_),
    .C(_2961_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6855_ (.A1(_2950_),
    .A2(_1671_),
    .B(_2952_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6856_ (.A1(_0787_),
    .A2(_2963_),
    .B(_2964_),
    .C(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6857_ (.A1(_2921_),
    .A2(_2924_),
    .A3(_2962_),
    .B(_2966_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6858_ (.A1(_2960_),
    .A2(_2967_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6859_ (.A1(net95),
    .A2(_2959_),
    .B1(_2949_),
    .B2(_2968_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6860_ (.A1(_2928_),
    .A2(_2958_),
    .B(_2969_),
    .ZN(\pc_next[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6861_ (.I(_2927_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6862_ (.I(\pc[9] ),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6863_ (.A1(_2971_),
    .A2(\pc[8] ),
    .A3(_2946_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6864_ (.A1(_2957_),
    .A2(_2946_),
    .B(_2971_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6865_ (.A1(_2972_),
    .A2(_2973_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6866_ (.I(_2971_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6867_ (.A1(_2957_),
    .A2(net21),
    .A3(_2939_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6868_ (.A1(_2960_),
    .A2(_2967_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6869_ (.A1(_2976_),
    .A2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6870_ (.A1(_2975_),
    .A2(_1779_),
    .A3(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6871_ (.A1(net96),
    .A2(_2959_),
    .B1(_2949_),
    .B2(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6872_ (.A1(_2970_),
    .A2(_2974_),
    .B(_2980_),
    .ZN(\pc_next[9] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6873_ (.I(\pc[10] ),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6874_ (.A1(_2981_),
    .A2(_2972_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6875_ (.A1(net22),
    .A2(_2939_),
    .B(_2971_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6876_ (.A1(_2975_),
    .A2(_1779_),
    .B(_2976_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6877_ (.A1(_2960_),
    .A2(_2967_),
    .B(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6878_ (.A1(_2983_),
    .A2(_2985_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6879_ (.I(_1822_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6880_ (.A1(_2981_),
    .A2(_2987_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6881_ (.A1(_2986_),
    .A2(_2988_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6882_ (.A1(net66),
    .A2(_2959_),
    .B1(_2949_),
    .B2(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6883_ (.A1(_2970_),
    .A2(_2982_),
    .B(_2990_),
    .ZN(\pc_next[10] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6884_ (.I(_2886_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6885_ (.A1(\pc[11] ),
    .A2(\pc[10] ),
    .A3(_2972_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6886_ (.I(\pc[11] ),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6887_ (.A1(\pc[10] ),
    .A2(_2972_),
    .B(_2993_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6888_ (.A1(_2992_),
    .A2(_2994_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6889_ (.A1(_2993_),
    .A2(net104),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6890_ (.A1(_2981_),
    .A2(_2987_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6891_ (.A1(_2986_),
    .A2(_2988_),
    .B(_2997_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6892_ (.A1(_2996_),
    .A2(_2998_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6893_ (.I(_2890_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6894_ (.A1(net67),
    .A2(_3000_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6895_ (.A1(_2991_),
    .A2(_2995_),
    .B1(_2999_),
    .B2(_2884_),
    .C(_3001_),
    .ZN(\pc_next[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6896_ (.I(\pc[12] ),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6897_ (.I(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6898_ (.A1(_3003_),
    .A2(_2992_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6899_ (.I(_2905_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6900_ (.A1(_0535_),
    .A2(_2167_),
    .B(_2168_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6901_ (.A1(_3002_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6902_ (.A1(_3003_),
    .A2(_1928_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6903_ (.A1(_3007_),
    .A2(_3008_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6904_ (.I(net104),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6905_ (.A1(_2993_),
    .A2(_3010_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6906_ (.A1(_2981_),
    .A2(_2987_),
    .B(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6907_ (.A1(_2993_),
    .A2(_3010_),
    .B(_3012_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6908_ (.I(_2988_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6909_ (.A1(_2983_),
    .A2(_2985_),
    .A3(_3014_),
    .A4(_2996_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6910_ (.A1(_3013_),
    .A2(_3015_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6911_ (.A1(_3009_),
    .A2(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6912_ (.A1(net68),
    .A2(_2959_),
    .B1(_3005_),
    .B2(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6913_ (.A1(_2970_),
    .A2(_3004_),
    .B(_3018_),
    .ZN(\pc_next[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6914_ (.I(\pc[13] ),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6915_ (.A1(_3019_),
    .A2(_3002_),
    .A3(_2992_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6916_ (.A1(_3002_),
    .A2(_2992_),
    .B(_3019_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6917_ (.A1(_3020_),
    .A2(_3021_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6918_ (.I(_2889_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6919_ (.A1(_0519_),
    .A2(_2167_),
    .B(_2168_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6920_ (.A1(_3019_),
    .A2(_3024_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6921_ (.A1(_3009_),
    .A2(_3016_),
    .B(_3007_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6922_ (.A1(_3025_),
    .A2(_3026_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6923_ (.A1(net69),
    .A2(_3023_),
    .B1(_3005_),
    .B2(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6924_ (.A1(_2970_),
    .A2(_3022_),
    .B(_3028_),
    .ZN(\pc_next[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6925_ (.I(\pc[14] ),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6926_ (.I(_3029_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6927_ (.A1(_3030_),
    .A2(_3020_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6928_ (.I(_3019_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6929_ (.A1(_3032_),
    .A2(_1973_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6930_ (.A1(_3032_),
    .A2(_1973_),
    .B(_1928_),
    .C(_3003_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6931_ (.A1(_3007_),
    .A2(_3008_),
    .A3(_3025_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6932_ (.A1(_3013_),
    .A2(_3015_),
    .B(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6933_ (.A1(_0483_),
    .A2(_2167_),
    .B(_2168_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6934_ (.A1(_3029_),
    .A2(_3037_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6935_ (.A1(_3033_),
    .A2(_3034_),
    .A3(_3036_),
    .B(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6936_ (.A1(_3033_),
    .A2(_3038_),
    .A3(_3034_),
    .A4(_3036_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6937_ (.A1(_3039_),
    .A2(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6938_ (.A1(net70),
    .A2(_3000_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6939_ (.A1(_2991_),
    .A2(_3031_),
    .B1(_3041_),
    .B2(_2884_),
    .C(_3042_),
    .ZN(\pc_next[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6940_ (.I(_2927_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6941_ (.I(\pc[15] ),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6942_ (.A1(_3044_),
    .A2(\pc[14] ),
    .A3(_3020_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6943_ (.A1(_3029_),
    .A2(_3020_),
    .B(_3044_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6944_ (.A1(_3045_),
    .A2(_3046_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6945_ (.A1(_3044_),
    .A2(_2069_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6946_ (.A1(_3044_),
    .A2(_2069_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6947_ (.A1(_3048_),
    .A2(_3049_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6948_ (.A1(_3030_),
    .A2(_2027_),
    .B(_3039_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6949_ (.A1(_3050_),
    .A2(_3051_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6950_ (.A1(net71),
    .A2(_3023_),
    .B1(_3005_),
    .B2(_3052_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6951_ (.A1(_3043_),
    .A2(_3047_),
    .B(_3053_),
    .ZN(\pc_next[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6952_ (.I(\pc[16] ),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6953_ (.A1(_3054_),
    .A2(_3045_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6954_ (.A1(_3054_),
    .A2(_2098_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6955_ (.I(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6956_ (.A1(_3029_),
    .A2(_3037_),
    .A3(_3049_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6957_ (.A1(_3038_),
    .A2(_3050_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6958_ (.A1(_3033_),
    .A2(_3034_),
    .A3(_3036_),
    .B(_3059_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6959_ (.A1(_3048_),
    .A2(_3058_),
    .A3(_3060_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6960_ (.A1(_3057_),
    .A2(_3061_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6961_ (.A1(net72),
    .A2(_3023_),
    .B1(_3005_),
    .B2(_3062_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6962_ (.A1(_3043_),
    .A2(_3055_),
    .B(_3063_),
    .ZN(\pc_next[16] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6963_ (.A1(\pc[17] ),
    .A2(\pc[16] ),
    .A3(_3045_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6964_ (.I(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6965_ (.I(\pc[17] ),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6966_ (.A1(_3054_),
    .A2(_3045_),
    .B(_3066_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6967_ (.A1(_3065_),
    .A2(_3067_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6968_ (.I(_2893_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6969_ (.A1(\pc[17] ),
    .A2(_2169_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6970_ (.A1(_3054_),
    .A2(_2098_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6971_ (.A1(_3057_),
    .A2(_3061_),
    .B(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6972_ (.A1(_3070_),
    .A2(_3072_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6973_ (.A1(net73),
    .A2(_3023_),
    .B1(_3069_),
    .B2(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6974_ (.A1(_3043_),
    .A2(_3068_),
    .B(_3074_),
    .ZN(\pc_next[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6975_ (.I(\pc[18] ),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6976_ (.A1(_3075_),
    .A2(_3064_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6977_ (.I(_2889_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6978_ (.A1(_3075_),
    .A2(_2210_),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6979_ (.A1(_3057_),
    .A2(_3070_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6980_ (.I(_2169_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6981_ (.A1(_3066_),
    .A2(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6982_ (.A1(_3071_),
    .A2(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6983_ (.A1(_3066_),
    .A2(_3080_),
    .B(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6984_ (.A1(_3061_),
    .A2(_3079_),
    .B(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6985_ (.A1(_3078_),
    .A2(_3084_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6986_ (.A1(net74),
    .A2(_3077_),
    .B1(_3069_),
    .B2(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6987_ (.A1(_3043_),
    .A2(_3076_),
    .B(_3086_),
    .ZN(\pc_next[18] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6988_ (.I(_2927_),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6989_ (.A1(\pc[19] ),
    .A2(\pc[18] ),
    .A3(_3065_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6990_ (.I(\pc[19] ),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6991_ (.A1(_3075_),
    .A2(_3065_),
    .B(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6992_ (.A1(_3088_),
    .A2(_3090_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6993_ (.A1(\pc[19] ),
    .A2(_2251_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6994_ (.A1(_3075_),
    .A2(_2210_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6995_ (.A1(_3078_),
    .A2(_3084_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6996_ (.A1(_3093_),
    .A2(_3094_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6997_ (.A1(_3092_),
    .A2(_3095_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6998_ (.A1(net75),
    .A2(_3077_),
    .B1(_3069_),
    .B2(_3096_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6999_ (.A1(_3087_),
    .A2(_3091_),
    .B(_3097_),
    .ZN(\pc_next[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7000_ (.I(_2886_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7001_ (.I(\pc[20] ),
    .Z(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7002_ (.A1(_3099_),
    .A2(_3088_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7003_ (.A1(_3099_),
    .A2(_2291_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7004_ (.A1(_3048_),
    .A2(_3058_),
    .A3(_3060_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7005_ (.A1(_3057_),
    .A2(_3070_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7006_ (.A1(_3066_),
    .A2(_3080_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7007_ (.A1(_3071_),
    .A2(_3081_),
    .B(_3104_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7008_ (.A1(_3102_),
    .A2(_3103_),
    .B(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7009_ (.A1(_3078_),
    .A2(_3092_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7010_ (.I(_2251_),
    .Z(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7011_ (.A1(_3089_),
    .A2(_3108_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7012_ (.A1(_3093_),
    .A2(_3109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7013_ (.A1(_3089_),
    .A2(_3108_),
    .B(_3110_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7014_ (.A1(_3106_),
    .A2(_3107_),
    .B(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7015_ (.A1(_3101_),
    .A2(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7016_ (.A1(_3101_),
    .A2(_3112_),
    .B(_3113_),
    .C(_2905_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7017_ (.A1(_2336_),
    .A2(_2880_),
    .B1(_3098_),
    .B2(_3100_),
    .C(_3114_),
    .ZN(\pc_next[20] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7018_ (.A1(\pc[21] ),
    .A2(\pc[20] ),
    .A3(_3088_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7019_ (.I(\pc[21] ),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7020_ (.A1(_3099_),
    .A2(_3088_),
    .B(_3116_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7021_ (.A1(_3115_),
    .A2(_3117_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7022_ (.A1(\pc[21] ),
    .A2(_2339_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7023_ (.A1(_3099_),
    .A2(_2291_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7024_ (.A1(_3120_),
    .A2(_3113_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7025_ (.A1(_3119_),
    .A2(_3121_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7026_ (.A1(net78),
    .A2(_3077_),
    .B1(_3069_),
    .B2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7027_ (.A1(_3087_),
    .A2(_3118_),
    .B(_3123_),
    .ZN(\pc_next[21] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7028_ (.I(\pc[22] ),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7029_ (.A1(_3124_),
    .A2(_3115_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7030_ (.I(_2893_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7031_ (.A1(_3124_),
    .A2(_2379_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7032_ (.A1(_3078_),
    .A2(_3092_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7033_ (.A1(_3089_),
    .A2(_3108_),
    .B1(_3084_),
    .B2(_3128_),
    .C(_3110_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7034_ (.A1(_3101_),
    .A2(_3119_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7035_ (.I(_2339_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7036_ (.A1(_3116_),
    .A2(_3131_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7037_ (.A1(_3120_),
    .A2(_3132_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7038_ (.A1(_3116_),
    .A2(_3131_),
    .B(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7039_ (.A1(_3129_),
    .A2(_3130_),
    .B(_3134_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7040_ (.A1(_3127_),
    .A2(_3135_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7041_ (.A1(net79),
    .A2(_3077_),
    .B1(_3126_),
    .B2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7042_ (.A1(_3087_),
    .A2(_3125_),
    .B(_3137_),
    .ZN(\pc_next[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7043_ (.I(\pc[23] ),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7044_ (.A1(_3124_),
    .A2(_3115_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7045_ (.A1(_3138_),
    .A2(_3139_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7046_ (.A1(_3138_),
    .A2(_2423_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7047_ (.A1(_3138_),
    .A2(_2423_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7048_ (.A1(_3141_),
    .A2(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7049_ (.A1(_3124_),
    .A2(_2379_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7050_ (.A1(_3127_),
    .A2(_3135_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7051_ (.A1(_3144_),
    .A2(_3145_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7052_ (.A1(_3143_),
    .A2(_3146_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7053_ (.A1(_2894_),
    .A2(_3147_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7054_ (.A1(_2458_),
    .A2(_2880_),
    .B1(_2991_),
    .B2(_3140_),
    .C(_3148_),
    .ZN(\pc_next[23] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7055_ (.A1(_3138_),
    .A2(\pc[22] ),
    .A3(_3115_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7056_ (.A1(\pc[24] ),
    .A2(_3149_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7057_ (.I(_2889_),
    .Z(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7058_ (.A1(\pc[24] ),
    .A2(_2460_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _7059_ (.I(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7060_ (.A1(_3127_),
    .A2(_3143_),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7061_ (.A1(_3144_),
    .A2(_3142_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7062_ (.A1(_3135_),
    .A2(_3154_),
    .B(_3155_),
    .C(_3141_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7063_ (.A1(_3153_),
    .A2(_3156_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7064_ (.A1(net81),
    .A2(_3151_),
    .B1(_3126_),
    .B2(_3157_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7065_ (.A1(_3087_),
    .A2(_3150_),
    .B(_3158_),
    .ZN(\pc_next[24] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7066_ (.I(_2886_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7067_ (.I(\pc[25] ),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7068_ (.I(\pc[24] ),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7069_ (.A1(_3161_),
    .A2(_3149_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7070_ (.A1(_3160_),
    .A2(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7071_ (.I(_2511_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7072_ (.A1(_3160_),
    .A2(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7073_ (.A1(\pc[25] ),
    .A2(_3164_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7074_ (.I(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7075_ (.A1(_3165_),
    .A2(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7076_ (.A1(_3101_),
    .A2(_3119_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7077_ (.A1(_3116_),
    .A2(_3131_),
    .B1(_3112_),
    .B2(_3169_),
    .C(_3133_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7078_ (.A1(_3127_),
    .A2(_3143_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7079_ (.A1(_3141_),
    .A2(_3155_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7080_ (.A1(_3170_),
    .A2(_3171_),
    .B(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7081_ (.A1(_3161_),
    .A2(_2586_),
    .A3(_2459_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7082_ (.A1(_3152_),
    .A2(_3173_),
    .B(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7083_ (.A1(_3168_),
    .A2(_3175_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7084_ (.A1(net82),
    .A2(_3151_),
    .B1(_3126_),
    .B2(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7085_ (.A1(_3159_),
    .A2(_3163_),
    .B(_3177_),
    .ZN(\pc_next[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7086_ (.I(_2550_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7087_ (.A1(\pc[26] ),
    .A2(_3178_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7088_ (.I(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7089_ (.A1(_3165_),
    .A2(_3175_),
    .B(_3180_),
    .C(_3166_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7090_ (.A1(_3165_),
    .A2(_3175_),
    .B(_3166_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7091_ (.I(_2893_),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7092_ (.A1(_3179_),
    .A2(_3182_),
    .B(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7093_ (.I(\pc[26] ),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7094_ (.A1(_3160_),
    .A2(_3162_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7095_ (.A1(_3185_),
    .A2(_3186_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7096_ (.A1(net83),
    .A2(_3000_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7097_ (.A1(_3181_),
    .A2(_3184_),
    .B1(_3187_),
    .B2(_3159_),
    .C(_3188_),
    .ZN(\pc_next[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7098_ (.I(\pc[27] ),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7099_ (.I(_3189_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7100_ (.I(_2589_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7101_ (.A1(_3190_),
    .A2(_3191_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7102_ (.A1(_3185_),
    .A2(_3178_),
    .B(_3181_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7103_ (.A1(_3192_),
    .A2(_3193_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7104_ (.A1(_3192_),
    .A2(_3193_),
    .B(_3183_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7105_ (.A1(\pc[25] ),
    .A2(_3185_),
    .A3(_3162_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7106_ (.A1(_3189_),
    .A2(_3196_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7107_ (.A1(net84),
    .A2(_2891_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7108_ (.A1(_3194_),
    .A2(_3195_),
    .B1(_3197_),
    .B2(_3159_),
    .C(_3198_),
    .ZN(\pc_next[27] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7109_ (.I(\pc[28] ),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7110_ (.A1(_3190_),
    .A2(_3196_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7111_ (.A1(_3199_),
    .A2(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7112_ (.A1(_3180_),
    .A2(_3192_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7113_ (.A1(_3168_),
    .A2(_3202_),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7114_ (.A1(_3160_),
    .A2(_3164_),
    .B(_3174_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7115_ (.A1(_3185_),
    .A2(_3178_),
    .B1(_3191_),
    .B2(_3189_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7116_ (.A1(_3189_),
    .A2(_3191_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7117_ (.A1(_3166_),
    .A2(_3202_),
    .A3(_3204_),
    .B1(_3205_),
    .B2(_3206_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7118_ (.I(_3207_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _7119_ (.A1(_3153_),
    .A2(_3156_),
    .A3(_3203_),
    .B(_3208_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7120_ (.A1(\pc[28] ),
    .A2(_2637_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7121_ (.A1(_3209_),
    .A2(_3210_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7122_ (.A1(net85),
    .A2(_3151_),
    .B1(_3126_),
    .B2(_3211_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7123_ (.A1(_3159_),
    .A2(_3201_),
    .B(_3212_),
    .ZN(\pc_next[28] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7124_ (.I(\pc[29] ),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7125_ (.A1(_3199_),
    .A2(_3200_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7126_ (.A1(_3213_),
    .A2(_3214_),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7127_ (.I(_2683_),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7128_ (.A1(\pc[29] ),
    .A2(_3216_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7129_ (.A1(_3199_),
    .A2(_2637_),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7130_ (.A1(_3209_),
    .A2(_3210_),
    .B(_3218_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7131_ (.A1(_3217_),
    .A2(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7132_ (.A1(_2894_),
    .A2(_3220_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7133_ (.A1(_2710_),
    .A2(_2880_),
    .B1(_2991_),
    .B2(_3215_),
    .C(_3221_),
    .ZN(\pc_next[29] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7134_ (.I(\pc[30] ),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7135_ (.A1(_3213_),
    .A2(_3199_),
    .A3(_3200_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7136_ (.A1(_3222_),
    .A2(_3223_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7137_ (.A1(net88),
    .A2(_3000_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7138_ (.A1(_3210_),
    .A2(_3217_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7139_ (.A1(_3213_),
    .A2(_3216_),
    .B(_3218_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7140_ (.I(_3227_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7141_ (.A1(_3213_),
    .A2(_3216_),
    .B1(_3209_),
    .B2(_3226_),
    .C(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7142_ (.A1(_3222_),
    .A2(_2716_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7143_ (.A1(_3229_),
    .A2(_3230_),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7144_ (.A1(_2894_),
    .A2(_3231_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7145_ (.A1(_3098_),
    .A2(_3224_),
    .B(_3225_),
    .C(_3232_),
    .ZN(\pc_next[30] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7146_ (.A1(_2586_),
    .A2(_2715_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7147_ (.A1(_3222_),
    .A2(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7148_ (.A1(_3229_),
    .A2(_3230_),
    .B(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7149_ (.A1(_1874_),
    .A2(\pc[31] ),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7150_ (.A1(_3235_),
    .A2(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7151_ (.A1(_3235_),
    .A2(_3236_),
    .B(_3183_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7152_ (.A1(\pc[29] ),
    .A2(\pc[28] ),
    .A3(_3222_),
    .A4(_3200_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7153_ (.A1(\pc[31] ),
    .A2(_3239_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7154_ (.A1(net89),
    .A2(_2891_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7155_ (.A1(_3237_),
    .A2(_3238_),
    .B1(_3240_),
    .B2(_3098_),
    .C(_3241_),
    .ZN(\pc_next[31] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7156_ (.A1(_0497_),
    .A2(_0516_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7157_ (.I(_3242_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7158_ (.A1(_0496_),
    .A2(_0582_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7159_ (.A1(_3243_),
    .A2(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7160_ (.I(_3242_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7161_ (.A1(net33),
    .A2(_3246_),
    .B1(_3244_),
    .B2(\pc[0] ),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7162_ (.A1(_0554_),
    .A2(_3245_),
    .B(_3247_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7163_ (.A1(_0494_),
    .A2(_0484_),
    .A3(_0583_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7164_ (.A1(net106),
    .A2(_3249_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7165_ (.I(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7166_ (.I0(net65),
    .I1(_3248_),
    .S(_3251_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7167_ (.I(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7168_ (.I(_3253_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7169_ (.I(net31),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7170_ (.I(net30),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7171_ (.A1(_3255_),
    .A2(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7172_ (.I(net2),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7173_ (.I(net32),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7174_ (.A1(_3242_),
    .A2(_3244_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7175_ (.A1(_0489_),
    .A2(_0502_),
    .A3(_0501_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7176_ (.A1(_3260_),
    .A2(_3261_),
    .B(net3),
    .C(_2888_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7177_ (.I(_3262_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7178_ (.A1(_3258_),
    .A2(_3259_),
    .A3(_3263_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7179_ (.A1(_3257_),
    .A2(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7180_ (.I(_3265_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7181_ (.I(_3266_),
    .Z(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7182_ (.I0(\reg_file.reg_storage[11][0] ),
    .I1(_3254_),
    .S(_3267_),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7183_ (.I(_3268_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7184_ (.I(_3250_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7185_ (.A1(net44),
    .A2(_3246_),
    .B1(_3244_),
    .B2(\pc[1] ),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7186_ (.A1(_0642_),
    .A2(_3245_),
    .B(_3270_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_3251_),
    .A2(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7188_ (.A1(_2878_),
    .A2(_3269_),
    .B(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7189_ (.I(_3273_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7190_ (.I(_3274_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7191_ (.I0(\reg_file.reg_storage[11][1] ),
    .I1(_3275_),
    .S(_3267_),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7192_ (.I(_3276_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7193_ (.A1(net107),
    .A2(_3249_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7194_ (.I(_3277_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7195_ (.I(_3260_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7196_ (.I(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7197_ (.I(_2881_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7198_ (.A1(_2879_),
    .A2(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7199_ (.A1(net55),
    .A2(_3246_),
    .B1(_2895_),
    .B2(_3280_),
    .C(_3282_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7200_ (.A1(net87),
    .A2(_3278_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7201_ (.A1(_3278_),
    .A2(_3283_),
    .B(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7202_ (.I(_3285_),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7203_ (.I(_3286_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7204_ (.I0(\reg_file.reg_storage[11][2] ),
    .I1(_3287_),
    .S(_3267_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7205_ (.I(_3288_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7206_ (.I(_3280_),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7207_ (.A1(_2907_),
    .A2(_3289_),
    .A3(_3251_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7208_ (.I(_3277_),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7209_ (.A1(_3281_),
    .A2(_2904_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7210_ (.A1(net58),
    .A2(_3246_),
    .B(_3291_),
    .C(_3292_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7211_ (.A1(_1474_),
    .A2(_3278_),
    .B1(_3290_),
    .B2(_3293_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7212_ (.I(_3294_),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7213_ (.I(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7214_ (.I0(\reg_file.reg_storage[11][3] ),
    .I1(_3296_),
    .S(_3267_),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7215_ (.I(_3297_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7216_ (.I(_3265_),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7217_ (.I(_3298_),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7218_ (.I(_3299_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7219_ (.I(_3250_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7220_ (.I(_3301_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7221_ (.I(_3245_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7222_ (.I(_3242_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7223_ (.I(_3304_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7224_ (.A1(_3281_),
    .A2(_2917_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7225_ (.A1(net59),
    .A2(_3305_),
    .B(_3306_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7226_ (.A1(_1089_),
    .A2(_3303_),
    .B(_3269_),
    .C(_3307_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7227_ (.A1(net91),
    .A2(_3302_),
    .B(_3308_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7228_ (.I(_3309_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7229_ (.I(_3265_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7230_ (.I(_3311_),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7231_ (.A1(\reg_file.reg_storage[11][4] ),
    .A2(_3312_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7232_ (.A1(_3300_),
    .A2(_3310_),
    .B(_3313_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7233_ (.I(_3243_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7234_ (.A1(_3281_),
    .A2(_2930_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7235_ (.A1(net60),
    .A2(_3314_),
    .B(_3315_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7236_ (.A1(_1539_),
    .A2(_3303_),
    .B(_3269_),
    .C(_3316_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7237_ (.A1(net92),
    .A2(_3302_),
    .B(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7238_ (.I(_3318_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7239_ (.A1(\reg_file.reg_storage[11][5] ),
    .A2(_3312_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7240_ (.A1(_3300_),
    .A2(_3319_),
    .B(_3320_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _7241_ (.I(_3251_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7242_ (.I(_2881_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7243_ (.I(_3322_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7244_ (.A1(_3323_),
    .A2(_2938_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7245_ (.A1(net61),
    .A2(_3305_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7246_ (.A1(_1627_),
    .A2(_3303_),
    .B(_3269_),
    .C(_3325_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7247_ (.A1(net93),
    .A2(_3321_),
    .B1(_3324_),
    .B2(_3326_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7248_ (.I(_3327_),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7249_ (.A1(\reg_file.reg_storage[11][6] ),
    .A2(_3312_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7250_ (.A1(_3300_),
    .A2(_3328_),
    .B(_3329_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7251_ (.I(_2881_),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7252_ (.I(_3330_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7253_ (.A1(net62),
    .A2(_3314_),
    .B1(_2963_),
    .B2(_3289_),
    .C(_3278_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7254_ (.A1(_3331_),
    .A2(_2948_),
    .B(_3332_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7255_ (.A1(net94),
    .A2(_3302_),
    .B(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7256_ (.I(_3334_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7257_ (.A1(\reg_file.reg_storage[11][7] ),
    .A2(_3312_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7258_ (.A1(_3300_),
    .A2(_3335_),
    .B(_3336_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7259_ (.I(_3299_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7260_ (.A1(_3330_),
    .A2(_2958_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7261_ (.A1(net63),
    .A2(_3305_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7262_ (.A1(_1722_),
    .A2(_3303_),
    .B(_3301_),
    .C(_3339_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7263_ (.A1(net95),
    .A2(_3321_),
    .B1(_3338_),
    .B2(_3340_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7264_ (.I(_3341_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7265_ (.I(_3311_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7266_ (.A1(\reg_file.reg_storage[11][8] ),
    .A2(_3343_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7267_ (.A1(_3337_),
    .A2(_3342_),
    .B(_3344_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7268_ (.A1(_3330_),
    .A2(_2974_),
    .ZN(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7269_ (.A1(net64),
    .A2(_3305_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7270_ (.A1(_1779_),
    .A2(_3245_),
    .B(_3301_),
    .C(_3346_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7271_ (.A1(net96),
    .A2(_3321_),
    .B1(_3345_),
    .B2(_3347_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7272_ (.I(_3348_),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7273_ (.A1(\reg_file.reg_storage[11][9] ),
    .A2(_3343_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7274_ (.A1(_3337_),
    .A2(_3349_),
    .B(_3350_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7275_ (.I(_2987_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7276_ (.I(_3291_),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7277_ (.A1(net34),
    .A2(_3314_),
    .B1(_3351_),
    .B2(_3289_),
    .C(_3352_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7278_ (.A1(_3331_),
    .A2(_2982_),
    .B(_3353_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7279_ (.A1(net66),
    .A2(_3302_),
    .B(_3354_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7280_ (.I(_3355_),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7281_ (.A1(\reg_file.reg_storage[11][10] ),
    .A2(_3343_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7282_ (.A1(_3337_),
    .A2(_3356_),
    .B(_3357_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7283_ (.I(_3301_),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7284_ (.A1(net35),
    .A2(_3314_),
    .B1(_3010_),
    .B2(_3289_),
    .C(_3352_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7285_ (.A1(_3331_),
    .A2(_2995_),
    .B(_3359_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7286_ (.A1(net67),
    .A2(_3358_),
    .B(_3360_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7287_ (.I(_3361_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7288_ (.A1(\reg_file.reg_storage[11][11] ),
    .A2(_3343_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7289_ (.A1(_3337_),
    .A2(_3362_),
    .B(_3363_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7290_ (.I(_3299_),
    .Z(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7291_ (.I(_3304_),
    .Z(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7292_ (.I(_3280_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7293_ (.A1(net36),
    .A2(_3365_),
    .B1(_3006_),
    .B2(_3366_),
    .C(_3352_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7294_ (.A1(_3331_),
    .A2(_3004_),
    .B(_3367_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7295_ (.A1(net68),
    .A2(_3358_),
    .B(_3368_),
    .ZN(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7296_ (.I(_3369_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7297_ (.I(_3311_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7298_ (.A1(\reg_file.reg_storage[11][12] ),
    .A2(_3371_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7299_ (.A1(_3364_),
    .A2(_3370_),
    .B(_3372_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7300_ (.I(_3330_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7301_ (.A1(net37),
    .A2(_3365_),
    .B1(_3024_),
    .B2(_3366_),
    .C(_3352_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7302_ (.A1(_3373_),
    .A2(_3022_),
    .B(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7303_ (.A1(net69),
    .A2(_3358_),
    .B(_3375_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7304_ (.I(_3376_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7305_ (.A1(\reg_file.reg_storage[11][13] ),
    .A2(_3371_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7306_ (.A1(_3364_),
    .A2(_3377_),
    .B(_3378_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7307_ (.I(_3277_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7308_ (.I(_3379_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7309_ (.A1(net38),
    .A2(_3365_),
    .B1(_3037_),
    .B2(_3366_),
    .C(_3380_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7310_ (.A1(_3373_),
    .A2(_3031_),
    .B(_3381_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7311_ (.A1(net70),
    .A2(_3358_),
    .B(_3382_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7312_ (.I(_3383_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7313_ (.A1(\reg_file.reg_storage[11][14] ),
    .A2(_3371_),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7314_ (.A1(_3364_),
    .A2(_3384_),
    .B(_3385_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7315_ (.I(_3250_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7316_ (.I(_3386_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7317_ (.A1(net39),
    .A2(_3365_),
    .B1(_2069_),
    .B2(_3366_),
    .C(_3380_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7318_ (.A1(_3373_),
    .A2(_3047_),
    .B(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7319_ (.A1(net71),
    .A2(_3387_),
    .B(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7320_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7321_ (.A1(\reg_file.reg_storage[11][15] ),
    .A2(_3371_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7322_ (.A1(_3364_),
    .A2(_3391_),
    .B(_3392_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7323_ (.I(_3299_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7324_ (.I(_3304_),
    .Z(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7325_ (.I(_3280_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7326_ (.A1(net40),
    .A2(_3394_),
    .B1(_2098_),
    .B2(_3395_),
    .C(_3380_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7327_ (.A1(_3373_),
    .A2(_3055_),
    .B(_3396_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7328_ (.A1(net72),
    .A2(_3387_),
    .B(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7329_ (.I(_3398_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7330_ (.I(_3311_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7331_ (.A1(\reg_file.reg_storage[11][16] ),
    .A2(_3400_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7332_ (.A1(_3393_),
    .A2(_3399_),
    .B(_3401_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7333_ (.I(_3322_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7334_ (.A1(net41),
    .A2(_3394_),
    .B1(_3080_),
    .B2(_3395_),
    .C(_3380_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7335_ (.A1(_3402_),
    .A2(_3068_),
    .B(_3403_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7336_ (.A1(net73),
    .A2(_3387_),
    .B(_3404_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7337_ (.I(_3405_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7338_ (.A1(\reg_file.reg_storage[11][17] ),
    .A2(_3400_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7339_ (.A1(_3393_),
    .A2(_3406_),
    .B(_3407_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7340_ (.I(_3379_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7341_ (.A1(net42),
    .A2(_3394_),
    .B1(_2210_),
    .B2(_3395_),
    .C(_3408_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7342_ (.A1(_3402_),
    .A2(_3076_),
    .B(_3409_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7343_ (.A1(net74),
    .A2(_3387_),
    .B(_3410_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7344_ (.I(_3411_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7345_ (.A1(\reg_file.reg_storage[11][18] ),
    .A2(_3400_),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7346_ (.A1(_3393_),
    .A2(_3412_),
    .B(_3413_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7347_ (.I(_3386_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7348_ (.A1(net43),
    .A2(_3394_),
    .B1(_3108_),
    .B2(_3395_),
    .C(_3408_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7349_ (.A1(_3402_),
    .A2(_3091_),
    .B(_3415_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7350_ (.A1(net75),
    .A2(_3414_),
    .B(_3416_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7351_ (.I(_3417_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7352_ (.A1(\reg_file.reg_storage[11][19] ),
    .A2(_3400_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7353_ (.A1(_3393_),
    .A2(_3418_),
    .B(_3419_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7354_ (.I(_3266_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7355_ (.I(_3304_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7356_ (.I(_3279_),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7357_ (.A1(net45),
    .A2(_3421_),
    .B1(_2291_),
    .B2(_3422_),
    .C(_3408_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7358_ (.A1(_3402_),
    .A2(_3100_),
    .B(_3423_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7359_ (.A1(net77),
    .A2(_3414_),
    .B(_3424_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7360_ (.I(_3425_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7361_ (.I(_3298_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7362_ (.A1(\reg_file.reg_storage[11][20] ),
    .A2(_3427_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7363_ (.A1(_3420_),
    .A2(_3426_),
    .B(_3428_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7364_ (.I(_3322_),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7365_ (.A1(net46),
    .A2(_3421_),
    .B1(_3131_),
    .B2(_3422_),
    .C(_3408_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7366_ (.A1(_3429_),
    .A2(_3118_),
    .B(_3430_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7367_ (.A1(net78),
    .A2(_3414_),
    .B(_3431_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7368_ (.I(_3432_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7369_ (.A1(\reg_file.reg_storage[11][21] ),
    .A2(_3427_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7370_ (.A1(_3420_),
    .A2(_3433_),
    .B(_3434_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7371_ (.I(_3379_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7372_ (.A1(net47),
    .A2(_3421_),
    .B1(_2379_),
    .B2(_3422_),
    .C(_3435_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7373_ (.A1(_3429_),
    .A2(_3125_),
    .B(_3436_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7374_ (.A1(net79),
    .A2(_3414_),
    .B(_3437_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7375_ (.I(_3438_),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7376_ (.A1(\reg_file.reg_storage[11][22] ),
    .A2(_3427_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7377_ (.A1(_3420_),
    .A2(_3439_),
    .B(_3440_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7378_ (.I(_3386_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7379_ (.A1(net48),
    .A2(_3421_),
    .B1(_2423_),
    .B2(_3422_),
    .C(_3435_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7380_ (.A1(_3429_),
    .A2(_3140_),
    .B(_3442_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7381_ (.A1(net80),
    .A2(_3441_),
    .B(_3443_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7382_ (.I(_3444_),
    .Z(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7383_ (.A1(\reg_file.reg_storage[11][23] ),
    .A2(_3427_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7384_ (.A1(_3420_),
    .A2(_3445_),
    .B(_3446_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7385_ (.I(_3266_),
    .Z(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7386_ (.I(_3243_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7387_ (.I(_3279_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7388_ (.A1(net49),
    .A2(_3448_),
    .B1(_2460_),
    .B2(_3449_),
    .C(_3435_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7389_ (.A1(_3429_),
    .A2(_3150_),
    .B(_3450_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7390_ (.A1(net81),
    .A2(_3441_),
    .B(_3451_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7391_ (.I(_3452_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7392_ (.I(_3298_),
    .Z(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7393_ (.A1(\reg_file.reg_storage[11][24] ),
    .A2(_3454_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7394_ (.A1(_3447_),
    .A2(_3453_),
    .B(_3455_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7395_ (.I(_3322_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7396_ (.A1(net50),
    .A2(_3448_),
    .B1(_3164_),
    .B2(_3449_),
    .C(_3435_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7397_ (.A1(_3456_),
    .A2(_3163_),
    .B(_3457_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7398_ (.A1(net82),
    .A2(_3441_),
    .B(_3458_),
    .ZN(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7399_ (.I(_3459_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7400_ (.A1(\reg_file.reg_storage[11][25] ),
    .A2(_3454_),
    .ZN(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7401_ (.A1(_3447_),
    .A2(_3460_),
    .B(_3461_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7402_ (.I(_3379_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7403_ (.A1(net51),
    .A2(_3448_),
    .B1(_3178_),
    .B2(_3449_),
    .C(_3462_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7404_ (.A1(_3456_),
    .A2(_3187_),
    .B(_3463_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7405_ (.A1(net83),
    .A2(_3441_),
    .B(_3464_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7406_ (.I(_3465_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7407_ (.A1(\reg_file.reg_storage[11][26] ),
    .A2(_3454_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7408_ (.A1(_3447_),
    .A2(_3466_),
    .B(_3467_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7409_ (.I(_3386_),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7410_ (.A1(net52),
    .A2(_3448_),
    .B1(_3191_),
    .B2(_3449_),
    .C(_3462_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7411_ (.A1(_3456_),
    .A2(_3197_),
    .B(_3469_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7412_ (.A1(net84),
    .A2(_3468_),
    .B(_3470_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7413_ (.I(_3471_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7414_ (.A1(\reg_file.reg_storage[11][27] ),
    .A2(_3454_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7415_ (.A1(_3447_),
    .A2(_3472_),
    .B(_3473_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7416_ (.I(_3266_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7417_ (.I(_3243_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7418_ (.I(_3279_),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7419_ (.A1(net53),
    .A2(_3475_),
    .B1(_2637_),
    .B2(_3476_),
    .C(_3462_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7420_ (.A1(_3456_),
    .A2(_3201_),
    .B(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7421_ (.A1(net85),
    .A2(_3468_),
    .B(_3478_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7422_ (.I(_3479_),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7423_ (.I(_3298_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7424_ (.A1(\reg_file.reg_storage[11][28] ),
    .A2(_3481_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7425_ (.A1(_3474_),
    .A2(_3480_),
    .B(_3482_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7426_ (.A1(net54),
    .A2(_3475_),
    .B1(_3216_),
    .B2(_3476_),
    .C(_3462_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7427_ (.A1(_3323_),
    .A2(_3215_),
    .B(_3483_),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7428_ (.A1(net86),
    .A2(_3468_),
    .B(_3484_),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7429_ (.I(_3485_),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7430_ (.A1(\reg_file.reg_storage[11][29] ),
    .A2(_3481_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7431_ (.A1(_3474_),
    .A2(_3486_),
    .B(_3487_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7432_ (.A1(net56),
    .A2(_3475_),
    .B1(_3233_),
    .B2(_3476_),
    .C(_3291_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7433_ (.A1(_3323_),
    .A2(_3224_),
    .B(_3488_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7434_ (.A1(net88),
    .A2(_3468_),
    .B(_3489_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7435_ (.I(_3490_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7436_ (.A1(\reg_file.reg_storage[11][30] ),
    .A2(_3481_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7437_ (.A1(_3474_),
    .A2(_3491_),
    .B(_3492_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7438_ (.A1(net57),
    .A2(_3475_),
    .B1(_3476_),
    .B2(_1874_),
    .C(_3291_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7439_ (.A1(_3323_),
    .A2(_3240_),
    .B(_3493_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7440_ (.A1(net89),
    .A2(_3321_),
    .B(_3494_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7441_ (.I(_3495_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7442_ (.A1(\reg_file.reg_storage[11][31] ),
    .A2(_3481_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7443_ (.A1(_3474_),
    .A2(_3496_),
    .B(_3497_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7444_ (.I(_3262_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7445_ (.A1(net2),
    .A2(_3259_),
    .A3(_3498_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7446_ (.A1(_3257_),
    .A2(_3499_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7447_ (.I(_3500_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7448_ (.I(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7449_ (.I0(\reg_file.reg_storage[7][0] ),
    .I1(_3254_),
    .S(_3502_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7450_ (.I(_3503_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7451_ (.I(_3500_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7452_ (.I0(\reg_file.reg_storage[7][1] ),
    .I1(_3275_),
    .S(_3504_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7453_ (.I(_3505_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7454_ (.I0(\reg_file.reg_storage[7][2] ),
    .I1(_3287_),
    .S(_3504_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7455_ (.I(_3506_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7456_ (.I0(\reg_file.reg_storage[7][3] ),
    .I1(_3296_),
    .S(_3504_),
    .Z(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7457_ (.I(_3507_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7458_ (.I(_3501_),
    .Z(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7459_ (.I(_3508_),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7460_ (.I(_3504_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7461_ (.A1(\reg_file.reg_storage[7][4] ),
    .A2(_3510_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7462_ (.A1(_3310_),
    .A2(_3509_),
    .B(_3511_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7463_ (.A1(\reg_file.reg_storage[7][5] ),
    .A2(_3510_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7464_ (.A1(_3319_),
    .A2(_3509_),
    .B(_3512_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7465_ (.A1(\reg_file.reg_storage[7][6] ),
    .A2(_3510_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7466_ (.A1(_3328_),
    .A2(_3509_),
    .B(_3513_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7467_ (.A1(\reg_file.reg_storage[7][7] ),
    .A2(_3510_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7468_ (.A1(_3335_),
    .A2(_3509_),
    .B(_3514_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7469_ (.I(_3508_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7470_ (.I(_3500_),
    .Z(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7471_ (.I(_3516_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7472_ (.A1(\reg_file.reg_storage[7][8] ),
    .A2(_3517_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7473_ (.A1(_3342_),
    .A2(_3515_),
    .B(_3518_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7474_ (.A1(\reg_file.reg_storage[7][9] ),
    .A2(_3517_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7475_ (.A1(_3349_),
    .A2(_3515_),
    .B(_3519_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7476_ (.A1(\reg_file.reg_storage[7][10] ),
    .A2(_3517_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7477_ (.A1(_3356_),
    .A2(_3515_),
    .B(_3520_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7478_ (.A1(\reg_file.reg_storage[7][11] ),
    .A2(_3517_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7479_ (.A1(_3362_),
    .A2(_3515_),
    .B(_3521_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7480_ (.I(_3508_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7481_ (.I(_3516_),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7482_ (.A1(\reg_file.reg_storage[7][12] ),
    .A2(_3523_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7483_ (.A1(_3370_),
    .A2(_3522_),
    .B(_3524_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7484_ (.A1(\reg_file.reg_storage[7][13] ),
    .A2(_3523_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7485_ (.A1(_3377_),
    .A2(_3522_),
    .B(_3525_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7486_ (.A1(\reg_file.reg_storage[7][14] ),
    .A2(_3523_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7487_ (.A1(_3384_),
    .A2(_3522_),
    .B(_3526_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7488_ (.A1(\reg_file.reg_storage[7][15] ),
    .A2(_3523_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7489_ (.A1(_3391_),
    .A2(_3522_),
    .B(_3527_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7490_ (.I(_3508_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7491_ (.I(_3516_),
    .Z(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7492_ (.A1(\reg_file.reg_storage[7][16] ),
    .A2(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7493_ (.A1(_3399_),
    .A2(_3528_),
    .B(_3530_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7494_ (.A1(\reg_file.reg_storage[7][17] ),
    .A2(_3529_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7495_ (.A1(_3406_),
    .A2(_3528_),
    .B(_3531_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7496_ (.A1(\reg_file.reg_storage[7][18] ),
    .A2(_3529_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7497_ (.A1(_3412_),
    .A2(_3528_),
    .B(_3532_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7498_ (.A1(\reg_file.reg_storage[7][19] ),
    .A2(_3529_),
    .ZN(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7499_ (.A1(_3418_),
    .A2(_3528_),
    .B(_3533_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7500_ (.I(_3502_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7501_ (.I(_3516_),
    .Z(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7502_ (.A1(\reg_file.reg_storage[7][20] ),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7503_ (.A1(_3426_),
    .A2(_3534_),
    .B(_3536_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7504_ (.A1(\reg_file.reg_storage[7][21] ),
    .A2(_3535_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7505_ (.A1(_3433_),
    .A2(_3534_),
    .B(_3537_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7506_ (.A1(\reg_file.reg_storage[7][22] ),
    .A2(_3535_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7507_ (.A1(_3439_),
    .A2(_3534_),
    .B(_3538_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7508_ (.A1(\reg_file.reg_storage[7][23] ),
    .A2(_3535_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7509_ (.A1(_3445_),
    .A2(_3534_),
    .B(_3539_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7510_ (.I(_3502_),
    .Z(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7511_ (.I(_3501_),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7512_ (.A1(\reg_file.reg_storage[7][24] ),
    .A2(_3541_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7513_ (.A1(_3453_),
    .A2(_3540_),
    .B(_3542_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7514_ (.A1(\reg_file.reg_storage[7][25] ),
    .A2(_3541_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7515_ (.A1(_3460_),
    .A2(_3540_),
    .B(_3543_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7516_ (.A1(\reg_file.reg_storage[7][26] ),
    .A2(_3541_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7517_ (.A1(_3466_),
    .A2(_3540_),
    .B(_3544_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7518_ (.A1(\reg_file.reg_storage[7][27] ),
    .A2(_3541_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7519_ (.A1(_3472_),
    .A2(_3540_),
    .B(_3545_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7520_ (.I(_3502_),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7521_ (.I(_3501_),
    .Z(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7522_ (.A1(\reg_file.reg_storage[7][28] ),
    .A2(_3547_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7523_ (.A1(_3480_),
    .A2(_3546_),
    .B(_3548_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7524_ (.A1(\reg_file.reg_storage[7][29] ),
    .A2(_3547_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7525_ (.A1(_3486_),
    .A2(_3546_),
    .B(_3549_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7526_ (.A1(\reg_file.reg_storage[7][30] ),
    .A2(_3547_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7527_ (.A1(_3491_),
    .A2(_3546_),
    .B(_3550_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7528_ (.A1(\reg_file.reg_storage[7][31] ),
    .A2(_3547_),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7529_ (.A1(_3496_),
    .A2(_3546_),
    .B(_3551_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7530_ (.I(_3255_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7531_ (.I(net30),
    .Z(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7532_ (.A1(_3552_),
    .A2(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7533_ (.A1(_3264_),
    .A2(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7534_ (.I(_3555_),
    .Z(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7535_ (.I(_3556_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7536_ (.I0(\reg_file.reg_storage[9][0] ),
    .I1(_3254_),
    .S(_3557_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7537_ (.I(_3558_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7538_ (.I(_3555_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7539_ (.I0(\reg_file.reg_storage[9][1] ),
    .I1(_3275_),
    .S(_3559_),
    .Z(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7540_ (.I(_3560_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7541_ (.I0(\reg_file.reg_storage[9][2] ),
    .I1(_3287_),
    .S(_3559_),
    .Z(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7542_ (.I(_3561_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7543_ (.I0(\reg_file.reg_storage[9][3] ),
    .I1(_3296_),
    .S(_3559_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7544_ (.I(_3562_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7545_ (.I(_3556_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7546_ (.I(_3563_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7547_ (.I(_3559_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7548_ (.A1(\reg_file.reg_storage[9][4] ),
    .A2(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7549_ (.A1(_3310_),
    .A2(_3564_),
    .B(_3566_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7550_ (.A1(\reg_file.reg_storage[9][5] ),
    .A2(_3565_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7551_ (.A1(_3319_),
    .A2(_3564_),
    .B(_3567_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7552_ (.A1(\reg_file.reg_storage[9][6] ),
    .A2(_3565_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7553_ (.A1(_3328_),
    .A2(_3564_),
    .B(_3568_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7554_ (.A1(\reg_file.reg_storage[9][7] ),
    .A2(_3565_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7555_ (.A1(_3335_),
    .A2(_3564_),
    .B(_3569_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7556_ (.I(_3563_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7557_ (.I(_3555_),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7558_ (.I(_3571_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7559_ (.A1(\reg_file.reg_storage[9][8] ),
    .A2(_3572_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7560_ (.A1(_3342_),
    .A2(_3570_),
    .B(_3573_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7561_ (.A1(\reg_file.reg_storage[9][9] ),
    .A2(_3572_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7562_ (.A1(_3349_),
    .A2(_3570_),
    .B(_3574_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7563_ (.A1(\reg_file.reg_storage[9][10] ),
    .A2(_3572_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7564_ (.A1(_3356_),
    .A2(_3570_),
    .B(_3575_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7565_ (.A1(\reg_file.reg_storage[9][11] ),
    .A2(_3572_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7566_ (.A1(_3362_),
    .A2(_3570_),
    .B(_3576_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7567_ (.I(_3563_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7568_ (.I(_3571_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7569_ (.A1(\reg_file.reg_storage[9][12] ),
    .A2(_3578_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7570_ (.A1(_3370_),
    .A2(_3577_),
    .B(_3579_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7571_ (.A1(\reg_file.reg_storage[9][13] ),
    .A2(_3578_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7572_ (.A1(_3377_),
    .A2(_3577_),
    .B(_3580_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7573_ (.A1(\reg_file.reg_storage[9][14] ),
    .A2(_3578_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7574_ (.A1(_3384_),
    .A2(_3577_),
    .B(_3581_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7575_ (.A1(\reg_file.reg_storage[9][15] ),
    .A2(_3578_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7576_ (.A1(_3391_),
    .A2(_3577_),
    .B(_3582_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7577_ (.I(_3563_),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7578_ (.I(_3571_),
    .Z(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7579_ (.A1(\reg_file.reg_storage[9][16] ),
    .A2(_3584_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7580_ (.A1(_3399_),
    .A2(_3583_),
    .B(_3585_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7581_ (.A1(\reg_file.reg_storage[9][17] ),
    .A2(_3584_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7582_ (.A1(_3406_),
    .A2(_3583_),
    .B(_3586_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7583_ (.A1(\reg_file.reg_storage[9][18] ),
    .A2(_3584_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7584_ (.A1(_3412_),
    .A2(_3583_),
    .B(_3587_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7585_ (.A1(\reg_file.reg_storage[9][19] ),
    .A2(_3584_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7586_ (.A1(_3418_),
    .A2(_3583_),
    .B(_3588_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7587_ (.I(_3557_),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7588_ (.I(_3571_),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7589_ (.A1(\reg_file.reg_storage[9][20] ),
    .A2(_3590_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7590_ (.A1(_3426_),
    .A2(_3589_),
    .B(_3591_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7591_ (.A1(\reg_file.reg_storage[9][21] ),
    .A2(_3590_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7592_ (.A1(_3433_),
    .A2(_3589_),
    .B(_3592_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7593_ (.A1(\reg_file.reg_storage[9][22] ),
    .A2(_3590_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7594_ (.A1(_3439_),
    .A2(_3589_),
    .B(_3593_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7595_ (.A1(\reg_file.reg_storage[9][23] ),
    .A2(_3590_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7596_ (.A1(_3445_),
    .A2(_3589_),
    .B(_3594_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7597_ (.I(_3557_),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7598_ (.I(_3556_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7599_ (.A1(\reg_file.reg_storage[9][24] ),
    .A2(_3596_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7600_ (.A1(_3453_),
    .A2(_3595_),
    .B(_3597_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7601_ (.A1(\reg_file.reg_storage[9][25] ),
    .A2(_3596_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7602_ (.A1(_3460_),
    .A2(_3595_),
    .B(_3598_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7603_ (.A1(\reg_file.reg_storage[9][26] ),
    .A2(_3596_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7604_ (.A1(_3466_),
    .A2(_3595_),
    .B(_3599_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7605_ (.A1(\reg_file.reg_storage[9][27] ),
    .A2(_3596_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7606_ (.A1(_3472_),
    .A2(_3595_),
    .B(_3600_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7607_ (.I(_3557_),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7608_ (.I(_3556_),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7609_ (.A1(\reg_file.reg_storage[9][28] ),
    .A2(_3602_),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7610_ (.A1(_3480_),
    .A2(_3601_),
    .B(_3603_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7611_ (.A1(\reg_file.reg_storage[9][29] ),
    .A2(_3602_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7612_ (.A1(_3486_),
    .A2(_3601_),
    .B(_3604_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7613_ (.A1(\reg_file.reg_storage[9][30] ),
    .A2(_3602_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7614_ (.A1(_3491_),
    .A2(_3601_),
    .B(_3605_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7615_ (.A1(\reg_file.reg_storage[9][31] ),
    .A2(_3602_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7616_ (.A1(_3496_),
    .A2(_3601_),
    .B(_3606_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7617_ (.I(net31),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7618_ (.I(_3256_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7619_ (.A1(_3607_),
    .A2(_3608_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7620_ (.A1(_3264_),
    .A2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7621_ (.I(_3610_),
    .Z(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7622_ (.I(_3611_),
    .Z(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7623_ (.I0(\reg_file.reg_storage[10][0] ),
    .I1(_3254_),
    .S(_3612_),
    .Z(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7624_ (.I(_3613_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7625_ (.I(_3610_),
    .Z(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7626_ (.I0(\reg_file.reg_storage[10][1] ),
    .I1(_3275_),
    .S(_3614_),
    .Z(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7627_ (.I(_3615_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7628_ (.I0(\reg_file.reg_storage[10][2] ),
    .I1(_3287_),
    .S(_3614_),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7629_ (.I(_3616_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7630_ (.I0(\reg_file.reg_storage[10][3] ),
    .I1(_3296_),
    .S(_3614_),
    .Z(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7631_ (.I(_3617_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7632_ (.I(_3611_),
    .Z(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7633_ (.I(_3618_),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7634_ (.I(_3614_),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7635_ (.A1(\reg_file.reg_storage[10][4] ),
    .A2(_3620_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7636_ (.A1(_3310_),
    .A2(_3619_),
    .B(_3621_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7637_ (.A1(\reg_file.reg_storage[10][5] ),
    .A2(_3620_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7638_ (.A1(_3319_),
    .A2(_3619_),
    .B(_3622_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7639_ (.A1(\reg_file.reg_storage[10][6] ),
    .A2(_3620_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7640_ (.A1(_3328_),
    .A2(_3619_),
    .B(_3623_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7641_ (.A1(\reg_file.reg_storage[10][7] ),
    .A2(_3620_),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7642_ (.A1(_3335_),
    .A2(_3619_),
    .B(_3624_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7643_ (.I(_3618_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7644_ (.I(_3610_),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7645_ (.I(_3626_),
    .Z(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7646_ (.A1(\reg_file.reg_storage[10][8] ),
    .A2(_3627_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7647_ (.A1(_3342_),
    .A2(_3625_),
    .B(_3628_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7648_ (.A1(\reg_file.reg_storage[10][9] ),
    .A2(_3627_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7649_ (.A1(_3349_),
    .A2(_3625_),
    .B(_3629_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7650_ (.A1(\reg_file.reg_storage[10][10] ),
    .A2(_3627_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7651_ (.A1(_3356_),
    .A2(_3625_),
    .B(_3630_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7652_ (.A1(\reg_file.reg_storage[10][11] ),
    .A2(_3627_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7653_ (.A1(_3362_),
    .A2(_3625_),
    .B(_3631_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7654_ (.I(_3618_),
    .Z(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7655_ (.I(_3626_),
    .Z(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7656_ (.A1(\reg_file.reg_storage[10][12] ),
    .A2(_3633_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7657_ (.A1(_3370_),
    .A2(_3632_),
    .B(_3634_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7658_ (.A1(\reg_file.reg_storage[10][13] ),
    .A2(_3633_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7659_ (.A1(_3377_),
    .A2(_3632_),
    .B(_3635_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7660_ (.A1(\reg_file.reg_storage[10][14] ),
    .A2(_3633_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7661_ (.A1(_3384_),
    .A2(_3632_),
    .B(_3636_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7662_ (.A1(\reg_file.reg_storage[10][15] ),
    .A2(_3633_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7663_ (.A1(_3391_),
    .A2(_3632_),
    .B(_3637_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7664_ (.I(_3618_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7665_ (.I(_3626_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7666_ (.A1(\reg_file.reg_storage[10][16] ),
    .A2(_3639_),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7667_ (.A1(_3399_),
    .A2(_3638_),
    .B(_3640_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7668_ (.A1(\reg_file.reg_storage[10][17] ),
    .A2(_3639_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7669_ (.A1(_3406_),
    .A2(_3638_),
    .B(_3641_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7670_ (.A1(\reg_file.reg_storage[10][18] ),
    .A2(_3639_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7671_ (.A1(_3412_),
    .A2(_3638_),
    .B(_3642_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7672_ (.A1(\reg_file.reg_storage[10][19] ),
    .A2(_3639_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7673_ (.A1(_3418_),
    .A2(_3638_),
    .B(_3643_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7674_ (.I(_3612_),
    .Z(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7675_ (.I(_3626_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7676_ (.A1(\reg_file.reg_storage[10][20] ),
    .A2(_3645_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7677_ (.A1(_3426_),
    .A2(_3644_),
    .B(_3646_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7678_ (.A1(\reg_file.reg_storage[10][21] ),
    .A2(_3645_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7679_ (.A1(_3433_),
    .A2(_3644_),
    .B(_3647_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7680_ (.A1(\reg_file.reg_storage[10][22] ),
    .A2(_3645_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7681_ (.A1(_3439_),
    .A2(_3644_),
    .B(_3648_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7682_ (.A1(\reg_file.reg_storage[10][23] ),
    .A2(_3645_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7683_ (.A1(_3445_),
    .A2(_3644_),
    .B(_3649_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7684_ (.I(_3612_),
    .Z(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7685_ (.I(_3611_),
    .Z(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7686_ (.A1(\reg_file.reg_storage[10][24] ),
    .A2(_3651_),
    .ZN(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7687_ (.A1(_3453_),
    .A2(_3650_),
    .B(_3652_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7688_ (.A1(\reg_file.reg_storage[10][25] ),
    .A2(_3651_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7689_ (.A1(_3460_),
    .A2(_3650_),
    .B(_3653_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7690_ (.A1(\reg_file.reg_storage[10][26] ),
    .A2(_3651_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7691_ (.A1(_3466_),
    .A2(_3650_),
    .B(_3654_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7692_ (.A1(\reg_file.reg_storage[10][27] ),
    .A2(_3651_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7693_ (.A1(_3472_),
    .A2(_3650_),
    .B(_3655_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7694_ (.I(_3612_),
    .Z(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7695_ (.I(_3611_),
    .Z(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7696_ (.A1(\reg_file.reg_storage[10][28] ),
    .A2(_3657_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7697_ (.A1(_3480_),
    .A2(_3656_),
    .B(_3658_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7698_ (.A1(\reg_file.reg_storage[10][29] ),
    .A2(_3657_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7699_ (.A1(_3486_),
    .A2(_3656_),
    .B(_3659_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7700_ (.A1(\reg_file.reg_storage[10][30] ),
    .A2(_3657_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7701_ (.A1(_3491_),
    .A2(_3656_),
    .B(_3660_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7702_ (.A1(\reg_file.reg_storage[10][31] ),
    .A2(_3657_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7703_ (.A1(_3496_),
    .A2(_3656_),
    .B(_3661_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7704_ (.I(_3252_),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7705_ (.A1(_3607_),
    .A2(_3553_),
    .A3(_3499_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7706_ (.I(_3663_),
    .Z(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7707_ (.I(_3664_),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7708_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(_3662_),
    .S(_3665_),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7709_ (.I(_3666_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7710_ (.I(_3273_),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7711_ (.I(_3663_),
    .Z(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7712_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(_3667_),
    .S(_3668_),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7713_ (.I(_3669_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7714_ (.I(_3285_),
    .Z(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7715_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(_3670_),
    .S(_3668_),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7716_ (.I(_3671_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7717_ (.I(_3294_),
    .Z(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7718_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(_3672_),
    .S(_3668_),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7719_ (.I(_3673_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7720_ (.I(_3309_),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7721_ (.I(_3674_),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7722_ (.I(_3664_),
    .Z(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7723_ (.I(_3676_),
    .Z(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7724_ (.I(_3668_),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7725_ (.A1(\reg_file.reg_storage[4][4] ),
    .A2(_3678_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7726_ (.A1(_3675_),
    .A2(_3677_),
    .B(_3679_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7727_ (.I(_3318_),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7728_ (.I(_3680_),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7729_ (.A1(\reg_file.reg_storage[4][5] ),
    .A2(_3678_),
    .ZN(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7730_ (.A1(_3681_),
    .A2(_3677_),
    .B(_3682_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7731_ (.I(_3327_),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7732_ (.I(_3683_),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7733_ (.A1(\reg_file.reg_storage[4][6] ),
    .A2(_3678_),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7734_ (.A1(_3684_),
    .A2(_3677_),
    .B(_3685_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7735_ (.I(_3334_),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7736_ (.I(_3686_),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7737_ (.A1(\reg_file.reg_storage[4][7] ),
    .A2(_3678_),
    .ZN(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7738_ (.A1(_3687_),
    .A2(_3677_),
    .B(_3688_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7739_ (.I(_3341_),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7740_ (.I(_3689_),
    .Z(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7741_ (.I(_3676_),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7742_ (.I(_3663_),
    .Z(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7743_ (.I(_3692_),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7744_ (.A1(\reg_file.reg_storage[4][8] ),
    .A2(_3693_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7745_ (.A1(_3690_),
    .A2(_3691_),
    .B(_3694_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7746_ (.I(_3348_),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7747_ (.I(_3695_),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7748_ (.A1(\reg_file.reg_storage[4][9] ),
    .A2(_3693_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7749_ (.A1(_3696_),
    .A2(_3691_),
    .B(_3697_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7750_ (.I(_3355_),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7751_ (.I(_3698_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7752_ (.A1(\reg_file.reg_storage[4][10] ),
    .A2(_3693_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7753_ (.A1(_3699_),
    .A2(_3691_),
    .B(_3700_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7754_ (.I(_3361_),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7755_ (.I(_3701_),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7756_ (.A1(\reg_file.reg_storage[4][11] ),
    .A2(_3693_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7757_ (.A1(_3702_),
    .A2(_3691_),
    .B(_3703_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7758_ (.I(_3369_),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7759_ (.I(_3704_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7760_ (.I(_3676_),
    .Z(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7761_ (.I(_3692_),
    .Z(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7762_ (.A1(\reg_file.reg_storage[4][12] ),
    .A2(_3707_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7763_ (.A1(_3705_),
    .A2(_3706_),
    .B(_3708_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7764_ (.I(_3376_),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7765_ (.I(_3709_),
    .Z(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7766_ (.A1(\reg_file.reg_storage[4][13] ),
    .A2(_3707_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7767_ (.A1(_3710_),
    .A2(_3706_),
    .B(_3711_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7768_ (.I(_3383_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7769_ (.I(_3712_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7770_ (.A1(\reg_file.reg_storage[4][14] ),
    .A2(_3707_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7771_ (.A1(_3713_),
    .A2(_3706_),
    .B(_3714_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7772_ (.I(_3390_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7773_ (.I(_3715_),
    .Z(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7774_ (.A1(\reg_file.reg_storage[4][15] ),
    .A2(_3707_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7775_ (.A1(_3716_),
    .A2(_3706_),
    .B(_3717_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7776_ (.I(_3398_),
    .Z(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7777_ (.I(_3718_),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7778_ (.I(_3676_),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7779_ (.I(_3692_),
    .Z(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7780_ (.A1(\reg_file.reg_storage[4][16] ),
    .A2(_3721_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7781_ (.A1(_3719_),
    .A2(_3720_),
    .B(_3722_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7782_ (.I(_3405_),
    .Z(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7783_ (.I(_3723_),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7784_ (.A1(\reg_file.reg_storage[4][17] ),
    .A2(_3721_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7785_ (.A1(_3724_),
    .A2(_3720_),
    .B(_3725_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7786_ (.I(_3411_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7787_ (.I(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7788_ (.A1(\reg_file.reg_storage[4][18] ),
    .A2(_3721_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7789_ (.A1(_3727_),
    .A2(_3720_),
    .B(_3728_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7790_ (.I(_3417_),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7791_ (.I(_3729_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7792_ (.A1(\reg_file.reg_storage[4][19] ),
    .A2(_3721_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7793_ (.A1(_3730_),
    .A2(_3720_),
    .B(_3731_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7794_ (.I(_3425_),
    .Z(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7795_ (.I(_3732_),
    .Z(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7796_ (.I(_3665_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7797_ (.I(_3692_),
    .Z(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7798_ (.A1(\reg_file.reg_storage[4][20] ),
    .A2(_3735_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7799_ (.A1(_3733_),
    .A2(_3734_),
    .B(_3736_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7800_ (.I(_3432_),
    .Z(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7801_ (.I(_3737_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7802_ (.A1(\reg_file.reg_storage[4][21] ),
    .A2(_3735_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7803_ (.A1(_3738_),
    .A2(_3734_),
    .B(_3739_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7804_ (.I(_3438_),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7805_ (.I(_3740_),
    .Z(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7806_ (.A1(\reg_file.reg_storage[4][22] ),
    .A2(_3735_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7807_ (.A1(_3741_),
    .A2(_3734_),
    .B(_3742_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7808_ (.I(_3444_),
    .Z(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7809_ (.I(_3743_),
    .Z(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7810_ (.A1(\reg_file.reg_storage[4][23] ),
    .A2(_3735_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7811_ (.A1(_3744_),
    .A2(_3734_),
    .B(_3745_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7812_ (.I(_3452_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7813_ (.I(_3746_),
    .Z(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7814_ (.I(_3665_),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7815_ (.I(_3664_),
    .Z(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7816_ (.A1(\reg_file.reg_storage[4][24] ),
    .A2(_3749_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7817_ (.A1(_3747_),
    .A2(_3748_),
    .B(_3750_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7818_ (.I(_3459_),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7819_ (.I(_3751_),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7820_ (.A1(\reg_file.reg_storage[4][25] ),
    .A2(_3749_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7821_ (.A1(_3752_),
    .A2(_3748_),
    .B(_3753_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7822_ (.I(_3465_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7823_ (.I(_3754_),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7824_ (.A1(\reg_file.reg_storage[4][26] ),
    .A2(_3749_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7825_ (.A1(_3755_),
    .A2(_3748_),
    .B(_3756_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7826_ (.I(_3471_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7827_ (.I(_3757_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7828_ (.A1(\reg_file.reg_storage[4][27] ),
    .A2(_3749_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7829_ (.A1(_3758_),
    .A2(_3748_),
    .B(_3759_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7830_ (.I(_3479_),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7831_ (.I(_3760_),
    .Z(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7832_ (.I(_3665_),
    .Z(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7833_ (.I(_3664_),
    .Z(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7834_ (.A1(\reg_file.reg_storage[4][28] ),
    .A2(_3763_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7835_ (.A1(_3761_),
    .A2(_3762_),
    .B(_3764_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7836_ (.I(_3485_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7837_ (.I(_3765_),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7838_ (.A1(\reg_file.reg_storage[4][29] ),
    .A2(_3763_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7839_ (.A1(_3766_),
    .A2(_3762_),
    .B(_3767_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7840_ (.I(_3490_),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7841_ (.I(_3768_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7842_ (.A1(\reg_file.reg_storage[4][30] ),
    .A2(_3763_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7843_ (.A1(_3769_),
    .A2(_3762_),
    .B(_3770_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7844_ (.I(_3495_),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7845_ (.I(_3771_),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7846_ (.A1(\reg_file.reg_storage[4][31] ),
    .A2(_3763_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7847_ (.A1(_3772_),
    .A2(_3762_),
    .B(_3773_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7848_ (.A1(_3255_),
    .A2(_3256_),
    .A3(_3263_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7849_ (.I(net32),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7850_ (.A1(net2),
    .A2(_3775_),
    .ZN(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7851_ (.A1(_3774_),
    .A2(_3776_),
    .ZN(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7852_ (.I(_3777_),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7853_ (.I(_3778_),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7854_ (.I0(\reg_file.reg_storage[15][0] ),
    .I1(_3662_),
    .S(_3779_),
    .Z(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7855_ (.I(_3780_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7856_ (.I(_3777_),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7857_ (.I0(\reg_file.reg_storage[15][1] ),
    .I1(_3667_),
    .S(_3781_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7858_ (.I(_3782_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7859_ (.I0(\reg_file.reg_storage[15][2] ),
    .I1(_3670_),
    .S(_3781_),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7860_ (.I(_3783_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7861_ (.I0(\reg_file.reg_storage[15][3] ),
    .I1(_3672_),
    .S(_3781_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7862_ (.I(_3784_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7863_ (.I(_3778_),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7864_ (.I(_3785_),
    .Z(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7865_ (.I(_3781_),
    .Z(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7866_ (.A1(\reg_file.reg_storage[15][4] ),
    .A2(_3787_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7867_ (.A1(_3675_),
    .A2(_3786_),
    .B(_3788_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7868_ (.A1(\reg_file.reg_storage[15][5] ),
    .A2(_3787_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7869_ (.A1(_3681_),
    .A2(_3786_),
    .B(_3789_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7870_ (.A1(\reg_file.reg_storage[15][6] ),
    .A2(_3787_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7871_ (.A1(_3684_),
    .A2(_3786_),
    .B(_3790_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7872_ (.A1(\reg_file.reg_storage[15][7] ),
    .A2(_3787_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7873_ (.A1(_3687_),
    .A2(_3786_),
    .B(_3791_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7874_ (.I(_3785_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7875_ (.I(_3777_),
    .Z(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7876_ (.I(_3793_),
    .Z(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7877_ (.A1(\reg_file.reg_storage[15][8] ),
    .A2(_3794_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7878_ (.A1(_3690_),
    .A2(_3792_),
    .B(_3795_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7879_ (.A1(\reg_file.reg_storage[15][9] ),
    .A2(_3794_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7880_ (.A1(_3696_),
    .A2(_3792_),
    .B(_3796_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7881_ (.A1(\reg_file.reg_storage[15][10] ),
    .A2(_3794_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7882_ (.A1(_3699_),
    .A2(_3792_),
    .B(_3797_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7883_ (.A1(\reg_file.reg_storage[15][11] ),
    .A2(_3794_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7884_ (.A1(_3702_),
    .A2(_3792_),
    .B(_3798_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7885_ (.I(_3785_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7886_ (.I(_3793_),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7887_ (.A1(\reg_file.reg_storage[15][12] ),
    .A2(_3800_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7888_ (.A1(_3705_),
    .A2(_3799_),
    .B(_3801_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7889_ (.A1(\reg_file.reg_storage[15][13] ),
    .A2(_3800_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7890_ (.A1(_3710_),
    .A2(_3799_),
    .B(_3802_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7891_ (.A1(\reg_file.reg_storage[15][14] ),
    .A2(_3800_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7892_ (.A1(_3713_),
    .A2(_3799_),
    .B(_3803_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7893_ (.A1(\reg_file.reg_storage[15][15] ),
    .A2(_3800_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7894_ (.A1(_3716_),
    .A2(_3799_),
    .B(_3804_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7895_ (.I(_3785_),
    .Z(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7896_ (.I(_3793_),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7897_ (.A1(\reg_file.reg_storage[15][16] ),
    .A2(_3806_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7898_ (.A1(_3719_),
    .A2(_3805_),
    .B(_3807_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7899_ (.A1(\reg_file.reg_storage[15][17] ),
    .A2(_3806_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7900_ (.A1(_3724_),
    .A2(_3805_),
    .B(_3808_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7901_ (.A1(\reg_file.reg_storage[15][18] ),
    .A2(_3806_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7902_ (.A1(_3727_),
    .A2(_3805_),
    .B(_3809_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7903_ (.A1(\reg_file.reg_storage[15][19] ),
    .A2(_3806_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7904_ (.A1(_3730_),
    .A2(_3805_),
    .B(_3810_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7905_ (.I(_3779_),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7906_ (.I(_3793_),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7907_ (.A1(\reg_file.reg_storage[15][20] ),
    .A2(_3812_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7908_ (.A1(_3733_),
    .A2(_3811_),
    .B(_3813_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7909_ (.A1(\reg_file.reg_storage[15][21] ),
    .A2(_3812_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7910_ (.A1(_3738_),
    .A2(_3811_),
    .B(_3814_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7911_ (.A1(\reg_file.reg_storage[15][22] ),
    .A2(_3812_),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7912_ (.A1(_3741_),
    .A2(_3811_),
    .B(_3815_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7913_ (.A1(\reg_file.reg_storage[15][23] ),
    .A2(_3812_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7914_ (.A1(_3744_),
    .A2(_3811_),
    .B(_3816_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7915_ (.I(_3779_),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7916_ (.I(_3778_),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7917_ (.A1(\reg_file.reg_storage[15][24] ),
    .A2(_3818_),
    .ZN(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7918_ (.A1(_3747_),
    .A2(_3817_),
    .B(_3819_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7919_ (.A1(\reg_file.reg_storage[15][25] ),
    .A2(_3818_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7920_ (.A1(_3752_),
    .A2(_3817_),
    .B(_3820_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7921_ (.A1(\reg_file.reg_storage[15][26] ),
    .A2(_3818_),
    .ZN(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7922_ (.A1(_3755_),
    .A2(_3817_),
    .B(_3821_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7923_ (.A1(\reg_file.reg_storage[15][27] ),
    .A2(_3818_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7924_ (.A1(_3758_),
    .A2(_3817_),
    .B(_3822_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7925_ (.I(_3779_),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7926_ (.I(_3778_),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7927_ (.A1(\reg_file.reg_storage[15][28] ),
    .A2(_3824_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7928_ (.A1(_3761_),
    .A2(_3823_),
    .B(_3825_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7929_ (.A1(\reg_file.reg_storage[15][29] ),
    .A2(_3824_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7930_ (.A1(_3766_),
    .A2(_3823_),
    .B(_3826_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7931_ (.A1(\reg_file.reg_storage[15][30] ),
    .A2(_3824_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7932_ (.A1(_3769_),
    .A2(_3823_),
    .B(_3827_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7933_ (.A1(\reg_file.reg_storage[15][31] ),
    .A2(_3824_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7934_ (.A1(_3772_),
    .A2(_3823_),
    .B(_3828_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7935_ (.A1(_3255_),
    .A2(_3608_),
    .A3(_3263_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7936_ (.A1(_3258_),
    .A2(_3775_),
    .A3(_3829_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7937_ (.I(_3830_),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7938_ (.I(_3831_),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7939_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(_3662_),
    .S(_3832_),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7940_ (.I(_3833_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7941_ (.I(_3830_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7942_ (.I0(\reg_file.reg_storage[2][1] ),
    .I1(_3667_),
    .S(_3834_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7943_ (.I(_3835_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7944_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(_3670_),
    .S(_3834_),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7945_ (.I(_3836_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7946_ (.I0(\reg_file.reg_storage[2][3] ),
    .I1(_3672_),
    .S(_3834_),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7947_ (.I(_3837_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7948_ (.I(_3831_),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7949_ (.I(_3838_),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7950_ (.I(_3834_),
    .Z(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7951_ (.A1(\reg_file.reg_storage[2][4] ),
    .A2(_3840_),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7952_ (.A1(_3675_),
    .A2(_3839_),
    .B(_3841_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7953_ (.A1(\reg_file.reg_storage[2][5] ),
    .A2(_3840_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7954_ (.A1(_3681_),
    .A2(_3839_),
    .B(_3842_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7955_ (.A1(\reg_file.reg_storage[2][6] ),
    .A2(_3840_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7956_ (.A1(_3684_),
    .A2(_3839_),
    .B(_3843_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7957_ (.A1(\reg_file.reg_storage[2][7] ),
    .A2(_3840_),
    .ZN(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7958_ (.A1(_3687_),
    .A2(_3839_),
    .B(_3844_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7959_ (.I(_3838_),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7960_ (.I(_3830_),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7961_ (.I(_3846_),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7962_ (.A1(\reg_file.reg_storage[2][8] ),
    .A2(_3847_),
    .ZN(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7963_ (.A1(_3690_),
    .A2(_3845_),
    .B(_3848_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7964_ (.A1(\reg_file.reg_storage[2][9] ),
    .A2(_3847_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7965_ (.A1(_3696_),
    .A2(_3845_),
    .B(_3849_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7966_ (.A1(\reg_file.reg_storage[2][10] ),
    .A2(_3847_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7967_ (.A1(_3699_),
    .A2(_3845_),
    .B(_3850_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7968_ (.A1(\reg_file.reg_storage[2][11] ),
    .A2(_3847_),
    .ZN(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7969_ (.A1(_3702_),
    .A2(_3845_),
    .B(_3851_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7970_ (.I(_3838_),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7971_ (.I(_3846_),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7972_ (.A1(\reg_file.reg_storage[2][12] ),
    .A2(_3853_),
    .ZN(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7973_ (.A1(_3705_),
    .A2(_3852_),
    .B(_3854_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7974_ (.A1(\reg_file.reg_storage[2][13] ),
    .A2(_3853_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7975_ (.A1(_3710_),
    .A2(_3852_),
    .B(_3855_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7976_ (.A1(\reg_file.reg_storage[2][14] ),
    .A2(_3853_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7977_ (.A1(_3713_),
    .A2(_3852_),
    .B(_3856_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7978_ (.A1(\reg_file.reg_storage[2][15] ),
    .A2(_3853_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7979_ (.A1(_3716_),
    .A2(_3852_),
    .B(_3857_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7980_ (.I(_3838_),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7981_ (.I(_3846_),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7982_ (.A1(\reg_file.reg_storage[2][16] ),
    .A2(_3859_),
    .ZN(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7983_ (.A1(_3719_),
    .A2(_3858_),
    .B(_3860_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7984_ (.A1(\reg_file.reg_storage[2][17] ),
    .A2(_3859_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7985_ (.A1(_3724_),
    .A2(_3858_),
    .B(_3861_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7986_ (.A1(\reg_file.reg_storage[2][18] ),
    .A2(_3859_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7987_ (.A1(_3727_),
    .A2(_3858_),
    .B(_3862_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7988_ (.A1(\reg_file.reg_storage[2][19] ),
    .A2(_3859_),
    .ZN(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7989_ (.A1(_3730_),
    .A2(_3858_),
    .B(_3863_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7990_ (.I(_3832_),
    .Z(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7991_ (.I(_3846_),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7992_ (.A1(\reg_file.reg_storage[2][20] ),
    .A2(_3865_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7993_ (.A1(_3733_),
    .A2(_3864_),
    .B(_3866_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7994_ (.A1(\reg_file.reg_storage[2][21] ),
    .A2(_3865_),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7995_ (.A1(_3738_),
    .A2(_3864_),
    .B(_3867_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7996_ (.A1(\reg_file.reg_storage[2][22] ),
    .A2(_3865_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7997_ (.A1(_3741_),
    .A2(_3864_),
    .B(_3868_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7998_ (.A1(\reg_file.reg_storage[2][23] ),
    .A2(_3865_),
    .ZN(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7999_ (.A1(_3744_),
    .A2(_3864_),
    .B(_3869_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8000_ (.I(_3832_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8001_ (.I(_3831_),
    .Z(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8002_ (.A1(\reg_file.reg_storage[2][24] ),
    .A2(_3871_),
    .ZN(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8003_ (.A1(_3747_),
    .A2(_3870_),
    .B(_3872_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8004_ (.A1(\reg_file.reg_storage[2][25] ),
    .A2(_3871_),
    .ZN(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8005_ (.A1(_3752_),
    .A2(_3870_),
    .B(_3873_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8006_ (.A1(\reg_file.reg_storage[2][26] ),
    .A2(_3871_),
    .ZN(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8007_ (.A1(_3755_),
    .A2(_3870_),
    .B(_3874_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8008_ (.A1(\reg_file.reg_storage[2][27] ),
    .A2(_3871_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8009_ (.A1(_3758_),
    .A2(_3870_),
    .B(_3875_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8010_ (.I(_3832_),
    .Z(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8011_ (.I(_3831_),
    .Z(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8012_ (.A1(\reg_file.reg_storage[2][28] ),
    .A2(_3877_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8013_ (.A1(_3761_),
    .A2(_3876_),
    .B(_3878_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8014_ (.A1(\reg_file.reg_storage[2][29] ),
    .A2(_3877_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8015_ (.A1(_3766_),
    .A2(_3876_),
    .B(_3879_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8016_ (.A1(\reg_file.reg_storage[2][30] ),
    .A2(_3877_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8017_ (.A1(_3769_),
    .A2(_3876_),
    .B(_3880_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8018_ (.A1(\reg_file.reg_storage[2][31] ),
    .A2(_3877_),
    .ZN(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8019_ (.A1(_3772_),
    .A2(_3876_),
    .B(_3881_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8020_ (.A1(_3607_),
    .A2(_3553_),
    .A3(_3498_),
    .A4(_3776_),
    .ZN(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8021_ (.I(_3882_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8022_ (.I(_3883_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8023_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(_3662_),
    .S(_3884_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8024_ (.I(_3885_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8025_ (.I(_3882_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8026_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(_3667_),
    .S(_3886_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8027_ (.I(_3887_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8028_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(_3670_),
    .S(_3886_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8029_ (.I(_3888_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8030_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(_3672_),
    .S(_3886_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8031_ (.I(_3889_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8032_ (.I(_3883_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8033_ (.I(_3890_),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8034_ (.I(_3886_),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8035_ (.A1(\reg_file.reg_storage[12][4] ),
    .A2(_3892_),
    .ZN(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8036_ (.A1(_3675_),
    .A2(_3891_),
    .B(_3893_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8037_ (.A1(\reg_file.reg_storage[12][5] ),
    .A2(_3892_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8038_ (.A1(_3681_),
    .A2(_3891_),
    .B(_3894_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8039_ (.A1(\reg_file.reg_storage[12][6] ),
    .A2(_3892_),
    .ZN(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8040_ (.A1(_3684_),
    .A2(_3891_),
    .B(_3895_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8041_ (.A1(\reg_file.reg_storage[12][7] ),
    .A2(_3892_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8042_ (.A1(_3687_),
    .A2(_3891_),
    .B(_3896_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8043_ (.I(_3890_),
    .Z(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8044_ (.I(_3882_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8045_ (.I(_3898_),
    .Z(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8046_ (.A1(\reg_file.reg_storage[12][8] ),
    .A2(_3899_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8047_ (.A1(_3690_),
    .A2(_3897_),
    .B(_3900_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8048_ (.A1(\reg_file.reg_storage[12][9] ),
    .A2(_3899_),
    .ZN(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8049_ (.A1(_3696_),
    .A2(_3897_),
    .B(_3901_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8050_ (.A1(\reg_file.reg_storage[12][10] ),
    .A2(_3899_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8051_ (.A1(_3699_),
    .A2(_3897_),
    .B(_3902_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8052_ (.A1(\reg_file.reg_storage[12][11] ),
    .A2(_3899_),
    .ZN(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8053_ (.A1(_3702_),
    .A2(_3897_),
    .B(_3903_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8054_ (.I(_3890_),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8055_ (.I(_3898_),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8056_ (.A1(\reg_file.reg_storage[12][12] ),
    .A2(_3905_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8057_ (.A1(_3705_),
    .A2(_3904_),
    .B(_3906_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8058_ (.A1(\reg_file.reg_storage[12][13] ),
    .A2(_3905_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8059_ (.A1(_3710_),
    .A2(_3904_),
    .B(_3907_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8060_ (.A1(\reg_file.reg_storage[12][14] ),
    .A2(_3905_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8061_ (.A1(_3713_),
    .A2(_3904_),
    .B(_3908_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8062_ (.A1(\reg_file.reg_storage[12][15] ),
    .A2(_3905_),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8063_ (.A1(_3716_),
    .A2(_3904_),
    .B(_3909_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8064_ (.I(_3890_),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8065_ (.I(_3898_),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8066_ (.A1(\reg_file.reg_storage[12][16] ),
    .A2(_3911_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8067_ (.A1(_3719_),
    .A2(_3910_),
    .B(_3912_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8068_ (.A1(\reg_file.reg_storage[12][17] ),
    .A2(_3911_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8069_ (.A1(_3724_),
    .A2(_3910_),
    .B(_3913_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8070_ (.A1(\reg_file.reg_storage[12][18] ),
    .A2(_3911_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8071_ (.A1(_3727_),
    .A2(_3910_),
    .B(_3914_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8072_ (.A1(\reg_file.reg_storage[12][19] ),
    .A2(_3911_),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8073_ (.A1(_3730_),
    .A2(_3910_),
    .B(_3915_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8074_ (.I(_3884_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8075_ (.I(_3898_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8076_ (.A1(\reg_file.reg_storage[12][20] ),
    .A2(_3917_),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8077_ (.A1(_3733_),
    .A2(_3916_),
    .B(_3918_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8078_ (.A1(\reg_file.reg_storage[12][21] ),
    .A2(_3917_),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8079_ (.A1(_3738_),
    .A2(_3916_),
    .B(_3919_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8080_ (.A1(\reg_file.reg_storage[12][22] ),
    .A2(_3917_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8081_ (.A1(_3741_),
    .A2(_3916_),
    .B(_3920_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8082_ (.A1(\reg_file.reg_storage[12][23] ),
    .A2(_3917_),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8083_ (.A1(_3744_),
    .A2(_3916_),
    .B(_3921_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8084_ (.I(_3884_),
    .Z(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8085_ (.I(_3883_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8086_ (.A1(\reg_file.reg_storage[12][24] ),
    .A2(_3923_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8087_ (.A1(_3747_),
    .A2(_3922_),
    .B(_3924_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8088_ (.A1(\reg_file.reg_storage[12][25] ),
    .A2(_3923_),
    .ZN(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8089_ (.A1(_3752_),
    .A2(_3922_),
    .B(_3925_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8090_ (.A1(\reg_file.reg_storage[12][26] ),
    .A2(_3923_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8091_ (.A1(_3755_),
    .A2(_3922_),
    .B(_3926_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8092_ (.A1(\reg_file.reg_storage[12][27] ),
    .A2(_3923_),
    .ZN(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8093_ (.A1(_3758_),
    .A2(_3922_),
    .B(_3927_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8094_ (.I(_3884_),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8095_ (.I(_3883_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8096_ (.A1(\reg_file.reg_storage[12][28] ),
    .A2(_3929_),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8097_ (.A1(_3761_),
    .A2(_3928_),
    .B(_3930_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8098_ (.A1(\reg_file.reg_storage[12][29] ),
    .A2(_3929_),
    .ZN(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8099_ (.A1(_3766_),
    .A2(_3928_),
    .B(_3931_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8100_ (.A1(\reg_file.reg_storage[12][30] ),
    .A2(_3929_),
    .ZN(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8101_ (.A1(_3769_),
    .A2(_3928_),
    .B(_3932_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8102_ (.A1(\reg_file.reg_storage[12][31] ),
    .A2(_3929_),
    .ZN(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8103_ (.A1(_3772_),
    .A2(_3928_),
    .B(_3933_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8104_ (.I(_3252_),
    .Z(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8105_ (.A1(_3552_),
    .A2(_3256_),
    .A3(_3263_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8106_ (.A1(_3776_),
    .A2(_3935_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8107_ (.I(_3936_),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8108_ (.I(_3937_),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8109_ (.I0(\reg_file.reg_storage[13][0] ),
    .I1(_3934_),
    .S(_3938_),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8110_ (.I(_3939_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8111_ (.I(_3273_),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8112_ (.I(_3936_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8113_ (.I0(\reg_file.reg_storage[13][1] ),
    .I1(_3940_),
    .S(_3941_),
    .Z(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8114_ (.I(_3942_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8115_ (.I(_3285_),
    .Z(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8116_ (.I0(\reg_file.reg_storage[13][2] ),
    .I1(_3943_),
    .S(_3941_),
    .Z(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8117_ (.I(_3944_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8118_ (.I(_3294_),
    .Z(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8119_ (.I0(\reg_file.reg_storage[13][3] ),
    .I1(_3945_),
    .S(_3941_),
    .Z(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8120_ (.I(_3946_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8121_ (.I(_3309_),
    .Z(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8122_ (.I(_3937_),
    .Z(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8123_ (.I(_3948_),
    .Z(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8124_ (.I(_3941_),
    .Z(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8125_ (.A1(\reg_file.reg_storage[13][4] ),
    .A2(_3950_),
    .ZN(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8126_ (.A1(_3947_),
    .A2(_3949_),
    .B(_3951_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8127_ (.I(_3318_),
    .Z(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8128_ (.A1(\reg_file.reg_storage[13][5] ),
    .A2(_3950_),
    .ZN(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8129_ (.A1(_3952_),
    .A2(_3949_),
    .B(_3953_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8130_ (.I(_3327_),
    .Z(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8131_ (.A1(\reg_file.reg_storage[13][6] ),
    .A2(_3950_),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8132_ (.A1(_3954_),
    .A2(_3949_),
    .B(_3955_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8133_ (.I(_3334_),
    .Z(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8134_ (.A1(\reg_file.reg_storage[13][7] ),
    .A2(_3950_),
    .ZN(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8135_ (.A1(_3956_),
    .A2(_3949_),
    .B(_3957_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8136_ (.I(_3341_),
    .Z(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8137_ (.I(_3948_),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8138_ (.I(_3936_),
    .Z(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8139_ (.I(_3960_),
    .Z(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8140_ (.A1(\reg_file.reg_storage[13][8] ),
    .A2(_3961_),
    .ZN(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8141_ (.A1(_3958_),
    .A2(_3959_),
    .B(_3962_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8142_ (.I(_3348_),
    .Z(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8143_ (.A1(\reg_file.reg_storage[13][9] ),
    .A2(_3961_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8144_ (.A1(_3963_),
    .A2(_3959_),
    .B(_3964_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8145_ (.I(_3355_),
    .Z(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8146_ (.A1(\reg_file.reg_storage[13][10] ),
    .A2(_3961_),
    .ZN(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8147_ (.A1(_3965_),
    .A2(_3959_),
    .B(_3966_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8148_ (.I(_3361_),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8149_ (.A1(\reg_file.reg_storage[13][11] ),
    .A2(_3961_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8150_ (.A1(_3967_),
    .A2(_3959_),
    .B(_3968_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8151_ (.I(_3369_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8152_ (.I(_3948_),
    .Z(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8153_ (.I(_3960_),
    .Z(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8154_ (.A1(\reg_file.reg_storage[13][12] ),
    .A2(_3971_),
    .ZN(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8155_ (.A1(_3969_),
    .A2(_3970_),
    .B(_3972_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8156_ (.I(_3376_),
    .Z(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8157_ (.A1(\reg_file.reg_storage[13][13] ),
    .A2(_3971_),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8158_ (.A1(_3973_),
    .A2(_3970_),
    .B(_3974_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8159_ (.I(_3383_),
    .Z(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8160_ (.A1(\reg_file.reg_storage[13][14] ),
    .A2(_3971_),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8161_ (.A1(_3975_),
    .A2(_3970_),
    .B(_3976_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8162_ (.I(_3390_),
    .Z(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8163_ (.A1(\reg_file.reg_storage[13][15] ),
    .A2(_3971_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8164_ (.A1(_3977_),
    .A2(_3970_),
    .B(_3978_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8165_ (.I(_3398_),
    .Z(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8166_ (.I(_3948_),
    .Z(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8167_ (.I(_3960_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8168_ (.A1(\reg_file.reg_storage[13][16] ),
    .A2(_3981_),
    .ZN(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8169_ (.A1(_3979_),
    .A2(_3980_),
    .B(_3982_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8170_ (.I(_3405_),
    .Z(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8171_ (.A1(\reg_file.reg_storage[13][17] ),
    .A2(_3981_),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8172_ (.A1(_3983_),
    .A2(_3980_),
    .B(_3984_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8173_ (.I(_3411_),
    .Z(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8174_ (.A1(\reg_file.reg_storage[13][18] ),
    .A2(_3981_),
    .ZN(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8175_ (.A1(_3985_),
    .A2(_3980_),
    .B(_3986_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8176_ (.I(_3417_),
    .Z(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8177_ (.A1(\reg_file.reg_storage[13][19] ),
    .A2(_3981_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8178_ (.A1(_3987_),
    .A2(_3980_),
    .B(_3988_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8179_ (.I(_3425_),
    .Z(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8180_ (.I(_3938_),
    .Z(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8181_ (.I(_3960_),
    .Z(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8182_ (.A1(\reg_file.reg_storage[13][20] ),
    .A2(_3991_),
    .ZN(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8183_ (.A1(_3989_),
    .A2(_3990_),
    .B(_3992_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8184_ (.I(_3432_),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8185_ (.A1(\reg_file.reg_storage[13][21] ),
    .A2(_3991_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8186_ (.A1(_3993_),
    .A2(_3990_),
    .B(_3994_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8187_ (.I(_3438_),
    .Z(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8188_ (.A1(\reg_file.reg_storage[13][22] ),
    .A2(_3991_),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8189_ (.A1(_3995_),
    .A2(_3990_),
    .B(_3996_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8190_ (.I(_3444_),
    .Z(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8191_ (.A1(\reg_file.reg_storage[13][23] ),
    .A2(_3991_),
    .ZN(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8192_ (.A1(_3997_),
    .A2(_3990_),
    .B(_3998_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8193_ (.I(_3452_),
    .Z(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8194_ (.I(_3938_),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8195_ (.I(_3937_),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8196_ (.A1(\reg_file.reg_storage[13][24] ),
    .A2(_4001_),
    .ZN(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8197_ (.A1(_3999_),
    .A2(_4000_),
    .B(_4002_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8198_ (.I(_3459_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8199_ (.A1(\reg_file.reg_storage[13][25] ),
    .A2(_4001_),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8200_ (.A1(_4003_),
    .A2(_4000_),
    .B(_4004_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8201_ (.I(_3465_),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8202_ (.A1(\reg_file.reg_storage[13][26] ),
    .A2(_4001_),
    .ZN(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8203_ (.A1(_4005_),
    .A2(_4000_),
    .B(_4006_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8204_ (.I(_3471_),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8205_ (.A1(\reg_file.reg_storage[13][27] ),
    .A2(_4001_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8206_ (.A1(_4007_),
    .A2(_4000_),
    .B(_4008_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8207_ (.I(_3479_),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8208_ (.I(_3938_),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8209_ (.I(_3937_),
    .Z(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8210_ (.A1(\reg_file.reg_storage[13][28] ),
    .A2(_4011_),
    .ZN(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8211_ (.A1(_4009_),
    .A2(_4010_),
    .B(_4012_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8212_ (.I(_3485_),
    .Z(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8213_ (.A1(\reg_file.reg_storage[13][29] ),
    .A2(_4011_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8214_ (.A1(_4013_),
    .A2(_4010_),
    .B(_4014_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8215_ (.I(_3490_),
    .Z(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8216_ (.A1(\reg_file.reg_storage[13][30] ),
    .A2(_4011_),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8217_ (.A1(_4015_),
    .A2(_4010_),
    .B(_4016_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8218_ (.I(_3495_),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8219_ (.A1(\reg_file.reg_storage[13][31] ),
    .A2(_4011_),
    .ZN(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8220_ (.A1(_4017_),
    .A2(_4010_),
    .B(_4018_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8221_ (.A1(_3776_),
    .A2(_3829_),
    .ZN(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8222_ (.I(_4019_),
    .Z(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8223_ (.I(_4020_),
    .Z(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8224_ (.I0(\reg_file.reg_storage[14][0] ),
    .I1(_3934_),
    .S(_4021_),
    .Z(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8225_ (.I(_4022_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8226_ (.I(_4019_),
    .Z(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8227_ (.I0(\reg_file.reg_storage[14][1] ),
    .I1(_3940_),
    .S(_4023_),
    .Z(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8228_ (.I(_4024_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8229_ (.I0(\reg_file.reg_storage[14][2] ),
    .I1(_3943_),
    .S(_4023_),
    .Z(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8230_ (.I(_4025_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8231_ (.I0(\reg_file.reg_storage[14][3] ),
    .I1(_3945_),
    .S(_4023_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8232_ (.I(_4026_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8233_ (.I(_4020_),
    .Z(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8234_ (.I(_4027_),
    .Z(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8235_ (.I(_4023_),
    .Z(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8236_ (.A1(\reg_file.reg_storage[14][4] ),
    .A2(_4029_),
    .ZN(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8237_ (.A1(_3947_),
    .A2(_4028_),
    .B(_4030_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8238_ (.A1(\reg_file.reg_storage[14][5] ),
    .A2(_4029_),
    .ZN(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8239_ (.A1(_3952_),
    .A2(_4028_),
    .B(_4031_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8240_ (.A1(\reg_file.reg_storage[14][6] ),
    .A2(_4029_),
    .ZN(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8241_ (.A1(_3954_),
    .A2(_4028_),
    .B(_4032_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8242_ (.A1(\reg_file.reg_storage[14][7] ),
    .A2(_4029_),
    .ZN(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8243_ (.A1(_3956_),
    .A2(_4028_),
    .B(_4033_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8244_ (.I(_4027_),
    .Z(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8245_ (.I(_4019_),
    .Z(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8246_ (.I(_4035_),
    .Z(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8247_ (.A1(\reg_file.reg_storage[14][8] ),
    .A2(_4036_),
    .ZN(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8248_ (.A1(_3958_),
    .A2(_4034_),
    .B(_4037_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8249_ (.A1(\reg_file.reg_storage[14][9] ),
    .A2(_4036_),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8250_ (.A1(_3963_),
    .A2(_4034_),
    .B(_4038_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8251_ (.A1(\reg_file.reg_storage[14][10] ),
    .A2(_4036_),
    .ZN(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8252_ (.A1(_3965_),
    .A2(_4034_),
    .B(_4039_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8253_ (.A1(\reg_file.reg_storage[14][11] ),
    .A2(_4036_),
    .ZN(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8254_ (.A1(_3967_),
    .A2(_4034_),
    .B(_4040_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8255_ (.I(_4027_),
    .Z(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8256_ (.I(_4035_),
    .Z(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8257_ (.A1(\reg_file.reg_storage[14][12] ),
    .A2(_4042_),
    .ZN(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8258_ (.A1(_3969_),
    .A2(_4041_),
    .B(_4043_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8259_ (.A1(\reg_file.reg_storage[14][13] ),
    .A2(_4042_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8260_ (.A1(_3973_),
    .A2(_4041_),
    .B(_4044_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8261_ (.A1(\reg_file.reg_storage[14][14] ),
    .A2(_4042_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8262_ (.A1(_3975_),
    .A2(_4041_),
    .B(_4045_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8263_ (.A1(\reg_file.reg_storage[14][15] ),
    .A2(_4042_),
    .ZN(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8264_ (.A1(_3977_),
    .A2(_4041_),
    .B(_4046_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8265_ (.I(_4027_),
    .Z(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8266_ (.I(_4035_),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8267_ (.A1(\reg_file.reg_storage[14][16] ),
    .A2(_4048_),
    .ZN(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8268_ (.A1(_3979_),
    .A2(_4047_),
    .B(_4049_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8269_ (.A1(\reg_file.reg_storage[14][17] ),
    .A2(_4048_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8270_ (.A1(_3983_),
    .A2(_4047_),
    .B(_4050_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8271_ (.A1(\reg_file.reg_storage[14][18] ),
    .A2(_4048_),
    .ZN(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8272_ (.A1(_3985_),
    .A2(_4047_),
    .B(_4051_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8273_ (.A1(\reg_file.reg_storage[14][19] ),
    .A2(_4048_),
    .ZN(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8274_ (.A1(_3987_),
    .A2(_4047_),
    .B(_4052_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8275_ (.I(_4021_),
    .Z(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8276_ (.I(_4035_),
    .Z(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8277_ (.A1(\reg_file.reg_storage[14][20] ),
    .A2(_4054_),
    .ZN(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8278_ (.A1(_3989_),
    .A2(_4053_),
    .B(_4055_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8279_ (.A1(\reg_file.reg_storage[14][21] ),
    .A2(_4054_),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8280_ (.A1(_3993_),
    .A2(_4053_),
    .B(_4056_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8281_ (.A1(\reg_file.reg_storage[14][22] ),
    .A2(_4054_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8282_ (.A1(_3995_),
    .A2(_4053_),
    .B(_4057_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8283_ (.A1(\reg_file.reg_storage[14][23] ),
    .A2(_4054_),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8284_ (.A1(_3997_),
    .A2(_4053_),
    .B(_4058_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8285_ (.I(_4021_),
    .Z(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8286_ (.I(_4020_),
    .Z(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8287_ (.A1(\reg_file.reg_storage[14][24] ),
    .A2(_4060_),
    .ZN(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8288_ (.A1(_3999_),
    .A2(_4059_),
    .B(_4061_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8289_ (.A1(\reg_file.reg_storage[14][25] ),
    .A2(_4060_),
    .ZN(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8290_ (.A1(_4003_),
    .A2(_4059_),
    .B(_4062_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8291_ (.A1(\reg_file.reg_storage[14][26] ),
    .A2(_4060_),
    .ZN(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8292_ (.A1(_4005_),
    .A2(_4059_),
    .B(_4063_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8293_ (.A1(\reg_file.reg_storage[14][27] ),
    .A2(_4060_),
    .ZN(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8294_ (.A1(_4007_),
    .A2(_4059_),
    .B(_4064_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8295_ (.I(_4021_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8296_ (.I(_4020_),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8297_ (.A1(\reg_file.reg_storage[14][28] ),
    .A2(_4066_),
    .ZN(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8298_ (.A1(_4009_),
    .A2(_4065_),
    .B(_4067_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8299_ (.A1(\reg_file.reg_storage[14][29] ),
    .A2(_4066_),
    .ZN(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8300_ (.A1(_4013_),
    .A2(_4065_),
    .B(_4068_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8301_ (.A1(\reg_file.reg_storage[14][30] ),
    .A2(_4066_),
    .ZN(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8302_ (.A1(_4015_),
    .A2(_4065_),
    .B(_4069_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8303_ (.A1(\reg_file.reg_storage[14][31] ),
    .A2(_4066_),
    .ZN(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8304_ (.A1(_4017_),
    .A2(_4065_),
    .B(_4070_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8305_ (.A1(_3499_),
    .A2(_3609_),
    .ZN(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8306_ (.I(_4071_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8307_ (.I(_4072_),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8308_ (.I0(\reg_file.reg_storage[6][0] ),
    .I1(_3934_),
    .S(_4073_),
    .Z(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8309_ (.I(_4074_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8310_ (.I(_4071_),
    .Z(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8311_ (.I0(\reg_file.reg_storage[6][1] ),
    .I1(_3940_),
    .S(_4075_),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8312_ (.I(_4076_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8313_ (.I0(\reg_file.reg_storage[6][2] ),
    .I1(_3943_),
    .S(_4075_),
    .Z(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8314_ (.I(_4077_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8315_ (.I0(\reg_file.reg_storage[6][3] ),
    .I1(_3945_),
    .S(_4075_),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8316_ (.I(_4078_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8317_ (.I(_4072_),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8318_ (.I(_4079_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8319_ (.I(_4075_),
    .Z(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8320_ (.A1(\reg_file.reg_storage[6][4] ),
    .A2(_4081_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8321_ (.A1(_3947_),
    .A2(_4080_),
    .B(_4082_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8322_ (.A1(\reg_file.reg_storage[6][5] ),
    .A2(_4081_),
    .ZN(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8323_ (.A1(_3952_),
    .A2(_4080_),
    .B(_4083_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8324_ (.A1(\reg_file.reg_storage[6][6] ),
    .A2(_4081_),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8325_ (.A1(_3954_),
    .A2(_4080_),
    .B(_4084_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8326_ (.A1(\reg_file.reg_storage[6][7] ),
    .A2(_4081_),
    .ZN(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8327_ (.A1(_3956_),
    .A2(_4080_),
    .B(_4085_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8328_ (.I(_4079_),
    .Z(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8329_ (.I(_4071_),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8330_ (.I(_4087_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8331_ (.A1(\reg_file.reg_storage[6][8] ),
    .A2(_4088_),
    .ZN(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8332_ (.A1(_3958_),
    .A2(_4086_),
    .B(_4089_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8333_ (.A1(\reg_file.reg_storage[6][9] ),
    .A2(_4088_),
    .ZN(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8334_ (.A1(_3963_),
    .A2(_4086_),
    .B(_4090_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8335_ (.A1(\reg_file.reg_storage[6][10] ),
    .A2(_4088_),
    .ZN(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8336_ (.A1(_3965_),
    .A2(_4086_),
    .B(_4091_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8337_ (.A1(\reg_file.reg_storage[6][11] ),
    .A2(_4088_),
    .ZN(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8338_ (.A1(_3967_),
    .A2(_4086_),
    .B(_4092_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8339_ (.I(_4079_),
    .Z(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8340_ (.I(_4087_),
    .Z(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8341_ (.A1(\reg_file.reg_storage[6][12] ),
    .A2(_4094_),
    .ZN(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8342_ (.A1(_3969_),
    .A2(_4093_),
    .B(_4095_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8343_ (.A1(\reg_file.reg_storage[6][13] ),
    .A2(_4094_),
    .ZN(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8344_ (.A1(_3973_),
    .A2(_4093_),
    .B(_4096_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8345_ (.A1(\reg_file.reg_storage[6][14] ),
    .A2(_4094_),
    .ZN(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8346_ (.A1(_3975_),
    .A2(_4093_),
    .B(_4097_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8347_ (.A1(\reg_file.reg_storage[6][15] ),
    .A2(_4094_),
    .ZN(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8348_ (.A1(_3977_),
    .A2(_4093_),
    .B(_4098_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8349_ (.I(_4079_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8350_ (.I(_4087_),
    .Z(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8351_ (.A1(\reg_file.reg_storage[6][16] ),
    .A2(_4100_),
    .ZN(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8352_ (.A1(_3979_),
    .A2(_4099_),
    .B(_4101_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8353_ (.A1(\reg_file.reg_storage[6][17] ),
    .A2(_4100_),
    .ZN(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8354_ (.A1(_3983_),
    .A2(_4099_),
    .B(_4102_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8355_ (.A1(\reg_file.reg_storage[6][18] ),
    .A2(_4100_),
    .ZN(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8356_ (.A1(_3985_),
    .A2(_4099_),
    .B(_4103_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8357_ (.A1(\reg_file.reg_storage[6][19] ),
    .A2(_4100_),
    .ZN(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8358_ (.A1(_3987_),
    .A2(_4099_),
    .B(_4104_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8359_ (.I(_4073_),
    .Z(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8360_ (.I(_4087_),
    .Z(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8361_ (.A1(\reg_file.reg_storage[6][20] ),
    .A2(_4106_),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8362_ (.A1(_3989_),
    .A2(_4105_),
    .B(_4107_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8363_ (.A1(\reg_file.reg_storage[6][21] ),
    .A2(_4106_),
    .ZN(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8364_ (.A1(_3993_),
    .A2(_4105_),
    .B(_4108_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8365_ (.A1(\reg_file.reg_storage[6][22] ),
    .A2(_4106_),
    .ZN(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8366_ (.A1(_3995_),
    .A2(_4105_),
    .B(_4109_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8367_ (.A1(\reg_file.reg_storage[6][23] ),
    .A2(_4106_),
    .ZN(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8368_ (.A1(_3997_),
    .A2(_4105_),
    .B(_4110_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8369_ (.I(_4073_),
    .Z(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8370_ (.I(_4072_),
    .Z(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8371_ (.A1(\reg_file.reg_storage[6][24] ),
    .A2(_4112_),
    .ZN(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8372_ (.A1(_3999_),
    .A2(_4111_),
    .B(_4113_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8373_ (.A1(\reg_file.reg_storage[6][25] ),
    .A2(_4112_),
    .ZN(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8374_ (.A1(_4003_),
    .A2(_4111_),
    .B(_4114_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8375_ (.A1(\reg_file.reg_storage[6][26] ),
    .A2(_4112_),
    .ZN(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8376_ (.A1(_4005_),
    .A2(_4111_),
    .B(_4115_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8377_ (.A1(\reg_file.reg_storage[6][27] ),
    .A2(_4112_),
    .ZN(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8378_ (.A1(_4007_),
    .A2(_4111_),
    .B(_4116_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8379_ (.I(_4073_),
    .Z(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8380_ (.I(_4072_),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8381_ (.A1(\reg_file.reg_storage[6][28] ),
    .A2(_4118_),
    .ZN(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8382_ (.A1(_4009_),
    .A2(_4117_),
    .B(_4119_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8383_ (.A1(\reg_file.reg_storage[6][29] ),
    .A2(_4118_),
    .ZN(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8384_ (.A1(_4013_),
    .A2(_4117_),
    .B(_4120_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8385_ (.A1(\reg_file.reg_storage[6][30] ),
    .A2(_4118_),
    .ZN(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8386_ (.A1(_4015_),
    .A2(_4117_),
    .B(_4121_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8387_ (.A1(\reg_file.reg_storage[6][31] ),
    .A2(_4118_),
    .ZN(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8388_ (.A1(_4017_),
    .A2(_4117_),
    .B(_4122_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8389_ (.A1(_2896_),
    .A2(_0554_),
    .Z(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8390_ (.A1(_2884_),
    .A2(_2897_),
    .A3(_4123_),
    .B1(_3098_),
    .B2(_2896_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8391_ (.A1(_2897_),
    .A2(_2898_),
    .Z(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8392_ (.A1(net76),
    .A2(_3151_),
    .B1(_3183_),
    .B2(_4124_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8393_ (.A1(_0664_),
    .A2(_2887_),
    .B(_4125_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8394_ (.A1(_3258_),
    .A2(_3775_),
    .A3(_3935_),
    .ZN(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8395_ (.I(_4126_),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8396_ (.I(_4127_),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8397_ (.I0(\reg_file.reg_storage[1][0] ),
    .I1(_3934_),
    .S(_4128_),
    .Z(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8398_ (.I(_4129_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8399_ (.I(_4126_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8400_ (.I0(\reg_file.reg_storage[1][1] ),
    .I1(_3940_),
    .S(_4130_),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8401_ (.I(_4131_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8402_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_3943_),
    .S(_4130_),
    .Z(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8403_ (.I(_4132_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8404_ (.I0(\reg_file.reg_storage[1][3] ),
    .I1(_3945_),
    .S(_4130_),
    .Z(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8405_ (.I(_4133_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8406_ (.I(_4127_),
    .Z(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8407_ (.I(_4134_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8408_ (.I(_4130_),
    .Z(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8409_ (.A1(\reg_file.reg_storage[1][4] ),
    .A2(_4136_),
    .ZN(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8410_ (.A1(_3947_),
    .A2(_4135_),
    .B(_4137_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8411_ (.A1(\reg_file.reg_storage[1][5] ),
    .A2(_4136_),
    .ZN(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8412_ (.A1(_3952_),
    .A2(_4135_),
    .B(_4138_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8413_ (.A1(\reg_file.reg_storage[1][6] ),
    .A2(_4136_),
    .ZN(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8414_ (.A1(_3954_),
    .A2(_4135_),
    .B(_4139_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8415_ (.A1(\reg_file.reg_storage[1][7] ),
    .A2(_4136_),
    .ZN(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8416_ (.A1(_3956_),
    .A2(_4135_),
    .B(_4140_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8417_ (.I(_4134_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8418_ (.I(_4126_),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8419_ (.I(_4142_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8420_ (.A1(\reg_file.reg_storage[1][8] ),
    .A2(_4143_),
    .ZN(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8421_ (.A1(_3958_),
    .A2(_4141_),
    .B(_4144_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8422_ (.A1(\reg_file.reg_storage[1][9] ),
    .A2(_4143_),
    .ZN(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8423_ (.A1(_3963_),
    .A2(_4141_),
    .B(_4145_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8424_ (.A1(\reg_file.reg_storage[1][10] ),
    .A2(_4143_),
    .ZN(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8425_ (.A1(_3965_),
    .A2(_4141_),
    .B(_4146_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8426_ (.A1(\reg_file.reg_storage[1][11] ),
    .A2(_4143_),
    .ZN(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8427_ (.A1(_3967_),
    .A2(_4141_),
    .B(_4147_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8428_ (.I(_4134_),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8429_ (.I(_4142_),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8430_ (.A1(\reg_file.reg_storage[1][12] ),
    .A2(_4149_),
    .ZN(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8431_ (.A1(_3969_),
    .A2(_4148_),
    .B(_4150_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8432_ (.A1(\reg_file.reg_storage[1][13] ),
    .A2(_4149_),
    .ZN(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8433_ (.A1(_3973_),
    .A2(_4148_),
    .B(_4151_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8434_ (.A1(\reg_file.reg_storage[1][14] ),
    .A2(_4149_),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8435_ (.A1(_3975_),
    .A2(_4148_),
    .B(_4152_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8436_ (.A1(\reg_file.reg_storage[1][15] ),
    .A2(_4149_),
    .ZN(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8437_ (.A1(_3977_),
    .A2(_4148_),
    .B(_4153_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8438_ (.I(_4134_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8439_ (.I(_4142_),
    .Z(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8440_ (.A1(\reg_file.reg_storage[1][16] ),
    .A2(_4155_),
    .ZN(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8441_ (.A1(_3979_),
    .A2(_4154_),
    .B(_4156_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8442_ (.A1(\reg_file.reg_storage[1][17] ),
    .A2(_4155_),
    .ZN(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8443_ (.A1(_3983_),
    .A2(_4154_),
    .B(_4157_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8444_ (.A1(\reg_file.reg_storage[1][18] ),
    .A2(_4155_),
    .ZN(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8445_ (.A1(_3985_),
    .A2(_4154_),
    .B(_4158_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8446_ (.A1(\reg_file.reg_storage[1][19] ),
    .A2(_4155_),
    .ZN(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8447_ (.A1(_3987_),
    .A2(_4154_),
    .B(_4159_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8448_ (.I(_4128_),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8449_ (.I(_4142_),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8450_ (.A1(\reg_file.reg_storage[1][20] ),
    .A2(_4161_),
    .ZN(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8451_ (.A1(_3989_),
    .A2(_4160_),
    .B(_4162_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8452_ (.A1(\reg_file.reg_storage[1][21] ),
    .A2(_4161_),
    .ZN(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8453_ (.A1(_3993_),
    .A2(_4160_),
    .B(_4163_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8454_ (.A1(\reg_file.reg_storage[1][22] ),
    .A2(_4161_),
    .ZN(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8455_ (.A1(_3995_),
    .A2(_4160_),
    .B(_4164_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8456_ (.A1(\reg_file.reg_storage[1][23] ),
    .A2(_4161_),
    .ZN(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8457_ (.A1(_3997_),
    .A2(_4160_),
    .B(_4165_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8458_ (.I(_4128_),
    .Z(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8459_ (.I(_4127_),
    .Z(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8460_ (.A1(\reg_file.reg_storage[1][24] ),
    .A2(_4167_),
    .ZN(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8461_ (.A1(_3999_),
    .A2(_4166_),
    .B(_4168_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8462_ (.A1(\reg_file.reg_storage[1][25] ),
    .A2(_4167_),
    .ZN(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8463_ (.A1(_4003_),
    .A2(_4166_),
    .B(_4169_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8464_ (.A1(\reg_file.reg_storage[1][26] ),
    .A2(_4167_),
    .ZN(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8465_ (.A1(_4005_),
    .A2(_4166_),
    .B(_4170_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8466_ (.A1(\reg_file.reg_storage[1][27] ),
    .A2(_4167_),
    .ZN(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8467_ (.A1(_4007_),
    .A2(_4166_),
    .B(_4171_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8468_ (.I(_4128_),
    .Z(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8469_ (.I(_4127_),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8470_ (.A1(\reg_file.reg_storage[1][28] ),
    .A2(_4173_),
    .ZN(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8471_ (.A1(_4009_),
    .A2(_4172_),
    .B(_4174_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8472_ (.A1(\reg_file.reg_storage[1][29] ),
    .A2(_4173_),
    .ZN(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8473_ (.A1(_4013_),
    .A2(_4172_),
    .B(_4175_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8474_ (.A1(\reg_file.reg_storage[1][30] ),
    .A2(_4173_),
    .ZN(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8475_ (.A1(_4015_),
    .A2(_4172_),
    .B(_4176_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8476_ (.A1(\reg_file.reg_storage[1][31] ),
    .A2(_4173_),
    .ZN(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8477_ (.A1(_4017_),
    .A2(_4172_),
    .B(_4177_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8478_ (.A1(_3258_),
    .A2(_3775_),
    .A3(_3774_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8479_ (.I(_4178_),
    .Z(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8480_ (.I(_4179_),
    .Z(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8481_ (.I0(\reg_file.reg_storage[3][0] ),
    .I1(_3253_),
    .S(_4180_),
    .Z(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8482_ (.I(_4181_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8483_ (.I(_4178_),
    .Z(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8484_ (.I0(\reg_file.reg_storage[3][1] ),
    .I1(_3274_),
    .S(_4182_),
    .Z(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8485_ (.I(_4183_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8486_ (.I0(\reg_file.reg_storage[3][2] ),
    .I1(_3286_),
    .S(_4182_),
    .Z(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8487_ (.I(_4184_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8488_ (.I0(\reg_file.reg_storage[3][3] ),
    .I1(_3295_),
    .S(_4182_),
    .Z(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8489_ (.I(_4185_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8490_ (.I(_4179_),
    .Z(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8491_ (.I(_4186_),
    .Z(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8492_ (.I(_4182_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8493_ (.A1(\reg_file.reg_storage[3][4] ),
    .A2(_4188_),
    .ZN(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8494_ (.A1(_3674_),
    .A2(_4187_),
    .B(_4189_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8495_ (.A1(\reg_file.reg_storage[3][5] ),
    .A2(_4188_),
    .ZN(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8496_ (.A1(_3680_),
    .A2(_4187_),
    .B(_4190_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8497_ (.A1(\reg_file.reg_storage[3][6] ),
    .A2(_4188_),
    .ZN(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8498_ (.A1(_3683_),
    .A2(_4187_),
    .B(_4191_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8499_ (.A1(\reg_file.reg_storage[3][7] ),
    .A2(_4188_),
    .ZN(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8500_ (.A1(_3686_),
    .A2(_4187_),
    .B(_4192_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8501_ (.I(_4186_),
    .Z(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8502_ (.I(_4178_),
    .Z(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8503_ (.I(_4194_),
    .Z(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8504_ (.A1(\reg_file.reg_storage[3][8] ),
    .A2(_4195_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8505_ (.A1(_3689_),
    .A2(_4193_),
    .B(_4196_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8506_ (.A1(\reg_file.reg_storage[3][9] ),
    .A2(_4195_),
    .ZN(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8507_ (.A1(_3695_),
    .A2(_4193_),
    .B(_4197_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8508_ (.A1(\reg_file.reg_storage[3][10] ),
    .A2(_4195_),
    .ZN(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8509_ (.A1(_3698_),
    .A2(_4193_),
    .B(_4198_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8510_ (.A1(\reg_file.reg_storage[3][11] ),
    .A2(_4195_),
    .ZN(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8511_ (.A1(_3701_),
    .A2(_4193_),
    .B(_4199_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8512_ (.I(_4186_),
    .Z(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8513_ (.I(_4194_),
    .Z(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8514_ (.A1(\reg_file.reg_storage[3][12] ),
    .A2(_4201_),
    .ZN(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8515_ (.A1(_3704_),
    .A2(_4200_),
    .B(_4202_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8516_ (.A1(\reg_file.reg_storage[3][13] ),
    .A2(_4201_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8517_ (.A1(_3709_),
    .A2(_4200_),
    .B(_4203_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8518_ (.A1(\reg_file.reg_storage[3][14] ),
    .A2(_4201_),
    .ZN(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8519_ (.A1(_3712_),
    .A2(_4200_),
    .B(_4204_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8520_ (.A1(\reg_file.reg_storage[3][15] ),
    .A2(_4201_),
    .ZN(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8521_ (.A1(_3715_),
    .A2(_4200_),
    .B(_4205_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8522_ (.I(_4186_),
    .Z(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8523_ (.I(_4194_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8524_ (.A1(\reg_file.reg_storage[3][16] ),
    .A2(_4207_),
    .ZN(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8525_ (.A1(_3718_),
    .A2(_4206_),
    .B(_4208_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8526_ (.A1(\reg_file.reg_storage[3][17] ),
    .A2(_4207_),
    .ZN(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8527_ (.A1(_3723_),
    .A2(_4206_),
    .B(_4209_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8528_ (.A1(\reg_file.reg_storage[3][18] ),
    .A2(_4207_),
    .ZN(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8529_ (.A1(_3726_),
    .A2(_4206_),
    .B(_4210_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8530_ (.A1(\reg_file.reg_storage[3][19] ),
    .A2(_4207_),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8531_ (.A1(_3729_),
    .A2(_4206_),
    .B(_4211_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8532_ (.I(_4180_),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8533_ (.I(_4194_),
    .Z(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8534_ (.A1(\reg_file.reg_storage[3][20] ),
    .A2(_4213_),
    .ZN(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8535_ (.A1(_3732_),
    .A2(_4212_),
    .B(_4214_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8536_ (.A1(\reg_file.reg_storage[3][21] ),
    .A2(_4213_),
    .ZN(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8537_ (.A1(_3737_),
    .A2(_4212_),
    .B(_4215_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8538_ (.A1(\reg_file.reg_storage[3][22] ),
    .A2(_4213_),
    .ZN(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8539_ (.A1(_3740_),
    .A2(_4212_),
    .B(_4216_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8540_ (.A1(\reg_file.reg_storage[3][23] ),
    .A2(_4213_),
    .ZN(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8541_ (.A1(_3743_),
    .A2(_4212_),
    .B(_4217_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8542_ (.I(_4180_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8543_ (.I(_4179_),
    .Z(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8544_ (.A1(\reg_file.reg_storage[3][24] ),
    .A2(_4219_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8545_ (.A1(_3746_),
    .A2(_4218_),
    .B(_4220_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8546_ (.A1(\reg_file.reg_storage[3][25] ),
    .A2(_4219_),
    .ZN(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8547_ (.A1(_3751_),
    .A2(_4218_),
    .B(_4221_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8548_ (.A1(\reg_file.reg_storage[3][26] ),
    .A2(_4219_),
    .ZN(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8549_ (.A1(_3754_),
    .A2(_4218_),
    .B(_4222_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8550_ (.A1(\reg_file.reg_storage[3][27] ),
    .A2(_4219_),
    .ZN(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8551_ (.A1(_3757_),
    .A2(_4218_),
    .B(_4223_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8552_ (.I(_4180_),
    .Z(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8553_ (.I(_4179_),
    .Z(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8554_ (.A1(\reg_file.reg_storage[3][28] ),
    .A2(_4225_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8555_ (.A1(_3760_),
    .A2(_4224_),
    .B(_4226_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8556_ (.A1(\reg_file.reg_storage[3][29] ),
    .A2(_4225_),
    .ZN(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8557_ (.A1(_3765_),
    .A2(_4224_),
    .B(_4227_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8558_ (.A1(\reg_file.reg_storage[3][30] ),
    .A2(_4225_),
    .ZN(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8559_ (.A1(_3768_),
    .A2(_4224_),
    .B(_4228_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8560_ (.A1(\reg_file.reg_storage[3][31] ),
    .A2(_4225_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8561_ (.A1(_3771_),
    .A2(_4224_),
    .B(_4229_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8562_ (.A1(_3607_),
    .A2(_3553_),
    .A3(_3264_),
    .ZN(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8563_ (.I(_4230_),
    .Z(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8564_ (.I(_4231_),
    .Z(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8565_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(_3253_),
    .S(_4232_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8566_ (.I(_4233_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8567_ (.I(_4230_),
    .Z(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8568_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(_3274_),
    .S(_4234_),
    .Z(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8569_ (.I(_4235_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8570_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(_3286_),
    .S(_4234_),
    .Z(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8571_ (.I(_4236_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8572_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(_3295_),
    .S(_4234_),
    .Z(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8573_ (.I(_4237_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8574_ (.I(_4231_),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8575_ (.I(_4238_),
    .Z(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8576_ (.I(_4234_),
    .Z(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8577_ (.A1(\reg_file.reg_storage[8][4] ),
    .A2(_4240_),
    .ZN(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8578_ (.A1(_3674_),
    .A2(_4239_),
    .B(_4241_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8579_ (.A1(\reg_file.reg_storage[8][5] ),
    .A2(_4240_),
    .ZN(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8580_ (.A1(_3680_),
    .A2(_4239_),
    .B(_4242_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8581_ (.A1(\reg_file.reg_storage[8][6] ),
    .A2(_4240_),
    .ZN(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8582_ (.A1(_3683_),
    .A2(_4239_),
    .B(_4243_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8583_ (.A1(\reg_file.reg_storage[8][7] ),
    .A2(_4240_),
    .ZN(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8584_ (.A1(_3686_),
    .A2(_4239_),
    .B(_4244_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8585_ (.I(_4238_),
    .Z(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8586_ (.I(_4230_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8587_ (.I(_4246_),
    .Z(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8588_ (.A1(\reg_file.reg_storage[8][8] ),
    .A2(_4247_),
    .ZN(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8589_ (.A1(_3689_),
    .A2(_4245_),
    .B(_4248_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8590_ (.A1(\reg_file.reg_storage[8][9] ),
    .A2(_4247_),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8591_ (.A1(_3695_),
    .A2(_4245_),
    .B(_4249_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8592_ (.A1(\reg_file.reg_storage[8][10] ),
    .A2(_4247_),
    .ZN(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8593_ (.A1(_3698_),
    .A2(_4245_),
    .B(_4250_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8594_ (.A1(\reg_file.reg_storage[8][11] ),
    .A2(_4247_),
    .ZN(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8595_ (.A1(_3701_),
    .A2(_4245_),
    .B(_4251_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8596_ (.I(_4238_),
    .Z(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8597_ (.I(_4246_),
    .Z(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8598_ (.A1(\reg_file.reg_storage[8][12] ),
    .A2(_4253_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8599_ (.A1(_3704_),
    .A2(_4252_),
    .B(_4254_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8600_ (.A1(\reg_file.reg_storage[8][13] ),
    .A2(_4253_),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8601_ (.A1(_3709_),
    .A2(_4252_),
    .B(_4255_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8602_ (.A1(\reg_file.reg_storage[8][14] ),
    .A2(_4253_),
    .ZN(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8603_ (.A1(_3712_),
    .A2(_4252_),
    .B(_4256_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8604_ (.A1(\reg_file.reg_storage[8][15] ),
    .A2(_4253_),
    .ZN(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8605_ (.A1(_3715_),
    .A2(_4252_),
    .B(_4257_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8606_ (.I(_4238_),
    .Z(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8607_ (.I(_4246_),
    .Z(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8608_ (.A1(\reg_file.reg_storage[8][16] ),
    .A2(_4259_),
    .ZN(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8609_ (.A1(_3718_),
    .A2(_4258_),
    .B(_4260_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8610_ (.A1(\reg_file.reg_storage[8][17] ),
    .A2(_4259_),
    .ZN(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8611_ (.A1(_3723_),
    .A2(_4258_),
    .B(_4261_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8612_ (.A1(\reg_file.reg_storage[8][18] ),
    .A2(_4259_),
    .ZN(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8613_ (.A1(_3726_),
    .A2(_4258_),
    .B(_4262_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8614_ (.A1(\reg_file.reg_storage[8][19] ),
    .A2(_4259_),
    .ZN(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8615_ (.A1(_3729_),
    .A2(_4258_),
    .B(_4263_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8616_ (.I(_4232_),
    .Z(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8617_ (.I(_4246_),
    .Z(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8618_ (.A1(\reg_file.reg_storage[8][20] ),
    .A2(_4265_),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8619_ (.A1(_3732_),
    .A2(_4264_),
    .B(_4266_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8620_ (.A1(\reg_file.reg_storage[8][21] ),
    .A2(_4265_),
    .ZN(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8621_ (.A1(_3737_),
    .A2(_4264_),
    .B(_4267_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8622_ (.A1(\reg_file.reg_storage[8][22] ),
    .A2(_4265_),
    .ZN(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8623_ (.A1(_3740_),
    .A2(_4264_),
    .B(_4268_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8624_ (.A1(\reg_file.reg_storage[8][23] ),
    .A2(_4265_),
    .ZN(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8625_ (.A1(_3743_),
    .A2(_4264_),
    .B(_4269_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8626_ (.I(_4232_),
    .Z(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8627_ (.I(_4231_),
    .Z(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8628_ (.A1(\reg_file.reg_storage[8][24] ),
    .A2(_4271_),
    .ZN(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8629_ (.A1(_3746_),
    .A2(_4270_),
    .B(_4272_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8630_ (.A1(\reg_file.reg_storage[8][25] ),
    .A2(_4271_),
    .ZN(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8631_ (.A1(_3751_),
    .A2(_4270_),
    .B(_4273_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8632_ (.A1(\reg_file.reg_storage[8][26] ),
    .A2(_4271_),
    .ZN(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8633_ (.A1(_3754_),
    .A2(_4270_),
    .B(_4274_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8634_ (.A1(\reg_file.reg_storage[8][27] ),
    .A2(_4271_),
    .ZN(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8635_ (.A1(_3757_),
    .A2(_4270_),
    .B(_4275_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8636_ (.I(_4232_),
    .Z(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8637_ (.I(_4231_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8638_ (.A1(\reg_file.reg_storage[8][28] ),
    .A2(_4277_),
    .ZN(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8639_ (.A1(_3760_),
    .A2(_4276_),
    .B(_4278_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8640_ (.A1(\reg_file.reg_storage[8][29] ),
    .A2(_4277_),
    .ZN(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8641_ (.A1(_3765_),
    .A2(_4276_),
    .B(_4279_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8642_ (.A1(\reg_file.reg_storage[8][30] ),
    .A2(_4277_),
    .ZN(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8643_ (.A1(_3768_),
    .A2(_4276_),
    .B(_4280_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8644_ (.A1(\reg_file.reg_storage[8][31] ),
    .A2(_4277_),
    .ZN(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8645_ (.A1(_3771_),
    .A2(_4276_),
    .B(_4281_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8646_ (.A1(_3499_),
    .A2(_3554_),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8647_ (.I(_4282_),
    .Z(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8648_ (.I(_4283_),
    .Z(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8649_ (.I0(\reg_file.reg_storage[5][0] ),
    .I1(_3253_),
    .S(_4284_),
    .Z(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8650_ (.I(_4285_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8651_ (.I(_4282_),
    .Z(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8652_ (.I0(\reg_file.reg_storage[5][1] ),
    .I1(_3274_),
    .S(_4286_),
    .Z(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8653_ (.I(_4287_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8654_ (.I0(\reg_file.reg_storage[5][2] ),
    .I1(_3286_),
    .S(_4286_),
    .Z(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8655_ (.I(_4288_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8656_ (.I0(\reg_file.reg_storage[5][3] ),
    .I1(_3295_),
    .S(_4286_),
    .Z(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8657_ (.I(_4289_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8658_ (.I(_4283_),
    .Z(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8659_ (.I(_4290_),
    .Z(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8660_ (.I(_4286_),
    .Z(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8661_ (.A1(\reg_file.reg_storage[5][4] ),
    .A2(_4292_),
    .ZN(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8662_ (.A1(_3674_),
    .A2(_4291_),
    .B(_4293_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8663_ (.A1(\reg_file.reg_storage[5][5] ),
    .A2(_4292_),
    .ZN(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8664_ (.A1(_3680_),
    .A2(_4291_),
    .B(_4294_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8665_ (.A1(\reg_file.reg_storage[5][6] ),
    .A2(_4292_),
    .ZN(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8666_ (.A1(_3683_),
    .A2(_4291_),
    .B(_4295_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8667_ (.A1(\reg_file.reg_storage[5][7] ),
    .A2(_4292_),
    .ZN(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8668_ (.A1(_3686_),
    .A2(_4291_),
    .B(_4296_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8669_ (.I(_4290_),
    .Z(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8670_ (.I(_4282_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8671_ (.I(_4298_),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8672_ (.A1(\reg_file.reg_storage[5][8] ),
    .A2(_4299_),
    .ZN(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8673_ (.A1(_3689_),
    .A2(_4297_),
    .B(_4300_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8674_ (.A1(\reg_file.reg_storage[5][9] ),
    .A2(_4299_),
    .ZN(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8675_ (.A1(_3695_),
    .A2(_4297_),
    .B(_4301_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8676_ (.A1(\reg_file.reg_storage[5][10] ),
    .A2(_4299_),
    .ZN(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8677_ (.A1(_3698_),
    .A2(_4297_),
    .B(_4302_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8678_ (.A1(\reg_file.reg_storage[5][11] ),
    .A2(_4299_),
    .ZN(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8679_ (.A1(_3701_),
    .A2(_4297_),
    .B(_4303_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8680_ (.I(_4290_),
    .Z(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8681_ (.I(_4298_),
    .Z(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8682_ (.A1(\reg_file.reg_storage[5][12] ),
    .A2(_4305_),
    .ZN(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8683_ (.A1(_3704_),
    .A2(_4304_),
    .B(_4306_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8684_ (.A1(\reg_file.reg_storage[5][13] ),
    .A2(_4305_),
    .ZN(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8685_ (.A1(_3709_),
    .A2(_4304_),
    .B(_4307_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8686_ (.A1(\reg_file.reg_storage[5][14] ),
    .A2(_4305_),
    .ZN(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8687_ (.A1(_3712_),
    .A2(_4304_),
    .B(_4308_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8688_ (.A1(\reg_file.reg_storage[5][15] ),
    .A2(_4305_),
    .ZN(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8689_ (.A1(_3715_),
    .A2(_4304_),
    .B(_4309_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8690_ (.I(_4290_),
    .Z(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8691_ (.I(_4298_),
    .Z(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8692_ (.A1(\reg_file.reg_storage[5][16] ),
    .A2(_4311_),
    .ZN(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8693_ (.A1(_3718_),
    .A2(_4310_),
    .B(_4312_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8694_ (.A1(\reg_file.reg_storage[5][17] ),
    .A2(_4311_),
    .ZN(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8695_ (.A1(_3723_),
    .A2(_4310_),
    .B(_4313_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8696_ (.A1(\reg_file.reg_storage[5][18] ),
    .A2(_4311_),
    .ZN(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8697_ (.A1(_3726_),
    .A2(_4310_),
    .B(_4314_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8698_ (.A1(\reg_file.reg_storage[5][19] ),
    .A2(_4311_),
    .ZN(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8699_ (.A1(_3729_),
    .A2(_4310_),
    .B(_4315_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8700_ (.I(_4284_),
    .Z(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8701_ (.I(_4298_),
    .Z(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8702_ (.A1(\reg_file.reg_storage[5][20] ),
    .A2(_4317_),
    .ZN(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8703_ (.A1(_3732_),
    .A2(_4316_),
    .B(_4318_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8704_ (.A1(\reg_file.reg_storage[5][21] ),
    .A2(_4317_),
    .ZN(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8705_ (.A1(_3737_),
    .A2(_4316_),
    .B(_4319_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8706_ (.A1(\reg_file.reg_storage[5][22] ),
    .A2(_4317_),
    .ZN(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8707_ (.A1(_3740_),
    .A2(_4316_),
    .B(_4320_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8708_ (.A1(\reg_file.reg_storage[5][23] ),
    .A2(_4317_),
    .ZN(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8709_ (.A1(_3743_),
    .A2(_4316_),
    .B(_4321_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8710_ (.I(_4284_),
    .Z(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8711_ (.I(_4283_),
    .Z(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8712_ (.A1(\reg_file.reg_storage[5][24] ),
    .A2(_4323_),
    .ZN(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8713_ (.A1(_3746_),
    .A2(_4322_),
    .B(_4324_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8714_ (.A1(\reg_file.reg_storage[5][25] ),
    .A2(_4323_),
    .ZN(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8715_ (.A1(_3751_),
    .A2(_4322_),
    .B(_4325_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8716_ (.A1(\reg_file.reg_storage[5][26] ),
    .A2(_4323_),
    .ZN(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8717_ (.A1(_3754_),
    .A2(_4322_),
    .B(_4326_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8718_ (.A1(\reg_file.reg_storage[5][27] ),
    .A2(_4323_),
    .ZN(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8719_ (.A1(_3757_),
    .A2(_4322_),
    .B(_4327_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8720_ (.I(_4284_),
    .Z(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8721_ (.I(_4283_),
    .Z(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8722_ (.A1(\reg_file.reg_storage[5][28] ),
    .A2(_4329_),
    .ZN(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8723_ (.A1(_3760_),
    .A2(_4328_),
    .B(_4330_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8724_ (.A1(\reg_file.reg_storage[5][29] ),
    .A2(_4329_),
    .ZN(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8725_ (.A1(_3765_),
    .A2(_4328_),
    .B(_4331_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8726_ (.A1(\reg_file.reg_storage[5][30] ),
    .A2(_4329_),
    .ZN(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8727_ (.A1(_3768_),
    .A2(_4328_),
    .B(_4332_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8728_ (.A1(\reg_file.reg_storage[5][31] ),
    .A2(_4329_),
    .ZN(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8729_ (.A1(_3771_),
    .A2(_4328_),
    .B(_4333_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8730_ (.D(_0000_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8731_ (.D(_0001_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8732_ (.D(_0002_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8733_ (.D(_0003_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8734_ (.D(_0004_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8735_ (.D(_0005_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8736_ (.D(_0006_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8737_ (.D(_0007_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8738_ (.D(_0008_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8739_ (.D(_0009_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8740_ (.D(_0010_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8741_ (.D(_0011_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8742_ (.D(_0012_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8743_ (.D(_0013_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8744_ (.D(_0014_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8745_ (.D(_0015_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8746_ (.D(_0016_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[11][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8747_ (.D(_0017_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8748_ (.D(_0018_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8749_ (.D(_0019_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[11][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8750_ (.D(_0020_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8751_ (.D(_0021_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[11][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8752_ (.D(_0022_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8753_ (.D(_0023_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8754_ (.D(_0024_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8755_ (.D(_0025_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8756_ (.D(_0026_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[11][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8757_ (.D(_0027_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8758_ (.D(_0028_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8759_ (.D(_0029_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[11][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8760_ (.D(_0030_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8761_ (.D(_0031_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8762_ (.D(_0032_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8763_ (.D(_0033_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8764_ (.D(_0034_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8765_ (.D(_0035_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8766_ (.D(_0036_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8767_ (.D(_0037_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8768_ (.D(_0038_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8769_ (.D(_0039_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8770_ (.D(_0040_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8771_ (.D(_0041_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8772_ (.D(_0042_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8773_ (.D(_0043_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8774_ (.D(_0044_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8775_ (.D(_0045_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8776_ (.D(_0046_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8777_ (.D(_0047_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8778_ (.D(_0048_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8779_ (.D(_0049_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8780_ (.D(_0050_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8781_ (.D(_0051_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[7][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8782_ (.D(_0052_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8783_ (.D(_0053_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8784_ (.D(_0054_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8785_ (.D(_0055_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8786_ (.D(_0056_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8787_ (.D(_0057_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8788_ (.D(_0058_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8789_ (.D(_0059_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8790_ (.D(_0060_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8791_ (.D(_0061_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8792_ (.D(_0062_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8793_ (.D(_0063_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8794_ (.D(_0064_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8795_ (.D(_0065_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8796_ (.D(_0066_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8797_ (.D(_0067_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8798_ (.D(_0068_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8799_ (.D(_0069_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8800_ (.D(_0070_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8801_ (.D(_0071_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8802_ (.D(_0072_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8803_ (.D(_0073_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8804_ (.D(_0074_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8805_ (.D(_0075_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8806_ (.D(_0076_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8807_ (.D(_0077_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8808_ (.D(_0078_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8809_ (.D(_0079_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8810_ (.D(_0080_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[9][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8811_ (.D(_0081_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8812_ (.D(_0082_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8813_ (.D(_0083_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8814_ (.D(_0084_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8815_ (.D(_0085_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8816_ (.D(_0086_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8817_ (.D(_0087_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8818_ (.D(_0088_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8819_ (.D(_0089_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8820_ (.D(_0090_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8821_ (.D(_0091_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8822_ (.D(_0092_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[9][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8823_ (.D(_0093_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8824_ (.D(_0094_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8825_ (.D(_0095_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8826_ (.D(_0096_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8827_ (.D(_0097_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8828_ (.D(_0098_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8829_ (.D(_0099_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8830_ (.D(_0100_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8831_ (.D(_0101_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8832_ (.D(_0102_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8833_ (.D(_0103_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8834_ (.D(_0104_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8835_ (.D(_0105_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8836_ (.D(_0106_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8837_ (.D(_0107_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8838_ (.D(_0108_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8839_ (.D(_0109_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8840_ (.D(_0110_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8841_ (.D(_0111_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8842_ (.D(_0112_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[10][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8843_ (.D(_0113_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8844_ (.D(_0114_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8845_ (.D(_0115_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8846_ (.D(_0116_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[10][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8847_ (.D(_0117_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[10][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8848_ (.D(_0118_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[10][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8849_ (.D(_0119_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[10][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8850_ (.D(_0120_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8851_ (.D(_0121_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[10][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8852_ (.D(_0122_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[10][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8853_ (.D(_0123_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8854_ (.D(_0124_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[10][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8855_ (.D(_0125_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[10][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8856_ (.D(_0126_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8857_ (.D(_0127_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8858_ (.D(_0128_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8859_ (.D(_0129_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8860_ (.D(_0130_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8861_ (.D(_0131_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8862_ (.D(_0132_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8863_ (.D(_0133_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8864_ (.D(_0134_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8865_ (.D(_0135_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8866_ (.D(_0136_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8867_ (.D(_0137_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8868_ (.D(_0138_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8869_ (.D(_0139_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8870_ (.D(_0140_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8871_ (.D(_0141_),
    .CLK(clknet_leaf_63_clk),
    .Q(\reg_file.reg_storage[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8872_ (.D(_0142_),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\reg_file.reg_storage[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8873_ (.D(_0143_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8874_ (.D(_0144_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8875_ (.D(_0145_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8876_ (.D(_0146_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8877_ (.D(_0147_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8878_ (.D(_0148_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[4][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8879_ (.D(_0149_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8880_ (.D(_0150_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[4][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8881_ (.D(_0151_),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\reg_file.reg_storage[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8882_ (.D(_0152_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8883_ (.D(_0153_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8884_ (.D(_0154_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8885_ (.D(_0155_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[4][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8886_ (.D(_0156_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8887_ (.D(_0157_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[4][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8888_ (.D(_0158_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[4][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8889_ (.D(_0159_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[4][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8890_ (.D(_0160_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8891_ (.D(_0161_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8892_ (.D(_0162_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8893_ (.D(_0163_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8894_ (.D(_0164_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8895_ (.D(_0165_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8896_ (.D(_0166_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8897_ (.D(_0167_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8898_ (.D(_0168_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8899_ (.D(_0169_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8900_ (.D(_0170_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8901_ (.D(_0171_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8902_ (.D(_0172_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8903_ (.D(_0173_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8904_ (.D(_0174_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8905_ (.D(_0175_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8906_ (.D(_0176_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[15][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8907_ (.D(_0177_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8908_ (.D(_0178_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[15][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8909_ (.D(_0179_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[15][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8910_ (.D(_0180_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8911_ (.D(_0181_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8912_ (.D(_0182_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8913_ (.D(_0183_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8914_ (.D(_0184_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8915_ (.D(_0185_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8916_ (.D(_0186_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8917_ (.D(_0187_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8918_ (.D(_0188_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8919_ (.D(_0189_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8920_ (.D(_0190_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[15][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8921_ (.D(_0191_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8922_ (.D(_0192_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8923_ (.D(_0193_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8924_ (.D(_0194_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8925_ (.D(_0195_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8926_ (.D(_0196_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8927_ (.D(_0197_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8928_ (.D(_0198_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8929_ (.D(_0199_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8930_ (.D(_0200_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8931_ (.D(_0201_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8932_ (.D(_0202_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8933_ (.D(_0203_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8934_ (.D(_0204_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8935_ (.D(_0205_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8936_ (.D(_0206_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8937_ (.D(_0207_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8938_ (.D(_0208_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8939_ (.D(_0209_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8940_ (.D(_0210_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8941_ (.D(_0211_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8942_ (.D(_0212_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8943_ (.D(_0213_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8944_ (.D(_0214_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8945_ (.D(_0215_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8946_ (.D(_0216_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8947_ (.D(_0217_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8948_ (.D(_0218_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8949_ (.D(_0219_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8950_ (.D(_0220_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[2][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8951_ (.D(_0221_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[2][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8952_ (.D(_0222_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8953_ (.D(_0223_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[2][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8954_ (.D(_0224_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8955_ (.D(_0225_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8956_ (.D(_0226_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8957_ (.D(_0227_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8958_ (.D(_0228_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8959_ (.D(_0229_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8960_ (.D(_0230_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8961_ (.D(_0231_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8962_ (.D(_0232_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8963_ (.D(_0233_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8964_ (.D(_0234_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8965_ (.D(_0235_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8966_ (.D(_0236_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8967_ (.D(_0237_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8968_ (.D(_0238_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8969_ (.D(_0239_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8970_ (.D(_0240_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[12][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8971_ (.D(_0241_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8972_ (.D(_0242_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[12][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8973_ (.D(_0243_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[12][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8974_ (.D(_0244_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[12][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8975_ (.D(_0245_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[12][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8976_ (.D(_0246_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8977_ (.D(_0247_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8978_ (.D(_0248_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[12][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8979_ (.D(_0249_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8980_ (.D(_0250_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[12][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8981_ (.D(_0251_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8982_ (.D(_0252_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8983_ (.D(_0253_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[12][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8984_ (.D(_0254_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[12][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8985_ (.D(_0255_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[12][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8986_ (.D(_0256_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8987_ (.D(_0257_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8988_ (.D(_0258_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8989_ (.D(_0259_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8990_ (.D(_0260_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8991_ (.D(_0261_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8992_ (.D(_0262_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8993_ (.D(_0263_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8994_ (.D(_0264_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8995_ (.D(_0265_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8996_ (.D(_0266_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8997_ (.D(_0267_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8998_ (.D(_0268_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8999_ (.D(_0269_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9000_ (.D(_0270_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9001_ (.D(_0271_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9002_ (.D(_0272_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9003_ (.D(_0273_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9004_ (.D(_0274_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9005_ (.D(_0275_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9006_ (.D(_0276_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9007_ (.D(_0277_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9008_ (.D(_0278_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9009_ (.D(_0279_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9010_ (.D(_0280_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9011_ (.D(_0281_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9012_ (.D(_0282_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9013_ (.D(_0283_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9014_ (.D(_0284_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9015_ (.D(_0285_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[13][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9016_ (.D(_0286_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9017_ (.D(_0287_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9018_ (.D(_0288_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9019_ (.D(_0289_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9020_ (.D(_0290_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9021_ (.D(_0291_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9022_ (.D(_0292_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9023_ (.D(_0293_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9024_ (.D(_0294_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9025_ (.D(_0295_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9026_ (.D(_0296_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9027_ (.D(_0297_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9028_ (.D(_0298_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9029_ (.D(_0299_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9030_ (.D(_0300_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9031_ (.D(_0301_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9032_ (.D(_0302_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9033_ (.D(_0303_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9034_ (.D(_0304_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[14][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9035_ (.D(_0305_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9036_ (.D(_0306_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9037_ (.D(_0307_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9038_ (.D(_0308_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9039_ (.D(_0309_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9040_ (.D(_0310_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9041_ (.D(_0311_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9042_ (.D(_0312_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9043_ (.D(_0313_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9044_ (.D(_0314_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9045_ (.D(_0315_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9046_ (.D(_0316_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9047_ (.D(_0317_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9048_ (.D(_0318_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9049_ (.D(_0319_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9050_ (.D(_0320_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9051_ (.D(_0321_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9052_ (.D(_0322_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9053_ (.D(_0323_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9054_ (.D(_0324_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9055_ (.D(_0325_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9056_ (.D(_0326_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9057_ (.D(_0327_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9058_ (.D(_0328_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9059_ (.D(_0329_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9060_ (.D(_0330_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9061_ (.D(_0331_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9062_ (.D(_0332_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9063_ (.D(_0333_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9064_ (.D(_0334_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9065_ (.D(_0335_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9066_ (.D(_0336_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[6][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9067_ (.D(_0337_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[6][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9068_ (.D(_0338_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9069_ (.D(_0339_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[6][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9070_ (.D(_0340_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9071_ (.D(_0341_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9072_ (.D(_0342_),
    .CLK(clknet_leaf_109_clk),
    .Q(\reg_file.reg_storage[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9073_ (.D(_0343_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9074_ (.D(_0344_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9075_ (.D(_0345_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9076_ (.D(_0346_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9077_ (.D(_0347_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9078_ (.D(_0348_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9079_ (.D(_0349_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9080_ (.D(_0350_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9081_ (.D(_0351_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9082_ (.D(_0352_),
    .CLK(clknet_leaf_65_clk),
    .Q(\pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9083_ (.D(_0353_),
    .CLK(clknet_leaf_66_clk),
    .Q(\pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9084_ (.D(_0354_),
    .CLK(clknet_leaf_108_clk),
    .Q(\reg_file.reg_storage[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9085_ (.D(_0355_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9086_ (.D(_0356_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9087_ (.D(_0357_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9088_ (.D(_0358_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9089_ (.D(_0359_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9090_ (.D(_0360_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9091_ (.D(_0361_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9092_ (.D(_0362_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9093_ (.D(_0363_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9094_ (.D(_0364_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9095_ (.D(_0365_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9096_ (.D(_0366_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9097_ (.D(_0367_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9098_ (.D(_0368_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9099_ (.D(_0369_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9100_ (.D(_0370_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9101_ (.D(_0371_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9102_ (.D(_0372_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9103_ (.D(_0373_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9104_ (.D(_0374_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9105_ (.D(_0375_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9106_ (.D(_0376_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9107_ (.D(_0377_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9108_ (.D(_0378_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9109_ (.D(_0379_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9110_ (.D(_0380_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9111_ (.D(_0381_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9112_ (.D(_0382_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[1][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9113_ (.D(_0383_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[1][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9114_ (.D(_0384_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9115_ (.D(_0385_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[1][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9116_ (.D(_0386_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9117_ (.D(_0387_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9118_ (.D(_0388_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9119_ (.D(_0389_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9120_ (.D(_0390_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9121_ (.D(_0391_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9122_ (.D(_0392_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9123_ (.D(_0393_),
    .CLK(clknet_leaf_24_clk),
    .Q(\reg_file.reg_storage[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9124_ (.D(_0394_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9125_ (.D(_0395_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9126_ (.D(_0396_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9127_ (.D(_0397_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9128_ (.D(_0398_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9129_ (.D(_0399_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9130_ (.D(_0400_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9131_ (.D(_0401_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9132_ (.D(_0402_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9133_ (.D(_0403_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9134_ (.D(_0404_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9135_ (.D(_0405_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9136_ (.D(_0406_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9137_ (.D(_0407_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9138_ (.D(_0408_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9139_ (.D(_0409_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9140_ (.D(_0410_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[3][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9141_ (.D(_0411_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[3][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9142_ (.D(_0412_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[3][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9143_ (.D(_0413_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[3][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9144_ (.D(_0414_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9145_ (.D(_0415_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9146_ (.D(_0416_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9147_ (.D(_0417_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9148_ (.D(_0418_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9149_ (.D(_0419_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9150_ (.D(_0420_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9151_ (.D(_0421_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9152_ (.D(_0422_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9153_ (.D(_0423_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9154_ (.D(_0424_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9155_ (.D(_0425_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9156_ (.D(_0426_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9157_ (.D(_0427_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9158_ (.D(_0428_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9159_ (.D(_0429_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9160_ (.D(_0430_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9161_ (.D(_0431_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9162_ (.D(_0432_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9163_ (.D(_0433_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9164_ (.D(_0434_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9165_ (.D(_0435_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9166_ (.D(_0436_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9167_ (.D(_0437_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9168_ (.D(_0438_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9169_ (.D(_0439_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9170_ (.D(_0440_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9171_ (.D(_0441_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9172_ (.D(_0442_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9173_ (.D(_0443_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9174_ (.D(_0444_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9175_ (.D(_0445_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9176_ (.D(_0446_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9177_ (.D(_0447_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9178_ (.D(_0448_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9179_ (.D(_0449_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9180_ (.D(_0450_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9181_ (.D(_0451_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9182_ (.D(_0452_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9183_ (.D(_0453_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9184_ (.D(_0454_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9185_ (.D(_0455_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9186_ (.D(_0456_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9187_ (.D(_0457_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9188_ (.D(_0458_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9189_ (.D(_0459_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9190_ (.D(_0460_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9191_ (.D(_0461_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9192_ (.D(_0462_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9193_ (.D(_0463_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9194_ (.D(_0464_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9195_ (.D(_0465_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9196_ (.D(_0466_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9197_ (.D(_0467_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9198_ (.D(_0468_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9199_ (.D(_0469_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9200_ (.D(_0470_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9201_ (.D(_0471_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9202_ (.D(_0472_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9203_ (.D(_0473_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9204_ (.D(_0474_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9205_ (.D(_0475_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9206_ (.D(_0476_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9207_ (.D(_0477_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9208_ (.D(_0478_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9209_ (.D(_0479_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9210_ (.D(_0480_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[5][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9211_ (.D(_0481_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[5][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9212_ (.D(\pc_next[2] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9213_ (.D(\pc_next[3] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9214_ (.D(\pc_next[4] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9215_ (.D(\pc_next[5] ),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9216_ (.D(\pc_next[6] ),
    .CLK(clknet_leaf_63_clk),
    .Q(\pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9217_ (.D(\pc_next[7] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9218_ (.D(\pc_next[8] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9219_ (.D(\pc_next[9] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9220_ (.D(\pc_next[10] ),
    .CLK(clknet_leaf_61_clk),
    .Q(\pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9221_ (.D(\pc_next[11] ),
    .CLK(clknet_leaf_61_clk),
    .Q(\pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9222_ (.D(\pc_next[12] ),
    .CLK(clknet_leaf_61_clk),
    .Q(\pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9223_ (.D(\pc_next[13] ),
    .CLK(clknet_leaf_61_clk),
    .Q(\pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9224_ (.D(\pc_next[14] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9225_ (.D(\pc_next[15] ),
    .CLK(clknet_leaf_60_clk),
    .Q(\pc[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9226_ (.D(\pc_next[16] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\pc[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9227_ (.D(\pc_next[17] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\pc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9228_ (.D(\pc_next[18] ),
    .CLK(clknet_leaf_74_clk),
    .Q(\pc[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9229_ (.D(\pc_next[19] ),
    .CLK(clknet_leaf_74_clk),
    .Q(\pc[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9230_ (.D(\pc_next[20] ),
    .CLK(clknet_leaf_74_clk),
    .Q(\pc[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9231_ (.D(\pc_next[21] ),
    .CLK(clknet_leaf_75_clk),
    .Q(\pc[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9232_ (.D(\pc_next[22] ),
    .CLK(clknet_leaf_76_clk),
    .Q(\pc[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9233_ (.D(\pc_next[23] ),
    .CLK(clknet_leaf_76_clk),
    .Q(\pc[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9234_ (.D(\pc_next[24] ),
    .CLK(clknet_leaf_80_clk),
    .Q(\pc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9235_ (.D(\pc_next[25] ),
    .CLK(clknet_leaf_79_clk),
    .Q(\pc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9236_ (.D(\pc_next[26] ),
    .CLK(clknet_leaf_78_clk),
    .Q(\pc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9237_ (.D(\pc_next[27] ),
    .CLK(clknet_leaf_78_clk),
    .Q(\pc[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9238_ (.D(\pc_next[28] ),
    .CLK(clknet_leaf_78_clk),
    .Q(\pc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9239_ (.D(\pc_next[29] ),
    .CLK(clknet_leaf_77_clk),
    .Q(\pc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9240_ (.D(\pc_next[30] ),
    .CLK(clknet_leaf_77_clk),
    .Q(\pc[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9241_ (.D(\pc_next[31] ),
    .CLK(clknet_leaf_77_clk),
    .Q(\pc[31] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input1 (.I(inst_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(inst_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(inst_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(inst_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input13 (.I(inst_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(inst_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(inst_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(inst_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input17 (.I(inst_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(inst_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(inst_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(inst_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(inst_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(inst_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input22 (.I(inst_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input23 (.I(inst_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(inst_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(inst_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input26 (.I(inst_in[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input27 (.I(inst_in[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input28 (.I(inst_in[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input29 (.I(inst_in[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(inst_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(inst_in[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(inst_in[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input32 (.I(inst_in[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(mem_load_out[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(mem_load_out[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(mem_load_out[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(mem_load_out[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(mem_load_out[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(mem_load_out[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(mem_load_out[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(inst_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(mem_load_out[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(mem_load_out[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(mem_load_out[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(mem_load_out[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(mem_load_out[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(mem_load_out[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(mem_load_out[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(mem_load_out[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(mem_load_out[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(mem_load_out[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input5 (.I(inst_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(mem_load_out[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(mem_load_out[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(mem_load_out[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(mem_load_out[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(mem_load_out[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input55 (.I(mem_load_out[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(mem_load_out[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(mem_load_out[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input58 (.I(mem_load_out[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(mem_load_out[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(inst_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(mem_load_out[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(mem_load_out[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input62 (.I(mem_load_out[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(mem_load_out[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(mem_load_out[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(inst_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(inst_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(inst_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(alu_out_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output66 (.I(net66),
    .Z(alu_out_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output67 (.I(net67),
    .Z(alu_out_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output68 (.I(net68),
    .Z(alu_out_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output69 (.I(net69),
    .Z(alu_out_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output70 (.I(net70),
    .Z(alu_out_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output71 (.I(net71),
    .Z(alu_out_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output72 (.I(net72),
    .Z(alu_out_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output73 (.I(net73),
    .Z(alu_out_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output74 (.I(net74),
    .Z(alu_out_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(alu_out_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(alu_out_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output77 (.I(net77),
    .Z(alu_out_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output78 (.I(net78),
    .Z(alu_out_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output79 (.I(net79),
    .Z(alu_out_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output80 (.I(net80),
    .Z(alu_out_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output81 (.I(net81),
    .Z(alu_out_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output82 (.I(net82),
    .Z(alu_out_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output83 (.I(net83),
    .Z(alu_out_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output84 (.I(net84),
    .Z(alu_out_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output85 (.I(net85),
    .Z(alu_out_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output86 (.I(net86),
    .Z(alu_out_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output87 (.I(net87),
    .Z(alu_out_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output88 (.I(net88),
    .Z(alu_out_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output89 (.I(net89),
    .Z(alu_out_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output90 (.I(net90),
    .Z(alu_out_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output91 (.I(net91),
    .Z(alu_out_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output92 (.I(net92),
    .Z(alu_out_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output93 (.I(net93),
    .Z(alu_out_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output94 (.I(net94),
    .Z(alu_out_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output95 (.I(net95),
    .Z(alu_out_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output96 (.I(net96),
    .Z(alu_out_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer1 (.I(net98),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer10 (.I(_0513_),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(net106),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(_0549_),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(net108),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer14 (.I(_1956_),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(_0638_),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(_0545_),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer17 (.I(_0546_),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer18 (.I(_0546_),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer19 (.I(_0718_),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(net102),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer3 (.I(_1087_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer4 (.I(_1553_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(net100),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(_1553_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer7 (.I(_2133_),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer8 (.I(_1875_),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(_0932_),
    .Z(net105));
endmodule

