magic
tech gf180mcuD
magscale 1 5
timestamp 1700266060
<< obsm1 >>
rect 672 855 279328 174817
<< metal2 >>
rect 66640 175600 66696 176000
rect 66752 175600 66808 176000
rect 66864 175600 66920 176000
rect 68656 175600 68712 176000
rect 68768 175600 68824 176000
rect 68880 175600 68936 176000
rect 68992 175600 69048 176000
rect 69104 175600 69160 176000
rect 69216 175600 69272 176000
rect 71568 175600 71624 176000
rect 71680 175600 71736 176000
rect 71792 175600 71848 176000
rect 71904 175600 71960 176000
rect 72016 175600 72072 176000
rect 72128 175600 72184 176000
rect 72240 175600 72296 176000
rect 72352 175600 72408 176000
rect 75264 175600 75320 176000
rect 77056 175600 77112 176000
rect 77168 175600 77224 176000
rect 77280 175600 77336 176000
rect 77392 175600 77448 176000
rect 77504 175600 77560 176000
rect 78736 175600 78792 176000
rect 78848 175600 78904 176000
rect 78960 175600 79016 176000
rect 81312 175600 81368 176000
rect 81424 175600 81480 176000
rect 81536 175600 81592 176000
rect 81648 175600 81704 176000
rect 81760 175600 81816 176000
rect 81872 175600 81928 176000
rect 83104 175600 83160 176000
rect 83216 175600 83272 176000
rect 83328 175600 83384 176000
rect 85120 175600 85176 176000
rect 85232 175600 85288 176000
rect 85344 175600 85400 176000
rect 87136 175600 87192 176000
rect 87248 175600 87304 176000
rect 87360 175600 87416 176000
rect 87472 175600 87528 176000
rect 87584 175600 87640 176000
rect 87696 175600 87752 176000
rect 90048 175600 90104 176000
rect 90160 175600 90216 176000
rect 90272 175600 90328 176000
rect 90384 175600 90440 176000
rect 90496 175600 90552 176000
rect 90608 175600 90664 176000
rect 90720 175600 90776 176000
rect 90832 175600 90888 176000
rect 93744 175600 93800 176000
rect 95536 175600 95592 176000
rect 95648 175600 95704 176000
rect 95760 175600 95816 176000
rect 95872 175600 95928 176000
rect 95984 175600 96040 176000
rect 97216 175600 97272 176000
rect 97328 175600 97384 176000
rect 97440 175600 97496 176000
rect 99792 175600 99848 176000
rect 99904 175600 99960 176000
rect 100016 175600 100072 176000
rect 100128 175600 100184 176000
rect 100240 175600 100296 176000
rect 100352 175600 100408 176000
rect 101584 175600 101640 176000
rect 101696 175600 101752 176000
rect 101808 175600 101864 176000
rect 103600 175600 103656 176000
rect 103712 175600 103768 176000
rect 103824 175600 103880 176000
rect 105616 175600 105672 176000
rect 105728 175600 105784 176000
rect 105840 175600 105896 176000
rect 105952 175600 106008 176000
rect 106064 175600 106120 176000
rect 106176 175600 106232 176000
rect 108528 175600 108584 176000
rect 108640 175600 108696 176000
rect 108752 175600 108808 176000
rect 108864 175600 108920 176000
rect 108976 175600 109032 176000
rect 109088 175600 109144 176000
rect 109200 175600 109256 176000
rect 109312 175600 109368 176000
rect 112224 175600 112280 176000
rect 114016 175600 114072 176000
rect 114128 175600 114184 176000
rect 114240 175600 114296 176000
rect 114352 175600 114408 176000
rect 114464 175600 114520 176000
rect 115696 175600 115752 176000
rect 115808 175600 115864 176000
rect 115920 175600 115976 176000
rect 118272 175600 118328 176000
rect 118384 175600 118440 176000
rect 118496 175600 118552 176000
rect 118608 175600 118664 176000
rect 118720 175600 118776 176000
rect 118832 175600 118888 176000
rect 120064 175600 120120 176000
rect 120176 175600 120232 176000
rect 120288 175600 120344 176000
rect 122080 175600 122136 176000
rect 122192 175600 122248 176000
rect 122304 175600 122360 176000
rect 124096 175600 124152 176000
rect 124208 175600 124264 176000
rect 124320 175600 124376 176000
rect 124432 175600 124488 176000
rect 124544 175600 124600 176000
rect 124656 175600 124712 176000
rect 127008 175600 127064 176000
rect 127120 175600 127176 176000
rect 127232 175600 127288 176000
rect 127344 175600 127400 176000
rect 127456 175600 127512 176000
rect 127568 175600 127624 176000
rect 127680 175600 127736 176000
rect 127792 175600 127848 176000
rect 130704 175600 130760 176000
rect 132496 175600 132552 176000
rect 132608 175600 132664 176000
rect 132720 175600 132776 176000
rect 132832 175600 132888 176000
rect 132944 175600 133000 176000
rect 134176 175600 134232 176000
rect 134288 175600 134344 176000
rect 134400 175600 134456 176000
rect 136752 175600 136808 176000
rect 136864 175600 136920 176000
rect 136976 175600 137032 176000
rect 137088 175600 137144 176000
rect 137200 175600 137256 176000
rect 137312 175600 137368 176000
rect 138544 175600 138600 176000
rect 138656 175600 138712 176000
rect 138768 175600 138824 176000
rect 140560 175600 140616 176000
rect 140672 175600 140728 176000
rect 140784 175600 140840 176000
rect 142576 175600 142632 176000
rect 142688 175600 142744 176000
rect 142800 175600 142856 176000
rect 142912 175600 142968 176000
rect 143024 175600 143080 176000
rect 143136 175600 143192 176000
rect 145488 175600 145544 176000
rect 145600 175600 145656 176000
rect 145712 175600 145768 176000
rect 145824 175600 145880 176000
rect 145936 175600 145992 176000
rect 146048 175600 146104 176000
rect 146160 175600 146216 176000
rect 146272 175600 146328 176000
rect 149184 175600 149240 176000
rect 150976 175600 151032 176000
rect 151088 175600 151144 176000
rect 151200 175600 151256 176000
rect 151312 175600 151368 176000
rect 151424 175600 151480 176000
rect 152656 175600 152712 176000
rect 152768 175600 152824 176000
rect 152880 175600 152936 176000
rect 155232 175600 155288 176000
rect 155344 175600 155400 176000
rect 155456 175600 155512 176000
rect 155568 175600 155624 176000
rect 155680 175600 155736 176000
rect 155792 175600 155848 176000
rect 157024 175600 157080 176000
rect 157136 175600 157192 176000
rect 157248 175600 157304 176000
rect 159040 175600 159096 176000
rect 159152 175600 159208 176000
rect 159264 175600 159320 176000
rect 161056 175600 161112 176000
rect 161168 175600 161224 176000
rect 161280 175600 161336 176000
rect 161392 175600 161448 176000
rect 161504 175600 161560 176000
rect 161616 175600 161672 176000
rect 163968 175600 164024 176000
rect 164080 175600 164136 176000
rect 164192 175600 164248 176000
rect 164304 175600 164360 176000
rect 164416 175600 164472 176000
rect 164528 175600 164584 176000
rect 164640 175600 164696 176000
rect 164752 175600 164808 176000
rect 167664 175600 167720 176000
rect 169456 175600 169512 176000
rect 169568 175600 169624 176000
rect 169680 175600 169736 176000
rect 169792 175600 169848 176000
rect 169904 175600 169960 176000
rect 171136 175600 171192 176000
rect 171248 175600 171304 176000
rect 171360 175600 171416 176000
rect 173712 175600 173768 176000
rect 173824 175600 173880 176000
rect 173936 175600 173992 176000
rect 174048 175600 174104 176000
rect 174160 175600 174216 176000
rect 174272 175600 174328 176000
rect 175504 175600 175560 176000
rect 175616 175600 175672 176000
rect 175728 175600 175784 176000
rect 177520 175600 177576 176000
rect 177632 175600 177688 176000
rect 177744 175600 177800 176000
rect 179536 175600 179592 176000
rect 179648 175600 179704 176000
rect 179760 175600 179816 176000
rect 179872 175600 179928 176000
rect 179984 175600 180040 176000
rect 180096 175600 180152 176000
rect 182448 175600 182504 176000
rect 182560 175600 182616 176000
rect 182672 175600 182728 176000
rect 182784 175600 182840 176000
rect 182896 175600 182952 176000
rect 183008 175600 183064 176000
rect 183120 175600 183176 176000
rect 183232 175600 183288 176000
rect 186144 175600 186200 176000
rect 187936 175600 187992 176000
rect 188048 175600 188104 176000
rect 188160 175600 188216 176000
rect 188272 175600 188328 176000
rect 188384 175600 188440 176000
rect 189616 175600 189672 176000
rect 189728 175600 189784 176000
rect 189840 175600 189896 176000
rect 192192 175600 192248 176000
rect 192304 175600 192360 176000
rect 192416 175600 192472 176000
rect 192528 175600 192584 176000
rect 192640 175600 192696 176000
rect 192752 175600 192808 176000
rect 193984 175600 194040 176000
rect 194096 175600 194152 176000
rect 194208 175600 194264 176000
rect 196000 175600 196056 176000
rect 196112 175600 196168 176000
rect 196224 175600 196280 176000
rect 198016 175600 198072 176000
rect 198128 175600 198184 176000
rect 198240 175600 198296 176000
rect 198352 175600 198408 176000
rect 198464 175600 198520 176000
rect 198576 175600 198632 176000
rect 200928 175600 200984 176000
rect 201040 175600 201096 176000
rect 201152 175600 201208 176000
rect 201264 175600 201320 176000
rect 201376 175600 201432 176000
rect 201488 175600 201544 176000
rect 201600 175600 201656 176000
rect 201712 175600 201768 176000
rect 204624 175600 204680 176000
rect 206416 175600 206472 176000
rect 206528 175600 206584 176000
rect 206640 175600 206696 176000
rect 206752 175600 206808 176000
rect 206864 175600 206920 176000
rect 208096 175600 208152 176000
rect 208208 175600 208264 176000
rect 208320 175600 208376 176000
rect 210672 175600 210728 176000
rect 210784 175600 210840 176000
rect 210896 175600 210952 176000
rect 211008 175600 211064 176000
rect 211120 175600 211176 176000
rect 211232 175600 211288 176000
rect 212464 175600 212520 176000
rect 212576 175600 212632 176000
rect 212688 175600 212744 176000
rect 5488 0 5544 400
rect 6384 0 6440 400
rect 7280 0 7336 400
rect 8176 0 8232 400
rect 9072 0 9128 400
rect 9968 0 10024 400
rect 10864 0 10920 400
rect 11760 0 11816 400
rect 12656 0 12712 400
rect 13552 0 13608 400
rect 14448 0 14504 400
rect 15344 0 15400 400
rect 16240 0 16296 400
rect 17136 0 17192 400
rect 18032 0 18088 400
rect 18928 0 18984 400
rect 19824 0 19880 400
rect 20720 0 20776 400
rect 21616 0 21672 400
rect 22512 0 22568 400
rect 23408 0 23464 400
rect 24304 0 24360 400
rect 25200 0 25256 400
rect 26096 0 26152 400
rect 26992 0 27048 400
rect 27888 0 27944 400
rect 28784 0 28840 400
rect 29680 0 29736 400
rect 30576 0 30632 400
rect 31472 0 31528 400
rect 32368 0 32424 400
rect 33264 0 33320 400
rect 34160 0 34216 400
rect 35056 0 35112 400
rect 35952 0 36008 400
rect 36848 0 36904 400
rect 37744 0 37800 400
rect 38640 0 38696 400
rect 39536 0 39592 400
rect 40432 0 40488 400
rect 41328 0 41384 400
rect 42224 0 42280 400
rect 43120 0 43176 400
rect 44016 0 44072 400
rect 44912 0 44968 400
rect 45808 0 45864 400
rect 46704 0 46760 400
rect 47600 0 47656 400
rect 48496 0 48552 400
rect 49392 0 49448 400
rect 50288 0 50344 400
rect 51184 0 51240 400
rect 52080 0 52136 400
rect 52976 0 53032 400
rect 53872 0 53928 400
rect 54768 0 54824 400
rect 55664 0 55720 400
rect 56560 0 56616 400
rect 57456 0 57512 400
rect 58352 0 58408 400
rect 59248 0 59304 400
rect 60144 0 60200 400
rect 61040 0 61096 400
rect 61936 0 61992 400
rect 62832 0 62888 400
rect 63728 0 63784 400
rect 64624 0 64680 400
rect 65520 0 65576 400
rect 66416 0 66472 400
rect 67312 0 67368 400
rect 68208 0 68264 400
rect 69104 0 69160 400
rect 70000 0 70056 400
rect 70896 0 70952 400
rect 71792 0 71848 400
rect 72688 0 72744 400
rect 73584 0 73640 400
rect 74480 0 74536 400
rect 75376 0 75432 400
rect 76272 0 76328 400
rect 77168 0 77224 400
rect 78064 0 78120 400
rect 78960 0 79016 400
rect 79856 0 79912 400
rect 80752 0 80808 400
rect 81648 0 81704 400
rect 82544 0 82600 400
rect 83440 0 83496 400
rect 84336 0 84392 400
rect 85232 0 85288 400
rect 86128 0 86184 400
rect 87024 0 87080 400
rect 87920 0 87976 400
rect 88816 0 88872 400
rect 89712 0 89768 400
rect 90608 0 90664 400
rect 91504 0 91560 400
rect 92400 0 92456 400
rect 93296 0 93352 400
rect 94192 0 94248 400
rect 95088 0 95144 400
rect 95984 0 96040 400
rect 96880 0 96936 400
rect 97776 0 97832 400
rect 98672 0 98728 400
rect 99568 0 99624 400
rect 100464 0 100520 400
rect 101360 0 101416 400
rect 102256 0 102312 400
rect 103152 0 103208 400
rect 104048 0 104104 400
rect 104944 0 105000 400
rect 105840 0 105896 400
rect 106736 0 106792 400
rect 107632 0 107688 400
rect 108528 0 108584 400
rect 109424 0 109480 400
rect 110320 0 110376 400
rect 111216 0 111272 400
rect 112112 0 112168 400
rect 113008 0 113064 400
rect 113904 0 113960 400
rect 114800 0 114856 400
rect 115696 0 115752 400
rect 116592 0 116648 400
rect 117488 0 117544 400
rect 118384 0 118440 400
rect 119280 0 119336 400
rect 120176 0 120232 400
rect 121072 0 121128 400
rect 121968 0 122024 400
rect 122864 0 122920 400
rect 123760 0 123816 400
rect 124656 0 124712 400
rect 125552 0 125608 400
rect 126448 0 126504 400
rect 127344 0 127400 400
rect 128240 0 128296 400
rect 129136 0 129192 400
rect 130032 0 130088 400
rect 130928 0 130984 400
rect 131824 0 131880 400
rect 132720 0 132776 400
rect 133616 0 133672 400
rect 134512 0 134568 400
rect 135408 0 135464 400
rect 136304 0 136360 400
rect 137200 0 137256 400
rect 138096 0 138152 400
rect 138992 0 139048 400
rect 139888 0 139944 400
rect 140784 0 140840 400
rect 141680 0 141736 400
rect 142576 0 142632 400
rect 143472 0 143528 400
rect 144368 0 144424 400
rect 145264 0 145320 400
rect 146160 0 146216 400
rect 147056 0 147112 400
rect 147952 0 148008 400
rect 148848 0 148904 400
rect 149744 0 149800 400
rect 150640 0 150696 400
rect 151536 0 151592 400
rect 152432 0 152488 400
rect 153328 0 153384 400
rect 154224 0 154280 400
rect 155120 0 155176 400
rect 156016 0 156072 400
rect 156912 0 156968 400
rect 157808 0 157864 400
rect 158704 0 158760 400
rect 159600 0 159656 400
rect 160496 0 160552 400
rect 161392 0 161448 400
rect 162288 0 162344 400
rect 163184 0 163240 400
rect 164080 0 164136 400
rect 164976 0 165032 400
rect 165872 0 165928 400
rect 166768 0 166824 400
rect 167664 0 167720 400
rect 168560 0 168616 400
rect 169456 0 169512 400
rect 170352 0 170408 400
rect 171248 0 171304 400
rect 172144 0 172200 400
rect 173040 0 173096 400
rect 173936 0 173992 400
rect 174832 0 174888 400
rect 175728 0 175784 400
rect 176624 0 176680 400
rect 177520 0 177576 400
rect 178416 0 178472 400
rect 179312 0 179368 400
rect 180208 0 180264 400
rect 181104 0 181160 400
rect 182000 0 182056 400
rect 182896 0 182952 400
rect 183792 0 183848 400
rect 184688 0 184744 400
rect 185584 0 185640 400
rect 186480 0 186536 400
rect 187376 0 187432 400
rect 188272 0 188328 400
rect 189168 0 189224 400
rect 190064 0 190120 400
rect 190960 0 191016 400
rect 191856 0 191912 400
rect 192752 0 192808 400
rect 193648 0 193704 400
rect 194544 0 194600 400
rect 195440 0 195496 400
rect 196336 0 196392 400
rect 197232 0 197288 400
rect 198128 0 198184 400
rect 199024 0 199080 400
rect 199920 0 199976 400
rect 200816 0 200872 400
rect 201712 0 201768 400
rect 202608 0 202664 400
rect 203504 0 203560 400
rect 204400 0 204456 400
rect 205296 0 205352 400
rect 206192 0 206248 400
rect 207088 0 207144 400
rect 207984 0 208040 400
rect 208880 0 208936 400
rect 209776 0 209832 400
rect 210672 0 210728 400
rect 211568 0 211624 400
rect 212464 0 212520 400
rect 213360 0 213416 400
rect 214256 0 214312 400
rect 215152 0 215208 400
rect 216048 0 216104 400
rect 216944 0 217000 400
rect 217840 0 217896 400
rect 218736 0 218792 400
rect 219632 0 219688 400
rect 220528 0 220584 400
rect 221424 0 221480 400
rect 222320 0 222376 400
rect 223216 0 223272 400
rect 224112 0 224168 400
rect 225008 0 225064 400
rect 225904 0 225960 400
rect 226800 0 226856 400
rect 227696 0 227752 400
rect 228592 0 228648 400
rect 229488 0 229544 400
rect 230384 0 230440 400
rect 231280 0 231336 400
rect 232176 0 232232 400
rect 233072 0 233128 400
rect 233968 0 234024 400
rect 234864 0 234920 400
rect 235760 0 235816 400
rect 236656 0 236712 400
rect 237552 0 237608 400
rect 238448 0 238504 400
rect 239344 0 239400 400
rect 240240 0 240296 400
rect 241136 0 241192 400
rect 242032 0 242088 400
rect 242928 0 242984 400
rect 243824 0 243880 400
rect 244720 0 244776 400
rect 245616 0 245672 400
rect 246512 0 246568 400
rect 247408 0 247464 400
rect 248304 0 248360 400
rect 249200 0 249256 400
rect 250096 0 250152 400
rect 250992 0 251048 400
rect 251888 0 251944 400
rect 252784 0 252840 400
rect 253680 0 253736 400
rect 254576 0 254632 400
rect 255472 0 255528 400
rect 256368 0 256424 400
rect 257264 0 257320 400
rect 258160 0 258216 400
rect 259056 0 259112 400
rect 259952 0 260008 400
rect 260848 0 260904 400
rect 261744 0 261800 400
rect 262640 0 262696 400
rect 263536 0 263592 400
rect 264432 0 264488 400
rect 265328 0 265384 400
rect 266224 0 266280 400
rect 267120 0 267176 400
rect 268016 0 268072 400
rect 268912 0 268968 400
rect 269808 0 269864 400
rect 270704 0 270760 400
rect 271600 0 271656 400
rect 272496 0 272552 400
rect 273392 0 273448 400
rect 274288 0 274344 400
<< obsm2 >>
rect 854 175570 66610 175658
rect 66950 175570 68626 175658
rect 69302 175570 71538 175658
rect 72438 175570 75234 175658
rect 75350 175570 77026 175658
rect 77590 175570 78706 175658
rect 79046 175570 81282 175658
rect 81958 175570 83074 175658
rect 83414 175570 85090 175658
rect 85430 175570 87106 175658
rect 87782 175570 90018 175658
rect 90918 175570 93714 175658
rect 93830 175570 95506 175658
rect 96070 175570 97186 175658
rect 97526 175570 99762 175658
rect 100438 175570 101554 175658
rect 101894 175570 103570 175658
rect 103910 175570 105586 175658
rect 106262 175570 108498 175658
rect 109398 175570 112194 175658
rect 112310 175570 113986 175658
rect 114550 175570 115666 175658
rect 116006 175570 118242 175658
rect 118918 175570 120034 175658
rect 120374 175570 122050 175658
rect 122390 175570 124066 175658
rect 124742 175570 126978 175658
rect 127878 175570 130674 175658
rect 130790 175570 132466 175658
rect 133030 175570 134146 175658
rect 134486 175570 136722 175658
rect 137398 175570 138514 175658
rect 138854 175570 140530 175658
rect 140870 175570 142546 175658
rect 143222 175570 145458 175658
rect 146358 175570 149154 175658
rect 149270 175570 150946 175658
rect 151510 175570 152626 175658
rect 152966 175570 155202 175658
rect 155878 175570 156994 175658
rect 157334 175570 159010 175658
rect 159350 175570 161026 175658
rect 161702 175570 163938 175658
rect 164838 175570 167634 175658
rect 167750 175570 169426 175658
rect 169990 175570 171106 175658
rect 171446 175570 173682 175658
rect 174358 175570 175474 175658
rect 175814 175570 177490 175658
rect 177830 175570 179506 175658
rect 180182 175570 182418 175658
rect 183318 175570 186114 175658
rect 186230 175570 187906 175658
rect 188470 175570 189586 175658
rect 189926 175570 192162 175658
rect 192838 175570 193954 175658
rect 194294 175570 195970 175658
rect 196310 175570 197986 175658
rect 198662 175570 200898 175658
rect 201798 175570 204594 175658
rect 204710 175570 206386 175658
rect 206950 175570 208066 175658
rect 208406 175570 210642 175658
rect 211318 175570 212434 175658
rect 212774 175570 279146 175658
rect 854 430 279146 175570
rect 854 350 5458 430
rect 5574 350 6354 430
rect 6470 350 7250 430
rect 7366 350 8146 430
rect 8262 350 9042 430
rect 9158 350 9938 430
rect 10054 350 10834 430
rect 10950 350 11730 430
rect 11846 350 12626 430
rect 12742 350 13522 430
rect 13638 350 14418 430
rect 14534 350 15314 430
rect 15430 350 16210 430
rect 16326 350 17106 430
rect 17222 350 18002 430
rect 18118 350 18898 430
rect 19014 350 19794 430
rect 19910 350 20690 430
rect 20806 350 21586 430
rect 21702 350 22482 430
rect 22598 350 23378 430
rect 23494 350 24274 430
rect 24390 350 25170 430
rect 25286 350 26066 430
rect 26182 350 26962 430
rect 27078 350 27858 430
rect 27974 350 28754 430
rect 28870 350 29650 430
rect 29766 350 30546 430
rect 30662 350 31442 430
rect 31558 350 32338 430
rect 32454 350 33234 430
rect 33350 350 34130 430
rect 34246 350 35026 430
rect 35142 350 35922 430
rect 36038 350 36818 430
rect 36934 350 37714 430
rect 37830 350 38610 430
rect 38726 350 39506 430
rect 39622 350 40402 430
rect 40518 350 41298 430
rect 41414 350 42194 430
rect 42310 350 43090 430
rect 43206 350 43986 430
rect 44102 350 44882 430
rect 44998 350 45778 430
rect 45894 350 46674 430
rect 46790 350 47570 430
rect 47686 350 48466 430
rect 48582 350 49362 430
rect 49478 350 50258 430
rect 50374 350 51154 430
rect 51270 350 52050 430
rect 52166 350 52946 430
rect 53062 350 53842 430
rect 53958 350 54738 430
rect 54854 350 55634 430
rect 55750 350 56530 430
rect 56646 350 57426 430
rect 57542 350 58322 430
rect 58438 350 59218 430
rect 59334 350 60114 430
rect 60230 350 61010 430
rect 61126 350 61906 430
rect 62022 350 62802 430
rect 62918 350 63698 430
rect 63814 350 64594 430
rect 64710 350 65490 430
rect 65606 350 66386 430
rect 66502 350 67282 430
rect 67398 350 68178 430
rect 68294 350 69074 430
rect 69190 350 69970 430
rect 70086 350 70866 430
rect 70982 350 71762 430
rect 71878 350 72658 430
rect 72774 350 73554 430
rect 73670 350 74450 430
rect 74566 350 75346 430
rect 75462 350 76242 430
rect 76358 350 77138 430
rect 77254 350 78034 430
rect 78150 350 78930 430
rect 79046 350 79826 430
rect 79942 350 80722 430
rect 80838 350 81618 430
rect 81734 350 82514 430
rect 82630 350 83410 430
rect 83526 350 84306 430
rect 84422 350 85202 430
rect 85318 350 86098 430
rect 86214 350 86994 430
rect 87110 350 87890 430
rect 88006 350 88786 430
rect 88902 350 89682 430
rect 89798 350 90578 430
rect 90694 350 91474 430
rect 91590 350 92370 430
rect 92486 350 93266 430
rect 93382 350 94162 430
rect 94278 350 95058 430
rect 95174 350 95954 430
rect 96070 350 96850 430
rect 96966 350 97746 430
rect 97862 350 98642 430
rect 98758 350 99538 430
rect 99654 350 100434 430
rect 100550 350 101330 430
rect 101446 350 102226 430
rect 102342 350 103122 430
rect 103238 350 104018 430
rect 104134 350 104914 430
rect 105030 350 105810 430
rect 105926 350 106706 430
rect 106822 350 107602 430
rect 107718 350 108498 430
rect 108614 350 109394 430
rect 109510 350 110290 430
rect 110406 350 111186 430
rect 111302 350 112082 430
rect 112198 350 112978 430
rect 113094 350 113874 430
rect 113990 350 114770 430
rect 114886 350 115666 430
rect 115782 350 116562 430
rect 116678 350 117458 430
rect 117574 350 118354 430
rect 118470 350 119250 430
rect 119366 350 120146 430
rect 120262 350 121042 430
rect 121158 350 121938 430
rect 122054 350 122834 430
rect 122950 350 123730 430
rect 123846 350 124626 430
rect 124742 350 125522 430
rect 125638 350 126418 430
rect 126534 350 127314 430
rect 127430 350 128210 430
rect 128326 350 129106 430
rect 129222 350 130002 430
rect 130118 350 130898 430
rect 131014 350 131794 430
rect 131910 350 132690 430
rect 132806 350 133586 430
rect 133702 350 134482 430
rect 134598 350 135378 430
rect 135494 350 136274 430
rect 136390 350 137170 430
rect 137286 350 138066 430
rect 138182 350 138962 430
rect 139078 350 139858 430
rect 139974 350 140754 430
rect 140870 350 141650 430
rect 141766 350 142546 430
rect 142662 350 143442 430
rect 143558 350 144338 430
rect 144454 350 145234 430
rect 145350 350 146130 430
rect 146246 350 147026 430
rect 147142 350 147922 430
rect 148038 350 148818 430
rect 148934 350 149714 430
rect 149830 350 150610 430
rect 150726 350 151506 430
rect 151622 350 152402 430
rect 152518 350 153298 430
rect 153414 350 154194 430
rect 154310 350 155090 430
rect 155206 350 155986 430
rect 156102 350 156882 430
rect 156998 350 157778 430
rect 157894 350 158674 430
rect 158790 350 159570 430
rect 159686 350 160466 430
rect 160582 350 161362 430
rect 161478 350 162258 430
rect 162374 350 163154 430
rect 163270 350 164050 430
rect 164166 350 164946 430
rect 165062 350 165842 430
rect 165958 350 166738 430
rect 166854 350 167634 430
rect 167750 350 168530 430
rect 168646 350 169426 430
rect 169542 350 170322 430
rect 170438 350 171218 430
rect 171334 350 172114 430
rect 172230 350 173010 430
rect 173126 350 173906 430
rect 174022 350 174802 430
rect 174918 350 175698 430
rect 175814 350 176594 430
rect 176710 350 177490 430
rect 177606 350 178386 430
rect 178502 350 179282 430
rect 179398 350 180178 430
rect 180294 350 181074 430
rect 181190 350 181970 430
rect 182086 350 182866 430
rect 182982 350 183762 430
rect 183878 350 184658 430
rect 184774 350 185554 430
rect 185670 350 186450 430
rect 186566 350 187346 430
rect 187462 350 188242 430
rect 188358 350 189138 430
rect 189254 350 190034 430
rect 190150 350 190930 430
rect 191046 350 191826 430
rect 191942 350 192722 430
rect 192838 350 193618 430
rect 193734 350 194514 430
rect 194630 350 195410 430
rect 195526 350 196306 430
rect 196422 350 197202 430
rect 197318 350 198098 430
rect 198214 350 198994 430
rect 199110 350 199890 430
rect 200006 350 200786 430
rect 200902 350 201682 430
rect 201798 350 202578 430
rect 202694 350 203474 430
rect 203590 350 204370 430
rect 204486 350 205266 430
rect 205382 350 206162 430
rect 206278 350 207058 430
rect 207174 350 207954 430
rect 208070 350 208850 430
rect 208966 350 209746 430
rect 209862 350 210642 430
rect 210758 350 211538 430
rect 211654 350 212434 430
rect 212550 350 213330 430
rect 213446 350 214226 430
rect 214342 350 215122 430
rect 215238 350 216018 430
rect 216134 350 216914 430
rect 217030 350 217810 430
rect 217926 350 218706 430
rect 218822 350 219602 430
rect 219718 350 220498 430
rect 220614 350 221394 430
rect 221510 350 222290 430
rect 222406 350 223186 430
rect 223302 350 224082 430
rect 224198 350 224978 430
rect 225094 350 225874 430
rect 225990 350 226770 430
rect 226886 350 227666 430
rect 227782 350 228562 430
rect 228678 350 229458 430
rect 229574 350 230354 430
rect 230470 350 231250 430
rect 231366 350 232146 430
rect 232262 350 233042 430
rect 233158 350 233938 430
rect 234054 350 234834 430
rect 234950 350 235730 430
rect 235846 350 236626 430
rect 236742 350 237522 430
rect 237638 350 238418 430
rect 238534 350 239314 430
rect 239430 350 240210 430
rect 240326 350 241106 430
rect 241222 350 242002 430
rect 242118 350 242898 430
rect 243014 350 243794 430
rect 243910 350 244690 430
rect 244806 350 245586 430
rect 245702 350 246482 430
rect 246598 350 247378 430
rect 247494 350 248274 430
rect 248390 350 249170 430
rect 249286 350 250066 430
rect 250182 350 250962 430
rect 251078 350 251858 430
rect 251974 350 252754 430
rect 252870 350 253650 430
rect 253766 350 254546 430
rect 254662 350 255442 430
rect 255558 350 256338 430
rect 256454 350 257234 430
rect 257350 350 258130 430
rect 258246 350 259026 430
rect 259142 350 259922 430
rect 260038 350 260818 430
rect 260934 350 261714 430
rect 261830 350 262610 430
rect 262726 350 263506 430
rect 263622 350 264402 430
rect 264518 350 265298 430
rect 265414 350 266194 430
rect 266310 350 267090 430
rect 267206 350 267986 430
rect 268102 350 268882 430
rect 268998 350 269778 430
rect 269894 350 270674 430
rect 270790 350 271570 430
rect 271686 350 272466 430
rect 272582 350 273362 430
rect 273478 350 274258 430
rect 274374 350 279146 430
<< metal3 >>
rect 0 171696 400 171752
rect 279600 171696 280000 171752
rect 0 164416 400 164472
rect 279600 164416 280000 164472
rect 0 157136 400 157192
rect 279600 157136 280000 157192
rect 0 149856 400 149912
rect 279600 149856 280000 149912
rect 0 142576 400 142632
rect 279600 142576 280000 142632
rect 0 135296 400 135352
rect 279600 135296 280000 135352
rect 0 128016 400 128072
rect 279600 128016 280000 128072
rect 0 120736 400 120792
rect 279600 120736 280000 120792
rect 0 113456 400 113512
rect 279600 113456 280000 113512
rect 0 106176 400 106232
rect 279600 106176 280000 106232
rect 0 98896 400 98952
rect 279600 98896 280000 98952
rect 0 91616 400 91672
rect 279600 91616 280000 91672
rect 0 84336 400 84392
rect 279600 84336 280000 84392
rect 0 77056 400 77112
rect 279600 77056 280000 77112
rect 0 69776 400 69832
rect 279600 69776 280000 69832
rect 0 62496 400 62552
rect 279600 62496 280000 62552
rect 0 55216 400 55272
rect 279600 55216 280000 55272
rect 0 47936 400 47992
rect 279600 47936 280000 47992
rect 0 40656 400 40712
rect 279600 40656 280000 40712
rect 0 33376 400 33432
rect 279600 33376 280000 33432
rect 0 26096 400 26152
rect 279600 26096 280000 26152
rect 0 18816 400 18872
rect 279600 18816 280000 18872
rect 0 11536 400 11592
rect 279600 11536 280000 11592
rect 0 4256 400 4312
rect 279600 4256 280000 4312
<< obsm3 >>
rect 400 171782 279600 174706
rect 430 171666 279570 171782
rect 400 164502 279600 171666
rect 430 164386 279570 164502
rect 400 157222 279600 164386
rect 430 157106 279570 157222
rect 400 149942 279600 157106
rect 430 149826 279570 149942
rect 400 142662 279600 149826
rect 430 142546 279570 142662
rect 400 135382 279600 142546
rect 430 135266 279570 135382
rect 400 128102 279600 135266
rect 430 127986 279570 128102
rect 400 120822 279600 127986
rect 430 120706 279570 120822
rect 400 113542 279600 120706
rect 430 113426 279570 113542
rect 400 106262 279600 113426
rect 430 106146 279570 106262
rect 400 98982 279600 106146
rect 430 98866 279570 98982
rect 400 91702 279600 98866
rect 430 91586 279570 91702
rect 400 84422 279600 91586
rect 430 84306 279570 84422
rect 400 77142 279600 84306
rect 430 77026 279570 77142
rect 400 69862 279600 77026
rect 430 69746 279570 69862
rect 400 62582 279600 69746
rect 430 62466 279570 62582
rect 400 55302 279600 62466
rect 430 55186 279570 55302
rect 400 48022 279600 55186
rect 430 47906 279570 48022
rect 400 40742 279600 47906
rect 430 40626 279570 40742
rect 400 33462 279600 40626
rect 430 33346 279570 33462
rect 400 26182 279600 33346
rect 430 26066 279570 26182
rect 400 18902 279600 26066
rect 430 18786 279570 18902
rect 400 11622 279600 18786
rect 430 11506 279570 11622
rect 400 4342 279600 11506
rect 430 4226 279570 4342
rect 400 1554 279600 4226
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< labels >>
rlabel metal3 s 279600 4256 280000 4312 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 128016 400 128072 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 106176 400 106232 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 84336 400 84392 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 62496 400 62552 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 40656 400 40712 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 279600 26096 280000 26152 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 279600 47936 280000 47992 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 279600 69776 280000 69832 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 279600 91616 280000 91672 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 279600 113456 280000 113512 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 279600 135296 280000 135352 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 279600 157136 280000 157192 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 171696 400 171752 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 149856 400 149912 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 279600 18816 280000 18872 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 113456 400 113512 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 91616 400 91672 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 69776 400 69832 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 47936 400 47992 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 26096 400 26152 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 279600 40656 280000 40712 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 279600 62496 280000 62552 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 279600 84336 280000 84392 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 279600 106176 280000 106232 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 279600 128016 280000 128072 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 279600 149856 280000 149912 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 279600 171696 280000 171752 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 157136 400 157192 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 135296 400 135352 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 279600 11536 280000 11592 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 120736 400 120792 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 98896 400 98952 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 77056 400 77112 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 55216 400 55272 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 33376 400 33432 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 279600 33376 280000 33432 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 279600 55216 280000 55272 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 279600 77056 280000 77112 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 279600 98896 280000 98952 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 279600 120736 280000 120792 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 279600 142576 280000 142632 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 279600 164416 280000 164472 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 164416 400 164472 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 142576 400 142632 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 272496 0 272552 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 273392 0 273448 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 274288 0 274344 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 100464 0 100520 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 127344 0 127400 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 130032 0 130088 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 132720 0 132776 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 138096 0 138152 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 140784 0 140840 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 143472 0 143528 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 146160 0 146216 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 148848 0 148904 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 151536 0 151592 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 103152 0 103208 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 154224 0 154280 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 156912 0 156968 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 159600 0 159656 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 162288 0 162344 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 164976 0 165032 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 167664 0 167720 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 170352 0 170408 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 173040 0 173096 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 175728 0 175784 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 178416 0 178472 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 105840 0 105896 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 181104 0 181160 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 183792 0 183848 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 186480 0 186536 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 189168 0 189224 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 191856 0 191912 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 194544 0 194600 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 197232 0 197288 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 199920 0 199976 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 202608 0 202664 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 205296 0 205352 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 108528 0 108584 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 207984 0 208040 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 210672 0 210728 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 213360 0 213416 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 216048 0 216104 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 218736 0 218792 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 221424 0 221480 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 224112 0 224168 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 226800 0 226856 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 229488 0 229544 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 232176 0 232232 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 111216 0 111272 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 234864 0 234920 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 237552 0 237608 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 240240 0 240296 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 242928 0 242984 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 245616 0 245672 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 248304 0 248360 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 250992 0 251048 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 253680 0 253736 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 256368 0 256424 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 259056 0 259112 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 113904 0 113960 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 261744 0 261800 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 264432 0 264488 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 267120 0 267176 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 269808 0 269864 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 116592 0 116648 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 119280 0 119336 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 121968 0 122024 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 124656 0 124712 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 101360 0 101416 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 128240 0 128296 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 130928 0 130984 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 133616 0 133672 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 136304 0 136360 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 138992 0 139048 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 141680 0 141736 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 144368 0 144424 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 147056 0 147112 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 149744 0 149800 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 152432 0 152488 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 104048 0 104104 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 155120 0 155176 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 157808 0 157864 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 160496 0 160552 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 163184 0 163240 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 165872 0 165928 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 168560 0 168616 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 171248 0 171304 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 173936 0 173992 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 176624 0 176680 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 179312 0 179368 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 106736 0 106792 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 182000 0 182056 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 184688 0 184744 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 187376 0 187432 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 190064 0 190120 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 192752 0 192808 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 195440 0 195496 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 198128 0 198184 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 200816 0 200872 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 203504 0 203560 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 206192 0 206248 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 208880 0 208936 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 211568 0 211624 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 214256 0 214312 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 216944 0 217000 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 219632 0 219688 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 222320 0 222376 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 225008 0 225064 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 227696 0 227752 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 230384 0 230440 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 233072 0 233128 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 112112 0 112168 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 235760 0 235816 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 238448 0 238504 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 241136 0 241192 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 243824 0 243880 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 246512 0 246568 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 249200 0 249256 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 251888 0 251944 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 254576 0 254632 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 257264 0 257320 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 259952 0 260008 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 114800 0 114856 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 262640 0 262696 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 265328 0 265384 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 268016 0 268072 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 270704 0 270760 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 120176 0 120232 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 122864 0 122920 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 125552 0 125608 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 102256 0 102312 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 129136 0 129192 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 131824 0 131880 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 134512 0 134568 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 137200 0 137256 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 142576 0 142632 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 145264 0 145320 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 147952 0 148008 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 150640 0 150696 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 153328 0 153384 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 104944 0 105000 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 156016 0 156072 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 158704 0 158760 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 161392 0 161448 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 164080 0 164136 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 166768 0 166824 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 169456 0 169512 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 172144 0 172200 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 174832 0 174888 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 177520 0 177576 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 180208 0 180264 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 107632 0 107688 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 182896 0 182952 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 185584 0 185640 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 188272 0 188328 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 190960 0 191016 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 193648 0 193704 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 196336 0 196392 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 199024 0 199080 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 201712 0 201768 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 204400 0 204456 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 207088 0 207144 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 110320 0 110376 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 209776 0 209832 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 212464 0 212520 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 215152 0 215208 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 217840 0 217896 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 220528 0 220584 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 223216 0 223272 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 225904 0 225960 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 228592 0 228648 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 231280 0 231336 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 233968 0 234024 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 113008 0 113064 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 236656 0 236712 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 239344 0 239400 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 242032 0 242088 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 244720 0 244776 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 247408 0 247464 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 250096 0 250152 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 252784 0 252840 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 255472 0 255528 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 258160 0 258216 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 260848 0 260904 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 115696 0 115752 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 263536 0 263592 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 266224 0 266280 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 268912 0 268968 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 271600 0 271656 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 118384 0 118440 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 121072 0 121128 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 123760 0 123816 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 126448 0 126504 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal2 s 132496 175600 132552 176000 6 line_a_buf_b_a[0]
port 244 nsew signal output
rlabel metal2 s 132608 175600 132664 176000 6 line_a_buf_b_a[1]
port 245 nsew signal output
rlabel metal2 s 132720 175600 132776 176000 6 line_a_buf_b_a[2]
port 246 nsew signal output
rlabel metal2 s 127344 175600 127400 176000 6 line_a_buf_b_a[3]
port 247 nsew signal output
rlabel metal2 s 127456 175600 127512 176000 6 line_a_buf_b_a[4]
port 248 nsew signal output
rlabel metal2 s 127568 175600 127624 176000 6 line_a_buf_b_a[5]
port 249 nsew signal output
rlabel metal2 s 127680 175600 127736 176000 6 line_a_buf_b_a[6]
port 250 nsew signal output
rlabel metal2 s 132832 175600 132888 176000 6 line_a_buf_b_a[7]
port 251 nsew signal output
rlabel metal2 s 127792 175600 127848 176000 6 line_a_buf_b_cen
port 252 nsew signal output
rlabel metal2 s 132944 175600 133000 176000 6 line_a_buf_b_clk
port 253 nsew signal output
rlabel metal2 s 138768 175600 138824 176000 6 line_a_buf_b_d[0]
port 254 nsew signal output
rlabel metal2 s 137200 175600 137256 176000 6 line_a_buf_b_d[1]
port 255 nsew signal output
rlabel metal2 s 136864 175600 136920 176000 6 line_a_buf_b_d[2]
port 256 nsew signal output
rlabel metal2 s 134176 175600 134232 176000 6 line_a_buf_b_d[3]
port 257 nsew signal output
rlabel metal2 s 127232 175600 127288 176000 6 line_a_buf_b_d[4]
port 258 nsew signal output
rlabel metal2 s 124544 175600 124600 176000 6 line_a_buf_b_d[5]
port 259 nsew signal output
rlabel metal2 s 124208 175600 124264 176000 6 line_a_buf_b_d[6]
port 260 nsew signal output
rlabel metal2 s 122080 175600 122136 176000 6 line_a_buf_b_d[7]
port 261 nsew signal output
rlabel metal2 s 130704 175600 130760 176000 6 line_a_buf_b_gwen
port 262 nsew signal output
rlabel metal2 s 138544 175600 138600 176000 6 line_a_buf_b_q[0]
port 263 nsew signal input
rlabel metal2 s 137312 175600 137368 176000 6 line_a_buf_b_q[1]
port 264 nsew signal input
rlabel metal2 s 136752 175600 136808 176000 6 line_a_buf_b_q[2]
port 265 nsew signal input
rlabel metal2 s 134400 175600 134456 176000 6 line_a_buf_b_q[3]
port 266 nsew signal input
rlabel metal2 s 127008 175600 127064 176000 6 line_a_buf_b_q[4]
port 267 nsew signal input
rlabel metal2 s 124656 175600 124712 176000 6 line_a_buf_b_q[5]
port 268 nsew signal input
rlabel metal2 s 124096 175600 124152 176000 6 line_a_buf_b_q[6]
port 269 nsew signal input
rlabel metal2 s 122304 175600 122360 176000 6 line_a_buf_b_q[7]
port 270 nsew signal input
rlabel metal2 s 138656 175600 138712 176000 6 line_a_buf_b_wen[0]
port 271 nsew signal output
rlabel metal2 s 137088 175600 137144 176000 6 line_a_buf_b_wen[1]
port 272 nsew signal output
rlabel metal2 s 136976 175600 137032 176000 6 line_a_buf_b_wen[2]
port 273 nsew signal output
rlabel metal2 s 134288 175600 134344 176000 6 line_a_buf_b_wen[3]
port 274 nsew signal output
rlabel metal2 s 127120 175600 127176 176000 6 line_a_buf_b_wen[4]
port 275 nsew signal output
rlabel metal2 s 124432 175600 124488 176000 6 line_a_buf_b_wen[5]
port 276 nsew signal output
rlabel metal2 s 124320 175600 124376 176000 6 line_a_buf_b_wen[6]
port 277 nsew signal output
rlabel metal2 s 122192 175600 122248 176000 6 line_a_buf_b_wen[7]
port 278 nsew signal output
rlabel metal2 s 95536 175600 95592 176000 6 line_a_buf_d_a[0]
port 279 nsew signal output
rlabel metal2 s 95648 175600 95704 176000 6 line_a_buf_d_a[1]
port 280 nsew signal output
rlabel metal2 s 95760 175600 95816 176000 6 line_a_buf_d_a[2]
port 281 nsew signal output
rlabel metal2 s 90384 175600 90440 176000 6 line_a_buf_d_a[3]
port 282 nsew signal output
rlabel metal2 s 90496 175600 90552 176000 6 line_a_buf_d_a[4]
port 283 nsew signal output
rlabel metal2 s 90608 175600 90664 176000 6 line_a_buf_d_a[5]
port 284 nsew signal output
rlabel metal2 s 90720 175600 90776 176000 6 line_a_buf_d_a[6]
port 285 nsew signal output
rlabel metal2 s 95872 175600 95928 176000 6 line_a_buf_d_a[7]
port 286 nsew signal output
rlabel metal2 s 90832 175600 90888 176000 6 line_a_buf_d_cen
port 287 nsew signal output
rlabel metal2 s 95984 175600 96040 176000 6 line_a_buf_d_clk
port 288 nsew signal output
rlabel metal2 s 101808 175600 101864 176000 6 line_a_buf_d_d[0]
port 289 nsew signal output
rlabel metal2 s 100240 175600 100296 176000 6 line_a_buf_d_d[1]
port 290 nsew signal output
rlabel metal2 s 99904 175600 99960 176000 6 line_a_buf_d_d[2]
port 291 nsew signal output
rlabel metal2 s 97216 175600 97272 176000 6 line_a_buf_d_d[3]
port 292 nsew signal output
rlabel metal2 s 90272 175600 90328 176000 6 line_a_buf_d_d[4]
port 293 nsew signal output
rlabel metal2 s 87584 175600 87640 176000 6 line_a_buf_d_d[5]
port 294 nsew signal output
rlabel metal2 s 87248 175600 87304 176000 6 line_a_buf_d_d[6]
port 295 nsew signal output
rlabel metal2 s 85120 175600 85176 176000 6 line_a_buf_d_d[7]
port 296 nsew signal output
rlabel metal2 s 93744 175600 93800 176000 6 line_a_buf_d_gwen
port 297 nsew signal output
rlabel metal2 s 101584 175600 101640 176000 6 line_a_buf_d_q[0]
port 298 nsew signal input
rlabel metal2 s 100352 175600 100408 176000 6 line_a_buf_d_q[1]
port 299 nsew signal input
rlabel metal2 s 99792 175600 99848 176000 6 line_a_buf_d_q[2]
port 300 nsew signal input
rlabel metal2 s 97440 175600 97496 176000 6 line_a_buf_d_q[3]
port 301 nsew signal input
rlabel metal2 s 90048 175600 90104 176000 6 line_a_buf_d_q[4]
port 302 nsew signal input
rlabel metal2 s 87696 175600 87752 176000 6 line_a_buf_d_q[5]
port 303 nsew signal input
rlabel metal2 s 87136 175600 87192 176000 6 line_a_buf_d_q[6]
port 304 nsew signal input
rlabel metal2 s 85344 175600 85400 176000 6 line_a_buf_d_q[7]
port 305 nsew signal input
rlabel metal2 s 101696 175600 101752 176000 6 line_a_buf_d_wen[0]
port 306 nsew signal output
rlabel metal2 s 100128 175600 100184 176000 6 line_a_buf_d_wen[1]
port 307 nsew signal output
rlabel metal2 s 100016 175600 100072 176000 6 line_a_buf_d_wen[2]
port 308 nsew signal output
rlabel metal2 s 97328 175600 97384 176000 6 line_a_buf_d_wen[3]
port 309 nsew signal output
rlabel metal2 s 90160 175600 90216 176000 6 line_a_buf_d_wen[4]
port 310 nsew signal output
rlabel metal2 s 87472 175600 87528 176000 6 line_a_buf_d_wen[5]
port 311 nsew signal output
rlabel metal2 s 87360 175600 87416 176000 6 line_a_buf_d_wen[6]
port 312 nsew signal output
rlabel metal2 s 85232 175600 85288 176000 6 line_a_buf_d_wen[7]
port 313 nsew signal output
rlabel metal2 s 169456 175600 169512 176000 6 line_a_buf_g_a[0]
port 314 nsew signal output
rlabel metal2 s 169568 175600 169624 176000 6 line_a_buf_g_a[1]
port 315 nsew signal output
rlabel metal2 s 169680 175600 169736 176000 6 line_a_buf_g_a[2]
port 316 nsew signal output
rlabel metal2 s 164304 175600 164360 176000 6 line_a_buf_g_a[3]
port 317 nsew signal output
rlabel metal2 s 164416 175600 164472 176000 6 line_a_buf_g_a[4]
port 318 nsew signal output
rlabel metal2 s 164528 175600 164584 176000 6 line_a_buf_g_a[5]
port 319 nsew signal output
rlabel metal2 s 164640 175600 164696 176000 6 line_a_buf_g_a[6]
port 320 nsew signal output
rlabel metal2 s 169792 175600 169848 176000 6 line_a_buf_g_a[7]
port 321 nsew signal output
rlabel metal2 s 164752 175600 164808 176000 6 line_a_buf_g_cen
port 322 nsew signal output
rlabel metal2 s 169904 175600 169960 176000 6 line_a_buf_g_clk
port 323 nsew signal output
rlabel metal2 s 175728 175600 175784 176000 6 line_a_buf_g_d[0]
port 324 nsew signal output
rlabel metal2 s 174160 175600 174216 176000 6 line_a_buf_g_d[1]
port 325 nsew signal output
rlabel metal2 s 173824 175600 173880 176000 6 line_a_buf_g_d[2]
port 326 nsew signal output
rlabel metal2 s 171136 175600 171192 176000 6 line_a_buf_g_d[3]
port 327 nsew signal output
rlabel metal2 s 164192 175600 164248 176000 6 line_a_buf_g_d[4]
port 328 nsew signal output
rlabel metal2 s 161504 175600 161560 176000 6 line_a_buf_g_d[5]
port 329 nsew signal output
rlabel metal2 s 161168 175600 161224 176000 6 line_a_buf_g_d[6]
port 330 nsew signal output
rlabel metal2 s 159040 175600 159096 176000 6 line_a_buf_g_d[7]
port 331 nsew signal output
rlabel metal2 s 167664 175600 167720 176000 6 line_a_buf_g_gwen
port 332 nsew signal output
rlabel metal2 s 175504 175600 175560 176000 6 line_a_buf_g_q[0]
port 333 nsew signal input
rlabel metal2 s 174272 175600 174328 176000 6 line_a_buf_g_q[1]
port 334 nsew signal input
rlabel metal2 s 173712 175600 173768 176000 6 line_a_buf_g_q[2]
port 335 nsew signal input
rlabel metal2 s 171360 175600 171416 176000 6 line_a_buf_g_q[3]
port 336 nsew signal input
rlabel metal2 s 163968 175600 164024 176000 6 line_a_buf_g_q[4]
port 337 nsew signal input
rlabel metal2 s 161616 175600 161672 176000 6 line_a_buf_g_q[5]
port 338 nsew signal input
rlabel metal2 s 161056 175600 161112 176000 6 line_a_buf_g_q[6]
port 339 nsew signal input
rlabel metal2 s 159264 175600 159320 176000 6 line_a_buf_g_q[7]
port 340 nsew signal input
rlabel metal2 s 175616 175600 175672 176000 6 line_a_buf_g_wen[0]
port 341 nsew signal output
rlabel metal2 s 174048 175600 174104 176000 6 line_a_buf_g_wen[1]
port 342 nsew signal output
rlabel metal2 s 173936 175600 173992 176000 6 line_a_buf_g_wen[2]
port 343 nsew signal output
rlabel metal2 s 171248 175600 171304 176000 6 line_a_buf_g_wen[3]
port 344 nsew signal output
rlabel metal2 s 164080 175600 164136 176000 6 line_a_buf_g_wen[4]
port 345 nsew signal output
rlabel metal2 s 161392 175600 161448 176000 6 line_a_buf_g_wen[5]
port 346 nsew signal output
rlabel metal2 s 161280 175600 161336 176000 6 line_a_buf_g_wen[6]
port 347 nsew signal output
rlabel metal2 s 159152 175600 159208 176000 6 line_a_buf_g_wen[7]
port 348 nsew signal output
rlabel metal2 s 206416 175600 206472 176000 6 line_a_buf_r_a[0]
port 349 nsew signal output
rlabel metal2 s 206528 175600 206584 176000 6 line_a_buf_r_a[1]
port 350 nsew signal output
rlabel metal2 s 206640 175600 206696 176000 6 line_a_buf_r_a[2]
port 351 nsew signal output
rlabel metal2 s 201264 175600 201320 176000 6 line_a_buf_r_a[3]
port 352 nsew signal output
rlabel metal2 s 201376 175600 201432 176000 6 line_a_buf_r_a[4]
port 353 nsew signal output
rlabel metal2 s 201488 175600 201544 176000 6 line_a_buf_r_a[5]
port 354 nsew signal output
rlabel metal2 s 201600 175600 201656 176000 6 line_a_buf_r_a[6]
port 355 nsew signal output
rlabel metal2 s 206752 175600 206808 176000 6 line_a_buf_r_a[7]
port 356 nsew signal output
rlabel metal2 s 201712 175600 201768 176000 6 line_a_buf_r_cen
port 357 nsew signal output
rlabel metal2 s 206864 175600 206920 176000 6 line_a_buf_r_clk
port 358 nsew signal output
rlabel metal2 s 212688 175600 212744 176000 6 line_a_buf_r_d[0]
port 359 nsew signal output
rlabel metal2 s 211120 175600 211176 176000 6 line_a_buf_r_d[1]
port 360 nsew signal output
rlabel metal2 s 210784 175600 210840 176000 6 line_a_buf_r_d[2]
port 361 nsew signal output
rlabel metal2 s 208096 175600 208152 176000 6 line_a_buf_r_d[3]
port 362 nsew signal output
rlabel metal2 s 201152 175600 201208 176000 6 line_a_buf_r_d[4]
port 363 nsew signal output
rlabel metal2 s 198464 175600 198520 176000 6 line_a_buf_r_d[5]
port 364 nsew signal output
rlabel metal2 s 198128 175600 198184 176000 6 line_a_buf_r_d[6]
port 365 nsew signal output
rlabel metal2 s 196000 175600 196056 176000 6 line_a_buf_r_d[7]
port 366 nsew signal output
rlabel metal2 s 204624 175600 204680 176000 6 line_a_buf_r_gwen
port 367 nsew signal output
rlabel metal2 s 212464 175600 212520 176000 6 line_a_buf_r_q[0]
port 368 nsew signal input
rlabel metal2 s 211232 175600 211288 176000 6 line_a_buf_r_q[1]
port 369 nsew signal input
rlabel metal2 s 210672 175600 210728 176000 6 line_a_buf_r_q[2]
port 370 nsew signal input
rlabel metal2 s 208320 175600 208376 176000 6 line_a_buf_r_q[3]
port 371 nsew signal input
rlabel metal2 s 200928 175600 200984 176000 6 line_a_buf_r_q[4]
port 372 nsew signal input
rlabel metal2 s 198576 175600 198632 176000 6 line_a_buf_r_q[5]
port 373 nsew signal input
rlabel metal2 s 198016 175600 198072 176000 6 line_a_buf_r_q[6]
port 374 nsew signal input
rlabel metal2 s 196224 175600 196280 176000 6 line_a_buf_r_q[7]
port 375 nsew signal input
rlabel metal2 s 212576 175600 212632 176000 6 line_a_buf_r_wen[0]
port 376 nsew signal output
rlabel metal2 s 211008 175600 211064 176000 6 line_a_buf_r_wen[1]
port 377 nsew signal output
rlabel metal2 s 210896 175600 210952 176000 6 line_a_buf_r_wen[2]
port 378 nsew signal output
rlabel metal2 s 208208 175600 208264 176000 6 line_a_buf_r_wen[3]
port 379 nsew signal output
rlabel metal2 s 201040 175600 201096 176000 6 line_a_buf_r_wen[4]
port 380 nsew signal output
rlabel metal2 s 198352 175600 198408 176000 6 line_a_buf_r_wen[5]
port 381 nsew signal output
rlabel metal2 s 198240 175600 198296 176000 6 line_a_buf_r_wen[6]
port 382 nsew signal output
rlabel metal2 s 196112 175600 196168 176000 6 line_a_buf_r_wen[7]
port 383 nsew signal output
rlabel metal2 s 114016 175600 114072 176000 6 line_b_buf_b_a[0]
port 384 nsew signal output
rlabel metal2 s 114128 175600 114184 176000 6 line_b_buf_b_a[1]
port 385 nsew signal output
rlabel metal2 s 114240 175600 114296 176000 6 line_b_buf_b_a[2]
port 386 nsew signal output
rlabel metal2 s 108864 175600 108920 176000 6 line_b_buf_b_a[3]
port 387 nsew signal output
rlabel metal2 s 108976 175600 109032 176000 6 line_b_buf_b_a[4]
port 388 nsew signal output
rlabel metal2 s 109088 175600 109144 176000 6 line_b_buf_b_a[5]
port 389 nsew signal output
rlabel metal2 s 109200 175600 109256 176000 6 line_b_buf_b_a[6]
port 390 nsew signal output
rlabel metal2 s 114352 175600 114408 176000 6 line_b_buf_b_a[7]
port 391 nsew signal output
rlabel metal2 s 109312 175600 109368 176000 6 line_b_buf_b_cen
port 392 nsew signal output
rlabel metal2 s 114464 175600 114520 176000 6 line_b_buf_b_clk
port 393 nsew signal output
rlabel metal2 s 120288 175600 120344 176000 6 line_b_buf_b_d[0]
port 394 nsew signal output
rlabel metal2 s 118720 175600 118776 176000 6 line_b_buf_b_d[1]
port 395 nsew signal output
rlabel metal2 s 118384 175600 118440 176000 6 line_b_buf_b_d[2]
port 396 nsew signal output
rlabel metal2 s 115696 175600 115752 176000 6 line_b_buf_b_d[3]
port 397 nsew signal output
rlabel metal2 s 108752 175600 108808 176000 6 line_b_buf_b_d[4]
port 398 nsew signal output
rlabel metal2 s 106064 175600 106120 176000 6 line_b_buf_b_d[5]
port 399 nsew signal output
rlabel metal2 s 105728 175600 105784 176000 6 line_b_buf_b_d[6]
port 400 nsew signal output
rlabel metal2 s 103600 175600 103656 176000 6 line_b_buf_b_d[7]
port 401 nsew signal output
rlabel metal2 s 112224 175600 112280 176000 6 line_b_buf_b_gwen
port 402 nsew signal output
rlabel metal2 s 120064 175600 120120 176000 6 line_b_buf_b_q[0]
port 403 nsew signal input
rlabel metal2 s 118832 175600 118888 176000 6 line_b_buf_b_q[1]
port 404 nsew signal input
rlabel metal2 s 118272 175600 118328 176000 6 line_b_buf_b_q[2]
port 405 nsew signal input
rlabel metal2 s 115920 175600 115976 176000 6 line_b_buf_b_q[3]
port 406 nsew signal input
rlabel metal2 s 108528 175600 108584 176000 6 line_b_buf_b_q[4]
port 407 nsew signal input
rlabel metal2 s 106176 175600 106232 176000 6 line_b_buf_b_q[5]
port 408 nsew signal input
rlabel metal2 s 105616 175600 105672 176000 6 line_b_buf_b_q[6]
port 409 nsew signal input
rlabel metal2 s 103824 175600 103880 176000 6 line_b_buf_b_q[7]
port 410 nsew signal input
rlabel metal2 s 120176 175600 120232 176000 6 line_b_buf_b_wen[0]
port 411 nsew signal output
rlabel metal2 s 118608 175600 118664 176000 6 line_b_buf_b_wen[1]
port 412 nsew signal output
rlabel metal2 s 118496 175600 118552 176000 6 line_b_buf_b_wen[2]
port 413 nsew signal output
rlabel metal2 s 115808 175600 115864 176000 6 line_b_buf_b_wen[3]
port 414 nsew signal output
rlabel metal2 s 108640 175600 108696 176000 6 line_b_buf_b_wen[4]
port 415 nsew signal output
rlabel metal2 s 105952 175600 106008 176000 6 line_b_buf_b_wen[5]
port 416 nsew signal output
rlabel metal2 s 105840 175600 105896 176000 6 line_b_buf_b_wen[6]
port 417 nsew signal output
rlabel metal2 s 103712 175600 103768 176000 6 line_b_buf_b_wen[7]
port 418 nsew signal output
rlabel metal2 s 77056 175600 77112 176000 6 line_b_buf_d_a[0]
port 419 nsew signal output
rlabel metal2 s 77168 175600 77224 176000 6 line_b_buf_d_a[1]
port 420 nsew signal output
rlabel metal2 s 77280 175600 77336 176000 6 line_b_buf_d_a[2]
port 421 nsew signal output
rlabel metal2 s 71904 175600 71960 176000 6 line_b_buf_d_a[3]
port 422 nsew signal output
rlabel metal2 s 72016 175600 72072 176000 6 line_b_buf_d_a[4]
port 423 nsew signal output
rlabel metal2 s 72128 175600 72184 176000 6 line_b_buf_d_a[5]
port 424 nsew signal output
rlabel metal2 s 72240 175600 72296 176000 6 line_b_buf_d_a[6]
port 425 nsew signal output
rlabel metal2 s 77392 175600 77448 176000 6 line_b_buf_d_a[7]
port 426 nsew signal output
rlabel metal2 s 72352 175600 72408 176000 6 line_b_buf_d_cen
port 427 nsew signal output
rlabel metal2 s 77504 175600 77560 176000 6 line_b_buf_d_clk
port 428 nsew signal output
rlabel metal2 s 83328 175600 83384 176000 6 line_b_buf_d_d[0]
port 429 nsew signal output
rlabel metal2 s 81760 175600 81816 176000 6 line_b_buf_d_d[1]
port 430 nsew signal output
rlabel metal2 s 81424 175600 81480 176000 6 line_b_buf_d_d[2]
port 431 nsew signal output
rlabel metal2 s 78736 175600 78792 176000 6 line_b_buf_d_d[3]
port 432 nsew signal output
rlabel metal2 s 71792 175600 71848 176000 6 line_b_buf_d_d[4]
port 433 nsew signal output
rlabel metal2 s 69104 175600 69160 176000 6 line_b_buf_d_d[5]
port 434 nsew signal output
rlabel metal2 s 68768 175600 68824 176000 6 line_b_buf_d_d[6]
port 435 nsew signal output
rlabel metal2 s 66640 175600 66696 176000 6 line_b_buf_d_d[7]
port 436 nsew signal output
rlabel metal2 s 75264 175600 75320 176000 6 line_b_buf_d_gwen
port 437 nsew signal output
rlabel metal2 s 83104 175600 83160 176000 6 line_b_buf_d_q[0]
port 438 nsew signal input
rlabel metal2 s 81872 175600 81928 176000 6 line_b_buf_d_q[1]
port 439 nsew signal input
rlabel metal2 s 81312 175600 81368 176000 6 line_b_buf_d_q[2]
port 440 nsew signal input
rlabel metal2 s 78960 175600 79016 176000 6 line_b_buf_d_q[3]
port 441 nsew signal input
rlabel metal2 s 71568 175600 71624 176000 6 line_b_buf_d_q[4]
port 442 nsew signal input
rlabel metal2 s 69216 175600 69272 176000 6 line_b_buf_d_q[5]
port 443 nsew signal input
rlabel metal2 s 68656 175600 68712 176000 6 line_b_buf_d_q[6]
port 444 nsew signal input
rlabel metal2 s 66864 175600 66920 176000 6 line_b_buf_d_q[7]
port 445 nsew signal input
rlabel metal2 s 83216 175600 83272 176000 6 line_b_buf_d_wen[0]
port 446 nsew signal output
rlabel metal2 s 81648 175600 81704 176000 6 line_b_buf_d_wen[1]
port 447 nsew signal output
rlabel metal2 s 81536 175600 81592 176000 6 line_b_buf_d_wen[2]
port 448 nsew signal output
rlabel metal2 s 78848 175600 78904 176000 6 line_b_buf_d_wen[3]
port 449 nsew signal output
rlabel metal2 s 71680 175600 71736 176000 6 line_b_buf_d_wen[4]
port 450 nsew signal output
rlabel metal2 s 68992 175600 69048 176000 6 line_b_buf_d_wen[5]
port 451 nsew signal output
rlabel metal2 s 68880 175600 68936 176000 6 line_b_buf_d_wen[6]
port 452 nsew signal output
rlabel metal2 s 66752 175600 66808 176000 6 line_b_buf_d_wen[7]
port 453 nsew signal output
rlabel metal2 s 150976 175600 151032 176000 6 line_b_buf_g_a[0]
port 454 nsew signal output
rlabel metal2 s 151088 175600 151144 176000 6 line_b_buf_g_a[1]
port 455 nsew signal output
rlabel metal2 s 151200 175600 151256 176000 6 line_b_buf_g_a[2]
port 456 nsew signal output
rlabel metal2 s 145824 175600 145880 176000 6 line_b_buf_g_a[3]
port 457 nsew signal output
rlabel metal2 s 145936 175600 145992 176000 6 line_b_buf_g_a[4]
port 458 nsew signal output
rlabel metal2 s 146048 175600 146104 176000 6 line_b_buf_g_a[5]
port 459 nsew signal output
rlabel metal2 s 146160 175600 146216 176000 6 line_b_buf_g_a[6]
port 460 nsew signal output
rlabel metal2 s 151312 175600 151368 176000 6 line_b_buf_g_a[7]
port 461 nsew signal output
rlabel metal2 s 146272 175600 146328 176000 6 line_b_buf_g_cen
port 462 nsew signal output
rlabel metal2 s 151424 175600 151480 176000 6 line_b_buf_g_clk
port 463 nsew signal output
rlabel metal2 s 157248 175600 157304 176000 6 line_b_buf_g_d[0]
port 464 nsew signal output
rlabel metal2 s 155680 175600 155736 176000 6 line_b_buf_g_d[1]
port 465 nsew signal output
rlabel metal2 s 155344 175600 155400 176000 6 line_b_buf_g_d[2]
port 466 nsew signal output
rlabel metal2 s 152656 175600 152712 176000 6 line_b_buf_g_d[3]
port 467 nsew signal output
rlabel metal2 s 145712 175600 145768 176000 6 line_b_buf_g_d[4]
port 468 nsew signal output
rlabel metal2 s 143024 175600 143080 176000 6 line_b_buf_g_d[5]
port 469 nsew signal output
rlabel metal2 s 142688 175600 142744 176000 6 line_b_buf_g_d[6]
port 470 nsew signal output
rlabel metal2 s 140560 175600 140616 176000 6 line_b_buf_g_d[7]
port 471 nsew signal output
rlabel metal2 s 149184 175600 149240 176000 6 line_b_buf_g_gwen
port 472 nsew signal output
rlabel metal2 s 157024 175600 157080 176000 6 line_b_buf_g_q[0]
port 473 nsew signal input
rlabel metal2 s 155792 175600 155848 176000 6 line_b_buf_g_q[1]
port 474 nsew signal input
rlabel metal2 s 155232 175600 155288 176000 6 line_b_buf_g_q[2]
port 475 nsew signal input
rlabel metal2 s 152880 175600 152936 176000 6 line_b_buf_g_q[3]
port 476 nsew signal input
rlabel metal2 s 145488 175600 145544 176000 6 line_b_buf_g_q[4]
port 477 nsew signal input
rlabel metal2 s 143136 175600 143192 176000 6 line_b_buf_g_q[5]
port 478 nsew signal input
rlabel metal2 s 142576 175600 142632 176000 6 line_b_buf_g_q[6]
port 479 nsew signal input
rlabel metal2 s 140784 175600 140840 176000 6 line_b_buf_g_q[7]
port 480 nsew signal input
rlabel metal2 s 157136 175600 157192 176000 6 line_b_buf_g_wen[0]
port 481 nsew signal output
rlabel metal2 s 155568 175600 155624 176000 6 line_b_buf_g_wen[1]
port 482 nsew signal output
rlabel metal2 s 155456 175600 155512 176000 6 line_b_buf_g_wen[2]
port 483 nsew signal output
rlabel metal2 s 152768 175600 152824 176000 6 line_b_buf_g_wen[3]
port 484 nsew signal output
rlabel metal2 s 145600 175600 145656 176000 6 line_b_buf_g_wen[4]
port 485 nsew signal output
rlabel metal2 s 142912 175600 142968 176000 6 line_b_buf_g_wen[5]
port 486 nsew signal output
rlabel metal2 s 142800 175600 142856 176000 6 line_b_buf_g_wen[6]
port 487 nsew signal output
rlabel metal2 s 140672 175600 140728 176000 6 line_b_buf_g_wen[7]
port 488 nsew signal output
rlabel metal2 s 187936 175600 187992 176000 6 line_b_buf_r_a[0]
port 489 nsew signal output
rlabel metal2 s 188048 175600 188104 176000 6 line_b_buf_r_a[1]
port 490 nsew signal output
rlabel metal2 s 188160 175600 188216 176000 6 line_b_buf_r_a[2]
port 491 nsew signal output
rlabel metal2 s 182784 175600 182840 176000 6 line_b_buf_r_a[3]
port 492 nsew signal output
rlabel metal2 s 182896 175600 182952 176000 6 line_b_buf_r_a[4]
port 493 nsew signal output
rlabel metal2 s 183008 175600 183064 176000 6 line_b_buf_r_a[5]
port 494 nsew signal output
rlabel metal2 s 183120 175600 183176 176000 6 line_b_buf_r_a[6]
port 495 nsew signal output
rlabel metal2 s 188272 175600 188328 176000 6 line_b_buf_r_a[7]
port 496 nsew signal output
rlabel metal2 s 183232 175600 183288 176000 6 line_b_buf_r_cen
port 497 nsew signal output
rlabel metal2 s 188384 175600 188440 176000 6 line_b_buf_r_clk
port 498 nsew signal output
rlabel metal2 s 194208 175600 194264 176000 6 line_b_buf_r_d[0]
port 499 nsew signal output
rlabel metal2 s 192640 175600 192696 176000 6 line_b_buf_r_d[1]
port 500 nsew signal output
rlabel metal2 s 192304 175600 192360 176000 6 line_b_buf_r_d[2]
port 501 nsew signal output
rlabel metal2 s 189616 175600 189672 176000 6 line_b_buf_r_d[3]
port 502 nsew signal output
rlabel metal2 s 182672 175600 182728 176000 6 line_b_buf_r_d[4]
port 503 nsew signal output
rlabel metal2 s 179984 175600 180040 176000 6 line_b_buf_r_d[5]
port 504 nsew signal output
rlabel metal2 s 179648 175600 179704 176000 6 line_b_buf_r_d[6]
port 505 nsew signal output
rlabel metal2 s 177520 175600 177576 176000 6 line_b_buf_r_d[7]
port 506 nsew signal output
rlabel metal2 s 186144 175600 186200 176000 6 line_b_buf_r_gwen
port 507 nsew signal output
rlabel metal2 s 193984 175600 194040 176000 6 line_b_buf_r_q[0]
port 508 nsew signal input
rlabel metal2 s 192752 175600 192808 176000 6 line_b_buf_r_q[1]
port 509 nsew signal input
rlabel metal2 s 192192 175600 192248 176000 6 line_b_buf_r_q[2]
port 510 nsew signal input
rlabel metal2 s 189840 175600 189896 176000 6 line_b_buf_r_q[3]
port 511 nsew signal input
rlabel metal2 s 182448 175600 182504 176000 6 line_b_buf_r_q[4]
port 512 nsew signal input
rlabel metal2 s 180096 175600 180152 176000 6 line_b_buf_r_q[5]
port 513 nsew signal input
rlabel metal2 s 179536 175600 179592 176000 6 line_b_buf_r_q[6]
port 514 nsew signal input
rlabel metal2 s 177744 175600 177800 176000 6 line_b_buf_r_q[7]
port 515 nsew signal input
rlabel metal2 s 194096 175600 194152 176000 6 line_b_buf_r_wen[0]
port 516 nsew signal output
rlabel metal2 s 192528 175600 192584 176000 6 line_b_buf_r_wen[1]
port 517 nsew signal output
rlabel metal2 s 192416 175600 192472 176000 6 line_b_buf_r_wen[2]
port 518 nsew signal output
rlabel metal2 s 189728 175600 189784 176000 6 line_b_buf_r_wen[3]
port 519 nsew signal output
rlabel metal2 s 182560 175600 182616 176000 6 line_b_buf_r_wen[4]
port 520 nsew signal output
rlabel metal2 s 179872 175600 179928 176000 6 line_b_buf_r_wen[5]
port 521 nsew signal output
rlabel metal2 s 179760 175600 179816 176000 6 line_b_buf_r_wen[6]
port 522 nsew signal output
rlabel metal2 s 177632 175600 177688 176000 6 line_b_buf_r_wen[7]
port 523 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 524 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 525 nsew ground bidirectional
rlabel metal2 s 5488 0 5544 400 6 wb_clk_i
port 526 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 wb_rst_i
port 527 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 wbs_ack_o
port 528 nsew signal output
rlabel metal2 s 10864 0 10920 400 6 wbs_adr_i[0]
port 529 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 wbs_adr_i[10]
port 530 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 wbs_adr_i[11]
port 531 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 wbs_adr_i[12]
port 532 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 wbs_adr_i[13]
port 533 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 wbs_adr_i[14]
port 534 nsew signal input
rlabel metal2 s 54768 0 54824 400 6 wbs_adr_i[15]
port 535 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 wbs_adr_i[16]
port 536 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 wbs_adr_i[17]
port 537 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 wbs_adr_i[18]
port 538 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 wbs_adr_i[19]
port 539 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_adr_i[1]
port 540 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 wbs_adr_i[20]
port 541 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 wbs_adr_i[21]
port 542 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 wbs_adr_i[22]
port 543 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 wbs_adr_i[23]
port 544 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 wbs_adr_i[24]
port 545 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 wbs_adr_i[25]
port 546 nsew signal input
rlabel metal2 s 84336 0 84392 400 6 wbs_adr_i[26]
port 547 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 wbs_adr_i[27]
port 548 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 wbs_adr_i[28]
port 549 nsew signal input
rlabel metal2 s 92400 0 92456 400 6 wbs_adr_i[29]
port 550 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_adr_i[2]
port 551 nsew signal input
rlabel metal2 s 95088 0 95144 400 6 wbs_adr_i[30]
port 552 nsew signal input
rlabel metal2 s 97776 0 97832 400 6 wbs_adr_i[31]
port 553 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_adr_i[3]
port 554 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 wbs_adr_i[4]
port 555 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 wbs_adr_i[5]
port 556 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 wbs_adr_i[6]
port 557 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 wbs_adr_i[7]
port 558 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 wbs_adr_i[8]
port 559 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 wbs_adr_i[9]
port 560 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_cyc_i
port 561 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_dat_i[0]
port 562 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 wbs_dat_i[10]
port 563 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 wbs_dat_i[11]
port 564 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 wbs_dat_i[12]
port 565 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 wbs_dat_i[13]
port 566 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 wbs_dat_i[14]
port 567 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 wbs_dat_i[15]
port 568 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 wbs_dat_i[16]
port 569 nsew signal input
rlabel metal2 s 61040 0 61096 400 6 wbs_dat_i[17]
port 570 nsew signal input
rlabel metal2 s 63728 0 63784 400 6 wbs_dat_i[18]
port 571 nsew signal input
rlabel metal2 s 66416 0 66472 400 6 wbs_dat_i[19]
port 572 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_dat_i[1]
port 573 nsew signal input
rlabel metal2 s 69104 0 69160 400 6 wbs_dat_i[20]
port 574 nsew signal input
rlabel metal2 s 71792 0 71848 400 6 wbs_dat_i[21]
port 575 nsew signal input
rlabel metal2 s 74480 0 74536 400 6 wbs_dat_i[22]
port 576 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 wbs_dat_i[23]
port 577 nsew signal input
rlabel metal2 s 79856 0 79912 400 6 wbs_dat_i[24]
port 578 nsew signal input
rlabel metal2 s 82544 0 82600 400 6 wbs_dat_i[25]
port 579 nsew signal input
rlabel metal2 s 85232 0 85288 400 6 wbs_dat_i[26]
port 580 nsew signal input
rlabel metal2 s 87920 0 87976 400 6 wbs_dat_i[27]
port 581 nsew signal input
rlabel metal2 s 90608 0 90664 400 6 wbs_dat_i[28]
port 582 nsew signal input
rlabel metal2 s 93296 0 93352 400 6 wbs_dat_i[29]
port 583 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_i[2]
port 584 nsew signal input
rlabel metal2 s 95984 0 96040 400 6 wbs_dat_i[30]
port 585 nsew signal input
rlabel metal2 s 98672 0 98728 400 6 wbs_dat_i[31]
port 586 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 wbs_dat_i[3]
port 587 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_i[4]
port 588 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[5]
port 589 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 wbs_dat_i[6]
port 590 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 wbs_dat_i[7]
port 591 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 wbs_dat_i[8]
port 592 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_i[9]
port 593 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_o[0]
port 594 nsew signal output
rlabel metal2 s 43120 0 43176 400 6 wbs_dat_o[10]
port 595 nsew signal output
rlabel metal2 s 45808 0 45864 400 6 wbs_dat_o[11]
port 596 nsew signal output
rlabel metal2 s 48496 0 48552 400 6 wbs_dat_o[12]
port 597 nsew signal output
rlabel metal2 s 51184 0 51240 400 6 wbs_dat_o[13]
port 598 nsew signal output
rlabel metal2 s 53872 0 53928 400 6 wbs_dat_o[14]
port 599 nsew signal output
rlabel metal2 s 56560 0 56616 400 6 wbs_dat_o[15]
port 600 nsew signal output
rlabel metal2 s 59248 0 59304 400 6 wbs_dat_o[16]
port 601 nsew signal output
rlabel metal2 s 61936 0 61992 400 6 wbs_dat_o[17]
port 602 nsew signal output
rlabel metal2 s 64624 0 64680 400 6 wbs_dat_o[18]
port 603 nsew signal output
rlabel metal2 s 67312 0 67368 400 6 wbs_dat_o[19]
port 604 nsew signal output
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_o[1]
port 605 nsew signal output
rlabel metal2 s 70000 0 70056 400 6 wbs_dat_o[20]
port 606 nsew signal output
rlabel metal2 s 72688 0 72744 400 6 wbs_dat_o[21]
port 607 nsew signal output
rlabel metal2 s 75376 0 75432 400 6 wbs_dat_o[22]
port 608 nsew signal output
rlabel metal2 s 78064 0 78120 400 6 wbs_dat_o[23]
port 609 nsew signal output
rlabel metal2 s 80752 0 80808 400 6 wbs_dat_o[24]
port 610 nsew signal output
rlabel metal2 s 83440 0 83496 400 6 wbs_dat_o[25]
port 611 nsew signal output
rlabel metal2 s 86128 0 86184 400 6 wbs_dat_o[26]
port 612 nsew signal output
rlabel metal2 s 88816 0 88872 400 6 wbs_dat_o[27]
port 613 nsew signal output
rlabel metal2 s 91504 0 91560 400 6 wbs_dat_o[28]
port 614 nsew signal output
rlabel metal2 s 94192 0 94248 400 6 wbs_dat_o[29]
port 615 nsew signal output
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_o[2]
port 616 nsew signal output
rlabel metal2 s 96880 0 96936 400 6 wbs_dat_o[30]
port 617 nsew signal output
rlabel metal2 s 99568 0 99624 400 6 wbs_dat_o[31]
port 618 nsew signal output
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_o[3]
port 619 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 wbs_dat_o[4]
port 620 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 wbs_dat_o[5]
port 621 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 wbs_dat_o[6]
port 622 nsew signal output
rlabel metal2 s 35056 0 35112 400 6 wbs_dat_o[7]
port 623 nsew signal output
rlabel metal2 s 37744 0 37800 400 6 wbs_dat_o[8]
port 624 nsew signal output
rlabel metal2 s 40432 0 40488 400 6 wbs_dat_o[9]
port 625 nsew signal output
rlabel metal2 s 13552 0 13608 400 6 wbs_sel_i[0]
port 626 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_sel_i[1]
port 627 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_sel_i[2]
port 628 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_sel_i[3]
port 629 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_stb_i
port 630 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_we_i
port 631 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15246040
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/tjrpu/runs/23_11_17_19_04/results/signoff/tjrpu.magic.gds
string GDS_START 65072
<< end >>

