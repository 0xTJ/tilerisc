magic
tech gf180mcuD
magscale 1 10
timestamp 1700950315
<< metal1 >>
rect 16818 76974 16830 77026
rect 16882 77023 16894 77026
rect 17938 77023 17950 77026
rect 16882 76977 17950 77023
rect 16882 76974 16894 76977
rect 17938 76974 17950 76977
rect 18002 76974 18014 77026
rect 18610 76974 18622 77026
rect 18674 77023 18686 77026
rect 19170 77023 19182 77026
rect 18674 76977 19182 77023
rect 18674 76974 18686 76977
rect 19170 76974 19182 76977
rect 19234 76974 19246 77026
rect 20402 76974 20414 77026
rect 20466 77023 20478 77026
rect 21522 77023 21534 77026
rect 20466 76977 21534 77023
rect 20466 76974 20478 76977
rect 21522 76974 21534 76977
rect 21586 76974 21598 77026
rect 22194 76974 22206 77026
rect 22258 77023 22270 77026
rect 23090 77023 23102 77026
rect 22258 76977 23102 77023
rect 22258 76974 22270 76977
rect 23090 76974 23102 76977
rect 23154 76974 23166 77026
rect 25778 76974 25790 77026
rect 25842 77023 25854 77026
rect 26338 77023 26350 77026
rect 25842 76977 26350 77023
rect 25842 76974 25854 76977
rect 26338 76974 26350 76977
rect 26402 76974 26414 77026
rect 43698 76974 43710 77026
rect 43762 77023 43774 77026
rect 44258 77023 44270 77026
rect 43762 76977 44270 77023
rect 43762 76974 43774 76977
rect 44258 76974 44270 76977
rect 44322 77023 44334 77026
rect 44706 77023 44718 77026
rect 44322 76977 44718 77023
rect 44322 76974 44334 76977
rect 44706 76974 44718 76977
rect 44770 76974 44782 77026
rect 45490 76974 45502 77026
rect 45554 77023 45566 77026
rect 46050 77023 46062 77026
rect 45554 76977 46062 77023
rect 45554 76974 45566 76977
rect 46050 76974 46062 76977
rect 46114 77023 46126 77026
rect 46498 77023 46510 77026
rect 46114 76977 46510 77023
rect 46114 76974 46126 76977
rect 46498 76974 46510 76977
rect 46562 76974 46574 77026
rect 1344 76858 48608 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 48608 76858
rect 1344 76772 48608 76806
rect 10222 76690 10274 76702
rect 10222 76626 10274 76638
rect 11790 76690 11842 76702
rect 11790 76626 11842 76638
rect 21534 76690 21586 76702
rect 21534 76626 21586 76638
rect 30382 76690 30434 76702
rect 30382 76626 30434 76638
rect 32622 76690 32674 76702
rect 32622 76626 32674 76638
rect 37550 76690 37602 76702
rect 37550 76626 37602 76638
rect 42926 76690 42978 76702
rect 42926 76626 42978 76638
rect 44270 76690 44322 76702
rect 44270 76626 44322 76638
rect 44718 76690 44770 76702
rect 44718 76626 44770 76638
rect 46062 76690 46114 76702
rect 46062 76626 46114 76638
rect 46510 76690 46562 76702
rect 46510 76626 46562 76638
rect 48190 76690 48242 76702
rect 48190 76626 48242 76638
rect 36094 76578 36146 76590
rect 2482 76526 2494 76578
rect 2546 76526 2558 76578
rect 7858 76526 7870 76578
rect 7922 76526 7934 76578
rect 17938 76526 17950 76578
rect 18002 76526 18014 76578
rect 19170 76526 19182 76578
rect 19234 76526 19246 76578
rect 26338 76526 26350 76578
rect 26402 76526 26414 76578
rect 36094 76514 36146 76526
rect 41470 76578 41522 76590
rect 41470 76514 41522 76526
rect 13470 76466 13522 76478
rect 3266 76414 3278 76466
rect 3330 76414 3342 76466
rect 3714 76414 3726 76466
rect 3778 76414 3790 76466
rect 6962 76414 6974 76466
rect 7026 76414 7038 76466
rect 8754 76414 8766 76466
rect 8818 76414 8830 76466
rect 10882 76414 10894 76466
rect 10946 76414 10958 76466
rect 12450 76414 12462 76466
rect 12514 76414 12526 76466
rect 13470 76402 13522 76414
rect 15150 76466 15202 76478
rect 20750 76466 20802 76478
rect 28814 76466 28866 76478
rect 17042 76414 17054 76466
rect 17106 76414 17118 76466
rect 20066 76414 20078 76466
rect 20130 76414 20142 76466
rect 22418 76414 22430 76466
rect 22482 76414 22494 76466
rect 27234 76414 27246 76466
rect 27298 76414 27310 76466
rect 15150 76402 15202 76414
rect 20750 76402 20802 76414
rect 28814 76402 28866 76414
rect 31166 76466 31218 76478
rect 31166 76402 31218 76414
rect 33406 76466 33458 76478
rect 43710 76466 43762 76478
rect 35074 76414 35086 76466
rect 35138 76414 35150 76466
rect 36978 76414 36990 76466
rect 37042 76414 37054 76466
rect 38770 76414 38782 76466
rect 38834 76414 38846 76466
rect 40786 76414 40798 76466
rect 40850 76414 40862 76466
rect 42354 76414 42366 76466
rect 42418 76414 42430 76466
rect 33406 76402 33458 76414
rect 43710 76402 43762 76414
rect 22094 76354 22146 76366
rect 36542 76354 36594 76366
rect 4386 76302 4398 76354
rect 4450 76302 4462 76354
rect 6178 76302 6190 76354
rect 6242 76302 6254 76354
rect 13906 76302 13918 76354
rect 13970 76302 13982 76354
rect 15586 76302 15598 76354
rect 15650 76302 15662 76354
rect 23090 76302 23102 76354
rect 23154 76302 23166 76354
rect 29250 76302 29262 76354
rect 29314 76302 29326 76354
rect 22094 76290 22146 76302
rect 36542 76290 36594 76302
rect 38334 76354 38386 76366
rect 45502 76354 45554 76366
rect 42018 76302 42030 76354
rect 42082 76302 42094 76354
rect 38334 76290 38386 76302
rect 45502 76290 45554 76302
rect 34302 76242 34354 76254
rect 34302 76178 34354 76190
rect 40014 76242 40066 76254
rect 40014 76178 40066 76190
rect 1344 76074 48608 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 48608 76074
rect 1344 75988 48608 76022
rect 3614 75794 3666 75806
rect 3614 75730 3666 75742
rect 19070 75794 19122 75806
rect 39118 75794 39170 75806
rect 24434 75742 24446 75794
rect 24498 75742 24510 75794
rect 34738 75742 34750 75794
rect 34802 75742 34814 75794
rect 19070 75730 19122 75742
rect 39118 75730 39170 75742
rect 2606 75682 2658 75694
rect 2606 75618 2658 75630
rect 3166 75682 3218 75694
rect 3166 75618 3218 75630
rect 9102 75682 9154 75694
rect 9102 75618 9154 75630
rect 20526 75682 20578 75694
rect 29262 75682 29314 75694
rect 25442 75630 25454 75682
rect 25506 75630 25518 75682
rect 20526 75618 20578 75630
rect 29262 75618 29314 75630
rect 31502 75682 31554 75694
rect 31938 75630 31950 75682
rect 32002 75630 32014 75682
rect 31502 75618 31554 75630
rect 1710 75570 1762 75582
rect 1710 75506 1762 75518
rect 2270 75570 2322 75582
rect 2270 75506 2322 75518
rect 15934 75570 15986 75582
rect 15934 75506 15986 75518
rect 16270 75570 16322 75582
rect 48190 75570 48242 75582
rect 32610 75518 32622 75570
rect 32674 75518 32686 75570
rect 16270 75506 16322 75518
rect 48190 75506 48242 75518
rect 13694 75458 13746 75470
rect 13694 75394 13746 75406
rect 17054 75458 17106 75470
rect 17054 75394 17106 75406
rect 26014 75458 26066 75470
rect 26014 75394 26066 75406
rect 1344 75290 48608 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 48608 75290
rect 1344 75204 48608 75238
rect 33294 75122 33346 75134
rect 33294 75058 33346 75070
rect 33518 75122 33570 75134
rect 33518 75058 33570 75070
rect 5406 75010 5458 75022
rect 25230 75010 25282 75022
rect 4050 74958 4062 75010
rect 4114 74958 4126 75010
rect 6626 74958 6638 75010
rect 6690 74958 6702 75010
rect 14690 74958 14702 75010
rect 14754 74958 14766 75010
rect 5406 74946 5458 74958
rect 25230 74946 25282 74958
rect 23998 74898 24050 74910
rect 4834 74846 4846 74898
rect 4898 74846 4910 74898
rect 5842 74846 5854 74898
rect 5906 74846 5918 74898
rect 10658 74846 10670 74898
rect 10722 74846 10734 74898
rect 14018 74846 14030 74898
rect 14082 74846 14094 74898
rect 17378 74846 17390 74898
rect 17442 74846 17454 74898
rect 23538 74846 23550 74898
rect 23602 74846 23614 74898
rect 23998 74834 24050 74846
rect 24670 74898 24722 74910
rect 25442 74846 25454 74898
rect 25506 74846 25518 74898
rect 26002 74846 26014 74898
rect 26066 74846 26078 74898
rect 31938 74846 31950 74898
rect 32002 74846 32014 74898
rect 24670 74834 24722 74846
rect 9662 74786 9714 74798
rect 1922 74734 1934 74786
rect 1986 74734 1998 74786
rect 8754 74734 8766 74786
rect 8818 74734 8830 74786
rect 11330 74734 11342 74786
rect 11394 74734 11406 74786
rect 13458 74734 13470 74786
rect 13522 74734 13534 74786
rect 16818 74734 16830 74786
rect 16882 74734 16894 74786
rect 18162 74734 18174 74786
rect 18226 74734 18238 74786
rect 20290 74734 20302 74786
rect 20354 74734 20366 74786
rect 20626 74734 20638 74786
rect 20690 74734 20702 74786
rect 22754 74734 22766 74786
rect 22818 74734 22830 74786
rect 26674 74734 26686 74786
rect 26738 74734 26750 74786
rect 28802 74734 28814 74786
rect 28866 74734 28878 74786
rect 29138 74734 29150 74786
rect 29202 74734 29214 74786
rect 31266 74734 31278 74786
rect 31330 74734 31342 74786
rect 33954 74734 33966 74786
rect 34018 74734 34030 74786
rect 9662 74722 9714 74734
rect 1344 74506 48608 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 48608 74506
rect 1344 74420 48608 74454
rect 1822 74226 1874 74238
rect 20190 74226 20242 74238
rect 12002 74174 12014 74226
rect 12066 74174 12078 74226
rect 13458 74174 13470 74226
rect 13522 74174 13534 74226
rect 15586 74174 15598 74226
rect 15650 74174 15662 74226
rect 1822 74162 1874 74174
rect 20190 74162 20242 74174
rect 22318 74226 22370 74238
rect 22318 74162 22370 74174
rect 22766 74226 22818 74238
rect 23874 74174 23886 74226
rect 23938 74174 23950 74226
rect 26002 74174 26014 74226
rect 26066 74174 26078 74226
rect 32386 74174 32398 74226
rect 32450 74174 32462 74226
rect 22766 74162 22818 74174
rect 3938 74062 3950 74114
rect 4002 74062 4014 74114
rect 9090 74062 9102 74114
rect 9154 74062 9166 74114
rect 16370 74062 16382 74114
rect 16434 74062 16446 74114
rect 17602 74062 17614 74114
rect 17666 74062 17678 74114
rect 18162 74062 18174 74114
rect 18226 74062 18238 74114
rect 23202 74062 23214 74114
rect 23266 74062 23278 74114
rect 26562 74062 26574 74114
rect 26626 74062 26638 74114
rect 29586 74062 29598 74114
rect 29650 74062 29662 74114
rect 33282 74062 33294 74114
rect 33346 74062 33358 74114
rect 3390 74002 3442 74014
rect 3390 73938 3442 73950
rect 4734 74002 4786 74014
rect 4734 73938 4786 73950
rect 5742 74002 5794 74014
rect 12462 74002 12514 74014
rect 9874 73950 9886 74002
rect 9938 73950 9950 74002
rect 5742 73938 5794 73950
rect 12462 73938 12514 73950
rect 16830 74002 16882 74014
rect 19406 74002 19458 74014
rect 18834 73950 18846 74002
rect 18898 73950 18910 74002
rect 16830 73938 16882 73950
rect 19406 73938 19458 73950
rect 19742 74002 19794 74014
rect 19742 73938 19794 73950
rect 20750 74002 20802 74014
rect 20750 73938 20802 73950
rect 26350 74002 26402 74014
rect 26350 73938 26402 73950
rect 27246 74002 27298 74014
rect 27246 73938 27298 73950
rect 27582 74002 27634 74014
rect 27582 73938 27634 73950
rect 28254 74002 28306 74014
rect 28254 73938 28306 73950
rect 28590 74002 28642 74014
rect 33070 74002 33122 74014
rect 30258 73950 30270 74002
rect 30322 73950 30334 74002
rect 28590 73938 28642 73950
rect 33070 73938 33122 73950
rect 4174 73890 4226 73902
rect 4174 73826 4226 73838
rect 1344 73722 48608 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 48608 73722
rect 1344 73636 48608 73670
rect 10334 73554 10386 73566
rect 10334 73490 10386 73502
rect 23102 73554 23154 73566
rect 23102 73490 23154 73502
rect 27694 73554 27746 73566
rect 27694 73490 27746 73502
rect 29150 73554 29202 73566
rect 29150 73490 29202 73502
rect 30606 73554 30658 73566
rect 30606 73490 30658 73502
rect 9550 73442 9602 73454
rect 9550 73378 9602 73390
rect 25454 73442 25506 73454
rect 25454 73378 25506 73390
rect 48190 73442 48242 73454
rect 48190 73378 48242 73390
rect 1710 73330 1762 73342
rect 9886 73330 9938 73342
rect 4050 73278 4062 73330
rect 4114 73278 4126 73330
rect 1710 73266 1762 73278
rect 9886 73266 9938 73278
rect 10670 73330 10722 73342
rect 19182 73330 19234 73342
rect 28030 73330 28082 73342
rect 13794 73278 13806 73330
rect 13858 73278 13870 73330
rect 18610 73278 18622 73330
rect 18674 73278 18686 73330
rect 20290 73278 20302 73330
rect 20354 73278 20366 73330
rect 20626 73278 20638 73330
rect 20690 73278 20702 73330
rect 21970 73278 21982 73330
rect 22034 73278 22046 73330
rect 22418 73278 22430 73330
rect 22482 73278 22494 73330
rect 23874 73278 23886 73330
rect 23938 73278 23950 73330
rect 24322 73278 24334 73330
rect 24386 73278 24398 73330
rect 25666 73278 25678 73330
rect 25730 73278 25742 73330
rect 30818 73278 30830 73330
rect 30882 73278 30894 73330
rect 10670 73266 10722 73278
rect 19182 73266 19234 73278
rect 28030 73266 28082 73278
rect 2270 73218 2322 73230
rect 7422 73218 7474 73230
rect 4834 73166 4846 73218
rect 4898 73166 4910 73218
rect 6962 73166 6974 73218
rect 7026 73166 7038 73218
rect 2270 73154 2322 73166
rect 7422 73154 7474 73166
rect 9102 73218 9154 73230
rect 9102 73154 9154 73166
rect 11118 73218 11170 73230
rect 17950 73218 18002 73230
rect 14466 73166 14478 73218
rect 14530 73166 14542 73218
rect 16594 73166 16606 73218
rect 16658 73166 16670 73218
rect 11118 73154 11170 73166
rect 17950 73154 18002 73166
rect 19294 73218 19346 73230
rect 22654 73218 22706 73230
rect 21298 73166 21310 73218
rect 21362 73166 21374 73218
rect 19294 73154 19346 73166
rect 22654 73154 22706 73166
rect 23662 73218 23714 73230
rect 23662 73154 23714 73166
rect 26238 73218 26290 73230
rect 26238 73154 26290 73166
rect 26686 73218 26738 73230
rect 26686 73154 26738 73166
rect 28478 73218 28530 73230
rect 28478 73154 28530 73166
rect 1344 72938 48608 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 48608 72938
rect 1344 72852 48608 72886
rect 10658 72718 10670 72770
rect 10722 72767 10734 72770
rect 10994 72767 11006 72770
rect 10722 72721 11006 72767
rect 10722 72718 10734 72721
rect 10994 72718 11006 72721
rect 11058 72718 11070 72770
rect 1822 72658 1874 72670
rect 10894 72658 10946 72670
rect 8306 72606 8318 72658
rect 8370 72606 8382 72658
rect 10434 72606 10446 72658
rect 10498 72606 10510 72658
rect 1822 72594 1874 72606
rect 10894 72594 10946 72606
rect 17166 72658 17218 72670
rect 17166 72594 17218 72606
rect 18174 72658 18226 72670
rect 25678 72658 25730 72670
rect 18946 72606 18958 72658
rect 19010 72606 19022 72658
rect 20626 72606 20638 72658
rect 20690 72606 20702 72658
rect 22418 72606 22430 72658
rect 22482 72606 22494 72658
rect 18174 72594 18226 72606
rect 25678 72594 25730 72606
rect 30494 72658 30546 72670
rect 30494 72594 30546 72606
rect 33182 72658 33234 72670
rect 33182 72594 33234 72606
rect 31390 72546 31442 72558
rect 33070 72546 33122 72558
rect 5842 72494 5854 72546
rect 5906 72494 5918 72546
rect 7522 72494 7534 72546
rect 7586 72494 7598 72546
rect 18722 72494 18734 72546
rect 18786 72494 18798 72546
rect 20290 72494 20302 72546
rect 20354 72494 20366 72546
rect 22194 72494 22206 72546
rect 22258 72494 22270 72546
rect 23986 72494 23998 72546
rect 24050 72494 24062 72546
rect 24546 72494 24558 72546
rect 24610 72494 24622 72546
rect 31154 72494 31166 72546
rect 31218 72494 31230 72546
rect 32498 72494 32510 72546
rect 32562 72494 32574 72546
rect 31390 72482 31442 72494
rect 33070 72482 33122 72494
rect 33854 72546 33906 72558
rect 33854 72482 33906 72494
rect 34078 72546 34130 72558
rect 34078 72482 34130 72494
rect 5630 72434 5682 72446
rect 5630 72370 5682 72382
rect 6526 72434 6578 72446
rect 6526 72370 6578 72382
rect 19406 72434 19458 72446
rect 19406 72370 19458 72382
rect 19742 72434 19794 72446
rect 19742 72370 19794 72382
rect 21646 72434 21698 72446
rect 21646 72370 21698 72382
rect 22878 72434 22930 72446
rect 25106 72382 25118 72434
rect 25170 72382 25182 72434
rect 33506 72382 33518 72434
rect 33570 72382 33582 72434
rect 22878 72370 22930 72382
rect 17054 72322 17106 72334
rect 17054 72258 17106 72270
rect 1344 72154 48608 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 48608 72154
rect 1344 72068 48608 72102
rect 25342 71986 25394 71998
rect 25342 71922 25394 71934
rect 31166 71986 31218 71998
rect 31166 71922 31218 71934
rect 31950 71986 32002 71998
rect 31950 71922 32002 71934
rect 18734 71874 18786 71886
rect 18734 71810 18786 71822
rect 20750 71874 20802 71886
rect 20750 71810 20802 71822
rect 29822 71874 29874 71886
rect 29822 71810 29874 71822
rect 30494 71874 30546 71886
rect 30494 71810 30546 71822
rect 31390 71874 31442 71886
rect 31390 71810 31442 71822
rect 32174 71874 32226 71886
rect 32174 71810 32226 71822
rect 32286 71874 32338 71886
rect 32286 71810 32338 71822
rect 19742 71762 19794 71774
rect 24334 71762 24386 71774
rect 21858 71710 21870 71762
rect 21922 71710 21934 71762
rect 22642 71710 22654 71762
rect 22706 71710 22718 71762
rect 19742 71698 19794 71710
rect 24334 71698 24386 71710
rect 30046 71762 30098 71774
rect 30046 71698 30098 71710
rect 30718 71762 30770 71774
rect 37102 71762 37154 71774
rect 33842 71710 33854 71762
rect 33906 71710 33918 71762
rect 35074 71710 35086 71762
rect 35138 71710 35150 71762
rect 35634 71710 35646 71762
rect 35698 71710 35710 71762
rect 35858 71710 35870 71762
rect 35922 71710 35934 71762
rect 30718 71698 30770 71710
rect 37102 71698 37154 71710
rect 37550 71762 37602 71774
rect 37550 71698 37602 71710
rect 37774 71762 37826 71774
rect 37774 71698 37826 71710
rect 30270 71650 30322 71662
rect 33182 71650 33234 71662
rect 37326 71650 37378 71662
rect 18498 71598 18510 71650
rect 18562 71598 18574 71650
rect 22754 71598 22766 71650
rect 22818 71598 22830 71650
rect 23762 71598 23774 71650
rect 23826 71598 23838 71650
rect 31042 71598 31054 71650
rect 31106 71598 31118 71650
rect 34066 71598 34078 71650
rect 34130 71598 34142 71650
rect 35746 71598 35758 71650
rect 35810 71598 35822 71650
rect 30270 71586 30322 71598
rect 33182 71586 33234 71598
rect 37326 71586 37378 71598
rect 1344 71370 48608 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 48608 71370
rect 1344 71284 48608 71318
rect 19854 71202 19906 71214
rect 19854 71138 19906 71150
rect 32510 71202 32562 71214
rect 35858 71150 35870 71202
rect 35922 71150 35934 71202
rect 32510 71138 32562 71150
rect 6302 71090 6354 71102
rect 6302 71026 6354 71038
rect 9214 71090 9266 71102
rect 26462 71090 26514 71102
rect 12786 71038 12798 71090
rect 12850 71038 12862 71090
rect 16594 71038 16606 71090
rect 16658 71038 16670 71090
rect 18946 71038 18958 71090
rect 19010 71038 19022 71090
rect 23090 71038 23102 71090
rect 23154 71038 23166 71090
rect 9214 71026 9266 71038
rect 26462 71026 26514 71038
rect 31390 71090 31442 71102
rect 31390 71026 31442 71038
rect 19630 70978 19682 70990
rect 8418 70926 8430 70978
rect 8482 70926 8494 70978
rect 9986 70926 9998 70978
rect 10050 70926 10062 70978
rect 13682 70926 13694 70978
rect 13746 70926 13758 70978
rect 17826 70926 17838 70978
rect 17890 70926 17902 70978
rect 18274 70926 18286 70978
rect 18338 70926 18350 70978
rect 19630 70914 19682 70926
rect 20078 70978 20130 70990
rect 20078 70914 20130 70926
rect 22430 70978 22482 70990
rect 26574 70978 26626 70990
rect 32958 70978 33010 70990
rect 24546 70926 24558 70978
rect 24610 70926 24622 70978
rect 26898 70926 26910 70978
rect 26962 70926 26974 70978
rect 29922 70926 29934 70978
rect 29986 70926 29998 70978
rect 30930 70926 30942 70978
rect 30994 70926 31006 70978
rect 22430 70914 22482 70926
rect 26574 70914 26626 70926
rect 32958 70914 33010 70926
rect 33182 70978 33234 70990
rect 33182 70914 33234 70926
rect 33406 70978 33458 70990
rect 33954 70926 33966 70978
rect 34018 70926 34030 70978
rect 34850 70926 34862 70978
rect 34914 70926 34926 70978
rect 35970 70926 35982 70978
rect 36034 70926 36046 70978
rect 37986 70926 37998 70978
rect 38050 70926 38062 70978
rect 38546 70926 38558 70978
rect 38610 70926 38622 70978
rect 33406 70914 33458 70926
rect 2270 70866 2322 70878
rect 2270 70802 2322 70814
rect 8206 70866 8258 70878
rect 19406 70866 19458 70878
rect 23550 70866 23602 70878
rect 10658 70814 10670 70866
rect 10722 70814 10734 70866
rect 14466 70814 14478 70866
rect 14530 70814 14542 70866
rect 20514 70814 20526 70866
rect 20578 70814 20590 70866
rect 8206 70802 8258 70814
rect 19406 70802 19458 70814
rect 23550 70802 23602 70814
rect 25006 70866 25058 70878
rect 29474 70814 29486 70866
rect 29538 70814 29550 70866
rect 36978 70814 36990 70866
rect 37042 70814 37054 70866
rect 25006 70802 25058 70814
rect 1710 70754 1762 70766
rect 1710 70690 1762 70702
rect 6190 70754 6242 70766
rect 6190 70690 6242 70702
rect 6974 70754 7026 70766
rect 6974 70690 7026 70702
rect 7422 70754 7474 70766
rect 7422 70690 7474 70702
rect 8654 70754 8706 70766
rect 8654 70690 8706 70702
rect 8766 70754 8818 70766
rect 8766 70690 8818 70702
rect 17166 70754 17218 70766
rect 17166 70690 17218 70702
rect 21422 70754 21474 70766
rect 21422 70690 21474 70702
rect 28702 70754 28754 70766
rect 28702 70690 28754 70702
rect 39118 70754 39170 70766
rect 39118 70690 39170 70702
rect 48190 70754 48242 70766
rect 48190 70690 48242 70702
rect 1344 70586 48608 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 48608 70586
rect 1344 70500 48608 70534
rect 1822 70418 1874 70430
rect 1822 70354 1874 70366
rect 7646 70418 7698 70430
rect 7646 70354 7698 70366
rect 10446 70418 10498 70430
rect 10446 70354 10498 70366
rect 22430 70418 22482 70430
rect 22430 70354 22482 70366
rect 25902 70418 25954 70430
rect 25902 70354 25954 70366
rect 34974 70418 35026 70430
rect 34974 70354 35026 70366
rect 35086 70418 35138 70430
rect 35086 70354 35138 70366
rect 38894 70418 38946 70430
rect 38894 70354 38946 70366
rect 8766 70306 8818 70318
rect 8766 70242 8818 70254
rect 8990 70306 9042 70318
rect 8990 70242 9042 70254
rect 18398 70306 18450 70318
rect 18398 70242 18450 70254
rect 19742 70306 19794 70318
rect 19742 70242 19794 70254
rect 20190 70306 20242 70318
rect 26014 70306 26066 70318
rect 24546 70254 24558 70306
rect 24610 70254 24622 70306
rect 20190 70242 20242 70254
rect 26014 70242 26066 70254
rect 26462 70306 26514 70318
rect 26462 70242 26514 70254
rect 28478 70306 28530 70318
rect 28478 70242 28530 70254
rect 30046 70306 30098 70318
rect 39006 70306 39058 70318
rect 33954 70254 33966 70306
rect 34018 70254 34030 70306
rect 35522 70254 35534 70306
rect 35586 70254 35598 70306
rect 37762 70254 37774 70306
rect 37826 70254 37838 70306
rect 30046 70242 30098 70254
rect 39006 70242 39058 70254
rect 8206 70194 8258 70206
rect 18286 70194 18338 70206
rect 21870 70194 21922 70206
rect 27358 70194 27410 70206
rect 30942 70194 30994 70206
rect 39566 70194 39618 70206
rect 7186 70142 7198 70194
rect 7250 70142 7262 70194
rect 10210 70142 10222 70194
rect 10274 70142 10286 70194
rect 12450 70142 12462 70194
rect 12514 70142 12526 70194
rect 17714 70142 17726 70194
rect 17778 70142 17790 70194
rect 19058 70142 19070 70194
rect 19122 70142 19134 70194
rect 21298 70142 21310 70194
rect 21362 70142 21374 70194
rect 23650 70142 23662 70194
rect 23714 70142 23726 70194
rect 27122 70142 27134 70194
rect 27186 70142 27198 70194
rect 29026 70142 29038 70194
rect 29090 70142 29102 70194
rect 30482 70142 30494 70194
rect 30546 70142 30558 70194
rect 32946 70142 32958 70194
rect 33010 70142 33022 70194
rect 33730 70142 33742 70194
rect 33794 70142 33806 70194
rect 36866 70142 36878 70194
rect 36930 70142 36942 70194
rect 37650 70142 37662 70194
rect 37714 70142 37726 70194
rect 8206 70130 8258 70142
rect 18286 70130 18338 70142
rect 21870 70130 21922 70142
rect 27358 70130 27410 70142
rect 30942 70130 30994 70142
rect 39566 70130 39618 70142
rect 9774 70082 9826 70094
rect 16830 70082 16882 70094
rect 20638 70082 20690 70094
rect 4274 70030 4286 70082
rect 4338 70030 4350 70082
rect 6402 70030 6414 70082
rect 6466 70030 6478 70082
rect 8642 70030 8654 70082
rect 8706 70030 8718 70082
rect 13122 70030 13134 70082
rect 13186 70030 13198 70082
rect 15250 70030 15262 70082
rect 15314 70030 15326 70082
rect 19282 70030 19294 70082
rect 19346 70030 19358 70082
rect 9774 70018 9826 70030
rect 16830 70018 16882 70030
rect 20638 70018 20690 70030
rect 21982 70082 22034 70094
rect 25454 70082 25506 70094
rect 23538 70030 23550 70082
rect 23602 70030 23614 70082
rect 29362 70030 29374 70082
rect 29426 70030 29438 70082
rect 33618 70030 33630 70082
rect 33682 70030 33694 70082
rect 21982 70018 22034 70030
rect 25454 70018 25506 70030
rect 8430 69970 8482 69982
rect 8430 69906 8482 69918
rect 25790 69970 25842 69982
rect 25790 69906 25842 69918
rect 35198 69970 35250 69982
rect 35198 69906 35250 69918
rect 38782 69970 38834 69982
rect 38782 69906 38834 69918
rect 1344 69802 48608 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 48608 69802
rect 1344 69716 48608 69750
rect 22542 69634 22594 69646
rect 22542 69570 22594 69582
rect 22766 69634 22818 69646
rect 22766 69570 22818 69582
rect 23438 69634 23490 69646
rect 23438 69570 23490 69582
rect 27806 69634 27858 69646
rect 27806 69570 27858 69582
rect 29374 69634 29426 69646
rect 29374 69570 29426 69582
rect 33406 69634 33458 69646
rect 33406 69570 33458 69582
rect 36430 69634 36482 69646
rect 38434 69582 38446 69634
rect 38498 69582 38510 69634
rect 36430 69570 36482 69582
rect 17726 69522 17778 69534
rect 12786 69470 12798 69522
rect 12850 69470 12862 69522
rect 17042 69470 17054 69522
rect 17106 69470 17118 69522
rect 17490 69470 17502 69522
rect 17554 69470 17566 69522
rect 17726 69458 17778 69470
rect 18734 69522 18786 69534
rect 18734 69458 18786 69470
rect 25006 69522 25058 69534
rect 28030 69522 28082 69534
rect 35646 69522 35698 69534
rect 25890 69470 25902 69522
rect 25954 69470 25966 69522
rect 29698 69470 29710 69522
rect 29762 69470 29774 69522
rect 25006 69458 25058 69470
rect 28030 69458 28082 69470
rect 35646 69458 35698 69470
rect 37998 69522 38050 69534
rect 41806 69522 41858 69534
rect 39106 69470 39118 69522
rect 39170 69470 39182 69522
rect 37998 69458 38050 69470
rect 41806 69458 41858 69470
rect 6190 69410 6242 69422
rect 6190 69346 6242 69358
rect 6414 69410 6466 69422
rect 6414 69346 6466 69358
rect 8430 69410 8482 69422
rect 8430 69346 8482 69358
rect 8766 69410 8818 69422
rect 22318 69410 22370 69422
rect 9986 69358 9998 69410
rect 10050 69358 10062 69410
rect 14130 69358 14142 69410
rect 14194 69358 14206 69410
rect 8766 69346 8818 69358
rect 22318 69346 22370 69358
rect 22990 69410 23042 69422
rect 26574 69410 26626 69422
rect 25666 69358 25678 69410
rect 25730 69358 25742 69410
rect 22990 69346 23042 69358
rect 26574 69346 26626 69358
rect 26798 69410 26850 69422
rect 37102 69410 37154 69422
rect 42702 69410 42754 69422
rect 33394 69358 33406 69410
rect 33458 69358 33470 69410
rect 37314 69358 37326 69410
rect 37378 69358 37390 69410
rect 39218 69358 39230 69410
rect 39282 69358 39294 69410
rect 42242 69358 42254 69410
rect 42306 69358 42318 69410
rect 26798 69346 26850 69358
rect 37102 69346 37154 69358
rect 42702 69346 42754 69358
rect 6638 69298 6690 69310
rect 6638 69234 6690 69246
rect 7982 69298 8034 69310
rect 27134 69298 27186 69310
rect 29598 69298 29650 69310
rect 10658 69246 10670 69298
rect 10722 69246 10734 69298
rect 14914 69246 14926 69298
rect 14978 69246 14990 69298
rect 27458 69246 27470 69298
rect 27522 69246 27534 69298
rect 7982 69234 8034 69246
rect 27134 69234 27186 69246
rect 29598 69234 29650 69246
rect 33070 69298 33122 69310
rect 33070 69234 33122 69246
rect 36318 69298 36370 69310
rect 36318 69234 36370 69246
rect 7086 69186 7138 69198
rect 5842 69134 5854 69186
rect 5906 69134 5918 69186
rect 7086 69122 7138 69134
rect 24222 69186 24274 69198
rect 24222 69122 24274 69134
rect 24670 69186 24722 69198
rect 24670 69122 24722 69134
rect 26686 69186 26738 69198
rect 26686 69122 26738 69134
rect 35198 69186 35250 69198
rect 35198 69122 35250 69134
rect 1344 69018 48608 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 48608 69018
rect 1344 68932 48608 68966
rect 27134 68850 27186 68862
rect 33730 68798 33742 68850
rect 33794 68798 33806 68850
rect 27134 68786 27186 68798
rect 6414 68738 6466 68750
rect 23438 68738 23490 68750
rect 6414 68674 6466 68686
rect 8082 68674 8094 68726
rect 8146 68674 8158 68726
rect 23438 68674 23490 68686
rect 25454 68738 25506 68750
rect 48190 68738 48242 68750
rect 34290 68686 34302 68738
rect 34354 68686 34366 68738
rect 25454 68674 25506 68686
rect 48190 68674 48242 68686
rect 5854 68626 5906 68638
rect 1810 68574 1822 68626
rect 1874 68574 1886 68626
rect 5854 68562 5906 68574
rect 6078 68626 6130 68638
rect 9550 68626 9602 68638
rect 24334 68626 24386 68638
rect 38670 68626 38722 68638
rect 8306 68574 8318 68626
rect 8370 68574 8382 68626
rect 23874 68574 23886 68626
rect 23938 68574 23950 68626
rect 26114 68574 26126 68626
rect 26178 68574 26190 68626
rect 33618 68574 33630 68626
rect 33682 68574 33694 68626
rect 34178 68574 34190 68626
rect 34242 68574 34254 68626
rect 39554 68574 39566 68626
rect 39618 68574 39630 68626
rect 6078 68562 6130 68574
rect 9550 68562 9602 68574
rect 24334 68562 24386 68574
rect 38670 68562 38722 68574
rect 2270 68514 2322 68526
rect 2270 68450 2322 68462
rect 5966 68514 6018 68526
rect 27918 68514 27970 68526
rect 7298 68462 7310 68514
rect 7362 68462 7374 68514
rect 7970 68462 7982 68514
rect 8034 68462 8046 68514
rect 9986 68462 9998 68514
rect 10050 68462 10062 68514
rect 26226 68462 26238 68514
rect 26290 68462 26302 68514
rect 5966 68450 6018 68462
rect 27918 68450 27970 68462
rect 35198 68514 35250 68526
rect 35198 68450 35250 68462
rect 35758 68514 35810 68526
rect 35758 68450 35810 68462
rect 39118 68514 39170 68526
rect 40002 68462 40014 68514
rect 40066 68462 40078 68514
rect 39118 68450 39170 68462
rect 35086 68402 35138 68414
rect 35086 68338 35138 68350
rect 38782 68402 38834 68414
rect 38782 68338 38834 68350
rect 1344 68234 48608 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 48608 68234
rect 1344 68148 48608 68182
rect 24322 68014 24334 68066
rect 24386 68063 24398 68066
rect 24770 68063 24782 68066
rect 24386 68017 24782 68063
rect 24386 68014 24398 68017
rect 24770 68014 24782 68017
rect 24834 68014 24846 68066
rect 1822 67954 1874 67966
rect 1822 67890 1874 67902
rect 6638 67954 6690 67966
rect 8206 67954 8258 67966
rect 24782 67954 24834 67966
rect 7634 67902 7646 67954
rect 7698 67902 7710 67954
rect 20738 67902 20750 67954
rect 20802 67902 20814 67954
rect 6638 67890 6690 67902
rect 8206 67890 8258 67902
rect 24782 67890 24834 67902
rect 29150 67954 29202 67966
rect 34066 67902 34078 67954
rect 34130 67902 34142 67954
rect 39778 67902 39790 67954
rect 39842 67902 39854 67954
rect 40450 67902 40462 67954
rect 40514 67902 40526 67954
rect 29150 67890 29202 67902
rect 7198 67842 7250 67854
rect 26238 67842 26290 67854
rect 10098 67790 10110 67842
rect 10162 67790 10174 67842
rect 17378 67790 17390 67842
rect 17442 67790 17454 67842
rect 17938 67790 17950 67842
rect 18002 67790 18014 67842
rect 7198 67778 7250 67790
rect 26238 67778 26290 67790
rect 26462 67842 26514 67854
rect 27022 67842 27074 67854
rect 26786 67790 26798 67842
rect 26850 67790 26862 67842
rect 26462 67778 26514 67790
rect 27022 67778 27074 67790
rect 27358 67842 27410 67854
rect 30046 67842 30098 67854
rect 32958 67842 33010 67854
rect 43150 67842 43202 67854
rect 29810 67790 29822 67842
rect 29874 67790 29886 67842
rect 32386 67790 32398 67842
rect 32450 67790 32462 67842
rect 34402 67790 34414 67842
rect 34466 67790 34478 67842
rect 35746 67790 35758 67842
rect 35810 67790 35822 67842
rect 39106 67790 39118 67842
rect 39170 67839 39182 67842
rect 39330 67839 39342 67842
rect 39170 67793 39342 67839
rect 39170 67790 39182 67793
rect 39330 67790 39342 67793
rect 39394 67790 39406 67842
rect 39666 67790 39678 67842
rect 39730 67790 39742 67842
rect 40562 67790 40574 67842
rect 40626 67790 40638 67842
rect 27358 67778 27410 67790
rect 30046 67778 30098 67790
rect 32958 67778 33010 67790
rect 43150 67778 43202 67790
rect 7534 67730 7586 67742
rect 7534 67666 7586 67678
rect 10334 67730 10386 67742
rect 33070 67730 33122 67742
rect 43598 67730 43650 67742
rect 18610 67678 18622 67730
rect 18674 67678 18686 67730
rect 33394 67678 33406 67730
rect 33458 67678 33470 67730
rect 40898 67678 40910 67730
rect 40962 67678 40974 67730
rect 10334 67666 10386 67678
rect 33070 67666 33122 67678
rect 43598 67666 43650 67678
rect 43822 67730 43874 67742
rect 43822 67666 43874 67678
rect 7758 67618 7810 67630
rect 7758 67554 7810 67566
rect 15262 67618 15314 67630
rect 15262 67554 15314 67566
rect 17390 67618 17442 67630
rect 17390 67554 17442 67566
rect 26350 67618 26402 67630
rect 26350 67554 26402 67566
rect 27246 67618 27298 67630
rect 27246 67554 27298 67566
rect 27918 67618 27970 67630
rect 27918 67554 27970 67566
rect 28366 67618 28418 67630
rect 28366 67554 28418 67566
rect 30718 67618 30770 67630
rect 30718 67554 30770 67566
rect 31054 67618 31106 67630
rect 31054 67554 31106 67566
rect 31726 67618 31778 67630
rect 31726 67554 31778 67566
rect 43486 67618 43538 67630
rect 43486 67554 43538 67566
rect 1344 67450 48608 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 48608 67450
rect 1344 67364 48608 67398
rect 36206 67282 36258 67294
rect 14578 67230 14590 67282
rect 14642 67230 14654 67282
rect 36206 67218 36258 67230
rect 39230 67282 39282 67294
rect 39230 67218 39282 67230
rect 6750 67170 6802 67182
rect 6750 67106 6802 67118
rect 18622 67170 18674 67182
rect 18622 67106 18674 67118
rect 23326 67170 23378 67182
rect 33182 67170 33234 67182
rect 30818 67118 30830 67170
rect 30882 67118 30894 67170
rect 23326 67106 23378 67118
rect 33182 67106 33234 67118
rect 33406 67170 33458 67182
rect 36318 67170 36370 67182
rect 34066 67118 34078 67170
rect 34130 67118 34142 67170
rect 33406 67106 33458 67118
rect 36318 67106 36370 67118
rect 41022 67170 41074 67182
rect 41022 67106 41074 67118
rect 42926 67170 42978 67182
rect 42926 67106 42978 67118
rect 7086 67058 7138 67070
rect 13918 67058 13970 67070
rect 15038 67058 15090 67070
rect 9874 67006 9886 67058
rect 9938 67006 9950 67058
rect 14466 67006 14478 67058
rect 14530 67006 14542 67058
rect 14802 67006 14814 67058
rect 14866 67006 14878 67058
rect 7086 66994 7138 67006
rect 13918 66994 13970 67006
rect 15038 66994 15090 67006
rect 18286 67058 18338 67070
rect 28366 67058 28418 67070
rect 33070 67058 33122 67070
rect 36094 67058 36146 67070
rect 20626 67006 20638 67058
rect 20690 67006 20702 67058
rect 26674 67006 26686 67058
rect 26738 67006 26750 67058
rect 27682 67006 27694 67058
rect 27746 67006 27758 67058
rect 29138 67006 29150 67058
rect 29202 67006 29214 67058
rect 30258 67006 30270 67058
rect 30322 67006 30334 67058
rect 30706 67006 30718 67058
rect 30770 67006 30782 67058
rect 35298 67006 35310 67058
rect 35362 67006 35374 67058
rect 35634 67006 35646 67058
rect 35698 67006 35710 67058
rect 18286 66994 18338 67006
rect 28366 66994 28418 67006
rect 33070 66994 33122 67006
rect 36094 66994 36146 67006
rect 39006 67058 39058 67070
rect 39006 66994 39058 67006
rect 39118 67058 39170 67070
rect 39118 66994 39170 67006
rect 39454 67058 39506 67070
rect 44382 67058 44434 67070
rect 41906 67006 41918 67058
rect 41970 67006 41982 67058
rect 43362 67006 43374 67058
rect 43426 67006 43438 67058
rect 44594 67006 44606 67058
rect 44658 67006 44670 67058
rect 39454 66994 39506 67006
rect 44382 66994 44434 67006
rect 15486 66946 15538 66958
rect 10546 66894 10558 66946
rect 10610 66894 10622 66946
rect 12674 66894 12686 66946
rect 12738 66894 12750 66946
rect 15486 66882 15538 66894
rect 15934 66946 15986 66958
rect 25454 66946 25506 66958
rect 31838 66946 31890 66958
rect 20738 66894 20750 66946
rect 20802 66894 20814 66946
rect 22978 66894 22990 66946
rect 23042 66894 23054 66946
rect 26562 66894 26574 66946
rect 26626 66894 26638 66946
rect 30818 66894 30830 66946
rect 30882 66894 30894 66946
rect 41346 66894 41358 66946
rect 41410 66894 41422 66946
rect 43250 66894 43262 66946
rect 43314 66894 43326 66946
rect 15934 66882 15986 66894
rect 25454 66882 25506 66894
rect 31838 66882 31890 66894
rect 44270 66834 44322 66846
rect 14466 66782 14478 66834
rect 14530 66782 14542 66834
rect 26226 66782 26238 66834
rect 26290 66782 26302 66834
rect 29362 66782 29374 66834
rect 29426 66782 29438 66834
rect 44270 66770 44322 66782
rect 1344 66666 48608 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 48608 66666
rect 1344 66580 48608 66614
rect 12238 66498 12290 66510
rect 12238 66434 12290 66446
rect 14142 66498 14194 66510
rect 37550 66498 37602 66510
rect 14690 66446 14702 66498
rect 14754 66446 14766 66498
rect 35634 66446 35646 66498
rect 35698 66446 35710 66498
rect 14142 66434 14194 66446
rect 37550 66434 37602 66446
rect 27358 66386 27410 66398
rect 6514 66334 6526 66386
rect 6578 66334 6590 66386
rect 19058 66334 19070 66386
rect 19122 66334 19134 66386
rect 24546 66334 24558 66386
rect 24610 66334 24622 66386
rect 27358 66322 27410 66334
rect 30158 66386 30210 66398
rect 32510 66386 32562 66398
rect 41358 66386 41410 66398
rect 32162 66334 32174 66386
rect 32226 66334 32238 66386
rect 34178 66334 34190 66386
rect 34242 66334 34254 66386
rect 36082 66334 36094 66386
rect 36146 66334 36158 66386
rect 38546 66334 38558 66386
rect 38610 66334 38622 66386
rect 39330 66334 39342 66386
rect 39394 66334 39406 66386
rect 30158 66322 30210 66334
rect 32510 66322 32562 66334
rect 41358 66322 41410 66334
rect 41918 66386 41970 66398
rect 41918 66322 41970 66334
rect 2270 66274 2322 66286
rect 15262 66274 15314 66286
rect 30606 66274 30658 66286
rect 32846 66274 32898 66286
rect 1810 66222 1822 66274
rect 1874 66222 1886 66274
rect 9426 66222 9438 66274
rect 9490 66222 9502 66274
rect 14466 66222 14478 66274
rect 14530 66222 14542 66274
rect 15026 66222 15038 66274
rect 15090 66222 15102 66274
rect 16258 66222 16270 66274
rect 16322 66222 16334 66274
rect 21634 66222 21646 66274
rect 21698 66222 21710 66274
rect 29474 66222 29486 66274
rect 29538 66222 29550 66274
rect 29922 66222 29934 66274
rect 29986 66222 29998 66274
rect 32050 66222 32062 66274
rect 32114 66222 32126 66274
rect 2270 66210 2322 66222
rect 15262 66210 15314 66222
rect 30606 66210 30658 66222
rect 32846 66210 32898 66222
rect 33406 66274 33458 66286
rect 42254 66274 42306 66286
rect 33730 66222 33742 66274
rect 33794 66222 33806 66274
rect 34290 66222 34302 66274
rect 34354 66222 34366 66274
rect 35858 66222 35870 66274
rect 35922 66222 35934 66274
rect 38434 66222 38446 66274
rect 38498 66222 38510 66274
rect 39218 66222 39230 66274
rect 39282 66222 39294 66274
rect 33406 66210 33458 66222
rect 42254 66210 42306 66222
rect 42590 66274 42642 66286
rect 42590 66210 42642 66222
rect 5966 66162 6018 66174
rect 11902 66162 11954 66174
rect 8642 66110 8654 66162
rect 8706 66110 8718 66162
rect 5966 66098 6018 66110
rect 11902 66098 11954 66110
rect 12238 66162 12290 66174
rect 12238 66098 12290 66110
rect 12350 66162 12402 66174
rect 12350 66098 12402 66110
rect 13806 66162 13858 66174
rect 13806 66098 13858 66110
rect 15710 66162 15762 66174
rect 37550 66162 37602 66174
rect 16930 66110 16942 66162
rect 16994 66110 17006 66162
rect 22418 66110 22430 66162
rect 22482 66110 22494 66162
rect 34402 66110 34414 66162
rect 34466 66110 34478 66162
rect 15710 66098 15762 66110
rect 37550 66098 37602 66110
rect 37662 66162 37714 66174
rect 42366 66162 42418 66174
rect 39554 66110 39566 66162
rect 39618 66110 39630 66162
rect 37662 66098 37714 66110
rect 42366 66098 42418 66110
rect 5630 66050 5682 66062
rect 5630 65986 5682 65998
rect 13022 66050 13074 66062
rect 13022 65986 13074 65998
rect 14030 66050 14082 66062
rect 15598 66050 15650 66062
rect 14914 65998 14926 66050
rect 14978 65998 14990 66050
rect 14030 65986 14082 65998
rect 15598 65986 15650 65998
rect 26462 66050 26514 66062
rect 26462 65986 26514 65998
rect 26798 66050 26850 66062
rect 26798 65986 26850 65998
rect 27806 66050 27858 66062
rect 27806 65986 27858 65998
rect 31054 66050 31106 66062
rect 31054 65986 31106 65998
rect 40574 66050 40626 66062
rect 40574 65986 40626 65998
rect 41022 66050 41074 66062
rect 41022 65986 41074 65998
rect 41246 66050 41298 66062
rect 41246 65986 41298 65998
rect 41470 66050 41522 66062
rect 41470 65986 41522 65998
rect 48190 66050 48242 66062
rect 48190 65986 48242 65998
rect 1344 65882 48608 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 48608 65882
rect 1344 65796 48608 65830
rect 1822 65714 1874 65726
rect 39230 65714 39282 65726
rect 13682 65662 13694 65714
rect 13746 65662 13758 65714
rect 14802 65662 14814 65714
rect 14866 65662 14878 65714
rect 15586 65662 15598 65714
rect 15650 65662 15662 65714
rect 38322 65662 38334 65714
rect 38386 65662 38398 65714
rect 1822 65650 1874 65662
rect 39230 65650 39282 65662
rect 39454 65714 39506 65726
rect 39454 65650 39506 65662
rect 7646 65602 7698 65614
rect 5058 65550 5070 65602
rect 5122 65550 5134 65602
rect 7646 65538 7698 65550
rect 7758 65602 7810 65614
rect 7758 65538 7810 65550
rect 12462 65602 12514 65614
rect 14142 65602 14194 65614
rect 13906 65550 13918 65602
rect 13970 65550 13982 65602
rect 12462 65538 12514 65550
rect 14142 65538 14194 65550
rect 15262 65602 15314 65614
rect 15262 65538 15314 65550
rect 16494 65602 16546 65614
rect 16494 65538 16546 65550
rect 18958 65602 19010 65614
rect 18958 65538 19010 65550
rect 20862 65602 20914 65614
rect 20862 65538 20914 65550
rect 20974 65602 21026 65614
rect 20974 65538 21026 65550
rect 24670 65602 24722 65614
rect 24670 65538 24722 65550
rect 32286 65602 32338 65614
rect 32286 65538 32338 65550
rect 34078 65602 34130 65614
rect 39678 65602 39730 65614
rect 35858 65550 35870 65602
rect 35922 65550 35934 65602
rect 38434 65550 38446 65602
rect 38498 65550 38510 65602
rect 34078 65538 34130 65550
rect 39678 65538 39730 65550
rect 40238 65602 40290 65614
rect 40238 65538 40290 65550
rect 41134 65602 41186 65614
rect 41134 65538 41186 65550
rect 41918 65602 41970 65614
rect 41918 65538 41970 65550
rect 8318 65490 8370 65502
rect 4386 65438 4398 65490
rect 4450 65438 4462 65490
rect 8318 65426 8370 65438
rect 11118 65490 11170 65502
rect 11118 65426 11170 65438
rect 11342 65490 11394 65502
rect 11342 65426 11394 65438
rect 11566 65490 11618 65502
rect 11566 65426 11618 65438
rect 11790 65490 11842 65502
rect 11790 65426 11842 65438
rect 12014 65490 12066 65502
rect 12014 65426 12066 65438
rect 12238 65490 12290 65502
rect 12238 65426 12290 65438
rect 12574 65490 12626 65502
rect 15934 65490 15986 65502
rect 32398 65490 32450 65502
rect 40014 65490 40066 65502
rect 13570 65438 13582 65490
rect 13634 65438 13646 65490
rect 14690 65438 14702 65490
rect 14754 65438 14766 65490
rect 15026 65438 15038 65490
rect 15090 65438 15102 65490
rect 20178 65438 20190 65490
rect 20242 65438 20254 65490
rect 20738 65438 20750 65490
rect 20802 65438 20814 65490
rect 21298 65438 21310 65490
rect 21362 65438 21374 65490
rect 22082 65438 22094 65490
rect 22146 65438 22158 65490
rect 30594 65438 30606 65490
rect 30658 65438 30670 65490
rect 33618 65438 33630 65490
rect 33682 65438 33694 65490
rect 36082 65438 36094 65490
rect 36146 65438 36158 65490
rect 36754 65438 36766 65490
rect 36818 65438 36830 65490
rect 37426 65438 37438 65490
rect 37490 65438 37502 65490
rect 37650 65438 37662 65490
rect 37714 65438 37726 65490
rect 38658 65438 38670 65490
rect 38722 65438 38734 65490
rect 12574 65426 12626 65438
rect 15934 65426 15986 65438
rect 32398 65426 32450 65438
rect 40014 65426 40066 65438
rect 40350 65490 40402 65502
rect 42354 65438 42366 65490
rect 42418 65438 42430 65490
rect 40350 65426 40402 65438
rect 8654 65378 8706 65390
rect 7186 65326 7198 65378
rect 7250 65326 7262 65378
rect 8654 65314 8706 65326
rect 10110 65378 10162 65390
rect 10110 65314 10162 65326
rect 10558 65378 10610 65390
rect 10558 65314 10610 65326
rect 10894 65378 10946 65390
rect 10894 65314 10946 65326
rect 16382 65378 16434 65390
rect 16382 65314 16434 65326
rect 18622 65378 18674 65390
rect 18622 65314 18674 65326
rect 19854 65378 19906 65390
rect 39566 65378 39618 65390
rect 24210 65326 24222 65378
rect 24274 65326 24286 65378
rect 30482 65326 30494 65378
rect 30546 65326 30558 65378
rect 33170 65326 33182 65378
rect 33234 65326 33246 65378
rect 36418 65326 36430 65378
rect 36482 65326 36494 65378
rect 41234 65326 41246 65378
rect 41298 65326 41310 65378
rect 42802 65326 42814 65378
rect 42866 65326 42878 65378
rect 19854 65314 19906 65326
rect 39566 65314 39618 65326
rect 7646 65266 7698 65278
rect 13694 65266 13746 65278
rect 8418 65214 8430 65266
rect 8482 65263 8494 65266
rect 8978 65263 8990 65266
rect 8482 65217 8990 65263
rect 8482 65214 8494 65217
rect 8978 65214 8990 65217
rect 9042 65214 9054 65266
rect 7646 65202 7698 65214
rect 13694 65202 13746 65214
rect 14814 65266 14866 65278
rect 14814 65202 14866 65214
rect 16270 65266 16322 65278
rect 16270 65202 16322 65214
rect 18846 65266 18898 65278
rect 24558 65266 24610 65278
rect 32510 65266 32562 65278
rect 20402 65214 20414 65266
rect 20466 65214 20478 65266
rect 30146 65214 30158 65266
rect 30210 65214 30222 65266
rect 18846 65202 18898 65214
rect 24558 65202 24610 65214
rect 32510 65202 32562 65214
rect 40910 65266 40962 65278
rect 40910 65202 40962 65214
rect 1344 65098 48608 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 48608 65098
rect 1344 65012 48608 65046
rect 8430 64930 8482 64942
rect 9886 64930 9938 64942
rect 5954 64878 5966 64930
rect 6018 64878 6030 64930
rect 9314 64878 9326 64930
rect 9378 64878 9390 64930
rect 8430 64866 8482 64878
rect 9886 64866 9938 64878
rect 13918 64930 13970 64942
rect 13918 64866 13970 64878
rect 14254 64930 14306 64942
rect 20414 64930 20466 64942
rect 17826 64878 17838 64930
rect 17890 64878 17902 64930
rect 14254 64866 14306 64878
rect 20414 64866 20466 64878
rect 35758 64930 35810 64942
rect 35758 64866 35810 64878
rect 8878 64818 8930 64830
rect 6178 64766 6190 64818
rect 6242 64766 6254 64818
rect 8878 64754 8930 64766
rect 11342 64818 11394 64830
rect 11342 64754 11394 64766
rect 15934 64818 15986 64830
rect 15934 64754 15986 64766
rect 25342 64818 25394 64830
rect 29822 64818 29874 64830
rect 35422 64818 35474 64830
rect 26114 64766 26126 64818
rect 26178 64766 26190 64818
rect 34402 64766 34414 64818
rect 34466 64766 34478 64818
rect 25342 64754 25394 64766
rect 29822 64754 29874 64766
rect 35422 64754 35474 64766
rect 37550 64818 37602 64830
rect 37550 64754 37602 64766
rect 37886 64818 37938 64830
rect 38210 64766 38222 64818
rect 38274 64766 38286 64818
rect 37886 64754 37938 64766
rect 11118 64706 11170 64718
rect 6514 64654 6526 64706
rect 6578 64654 6590 64706
rect 8978 64654 8990 64706
rect 9042 64654 9054 64706
rect 9538 64654 9550 64706
rect 9602 64654 9614 64706
rect 9874 64654 9886 64706
rect 9938 64654 9950 64706
rect 11118 64642 11170 64654
rect 12014 64706 12066 64718
rect 12014 64642 12066 64654
rect 12350 64706 12402 64718
rect 12350 64642 12402 64654
rect 12910 64706 12962 64718
rect 14926 64706 14978 64718
rect 19294 64706 19346 64718
rect 21646 64706 21698 64718
rect 14242 64654 14254 64706
rect 14306 64654 14318 64706
rect 17602 64654 17614 64706
rect 17666 64654 17678 64706
rect 19058 64654 19070 64706
rect 19122 64654 19134 64706
rect 20402 64654 20414 64706
rect 20466 64654 20478 64706
rect 21298 64654 21310 64706
rect 21362 64654 21374 64706
rect 12910 64642 12962 64654
rect 14926 64642 14978 64654
rect 19294 64642 19346 64654
rect 21646 64642 21698 64654
rect 22094 64706 22146 64718
rect 33742 64706 33794 64718
rect 25890 64654 25902 64706
rect 25954 64654 25966 64706
rect 34626 64654 34638 64706
rect 34690 64654 34702 64706
rect 38546 64654 38558 64706
rect 38610 64654 38622 64706
rect 40002 64654 40014 64706
rect 40066 64654 40078 64706
rect 40674 64654 40686 64706
rect 40738 64654 40750 64706
rect 22094 64642 22146 64654
rect 33742 64642 33794 64654
rect 7982 64594 8034 64606
rect 7982 64530 8034 64542
rect 8318 64594 8370 64606
rect 8318 64530 8370 64542
rect 8766 64594 8818 64606
rect 8766 64530 8818 64542
rect 10222 64594 10274 64606
rect 10222 64530 10274 64542
rect 10782 64594 10834 64606
rect 10782 64530 10834 64542
rect 10894 64594 10946 64606
rect 10894 64530 10946 64542
rect 11566 64594 11618 64606
rect 11566 64530 11618 64542
rect 11790 64594 11842 64606
rect 11790 64530 11842 64542
rect 12574 64594 12626 64606
rect 12574 64530 12626 64542
rect 14590 64594 14642 64606
rect 18398 64594 18450 64606
rect 19742 64594 19794 64606
rect 17266 64542 17278 64594
rect 17330 64542 17342 64594
rect 18162 64542 18174 64594
rect 18226 64542 18238 64594
rect 19506 64542 19518 64594
rect 19570 64542 19582 64594
rect 14590 64530 14642 64542
rect 18398 64530 18450 64542
rect 19742 64530 19794 64542
rect 20078 64594 20130 64606
rect 35198 64594 35250 64606
rect 21858 64542 21870 64594
rect 21922 64542 21934 64594
rect 41234 64542 41246 64594
rect 41298 64542 41310 64594
rect 20078 64530 20130 64542
rect 35198 64530 35250 64542
rect 7198 64482 7250 64494
rect 7198 64418 7250 64430
rect 10558 64482 10610 64494
rect 10558 64418 10610 64430
rect 12238 64482 12290 64494
rect 12238 64418 12290 64430
rect 12798 64482 12850 64494
rect 12798 64418 12850 64430
rect 13694 64482 13746 64494
rect 13694 64418 13746 64430
rect 15486 64482 15538 64494
rect 15486 64418 15538 64430
rect 16942 64482 16994 64494
rect 16942 64418 16994 64430
rect 17614 64482 17666 64494
rect 17614 64418 17666 64430
rect 18958 64482 19010 64494
rect 30270 64482 30322 64494
rect 21746 64430 21758 64482
rect 21810 64430 21822 64482
rect 18958 64418 19010 64430
rect 30270 64418 30322 64430
rect 31166 64482 31218 64494
rect 39666 64430 39678 64482
rect 39730 64430 39742 64482
rect 31166 64418 31218 64430
rect 1344 64314 48608 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 48608 64314
rect 1344 64228 48608 64262
rect 8990 64146 9042 64158
rect 8990 64082 9042 64094
rect 10334 64146 10386 64158
rect 10334 64082 10386 64094
rect 11006 64146 11058 64158
rect 11006 64082 11058 64094
rect 11230 64146 11282 64158
rect 11230 64082 11282 64094
rect 12014 64146 12066 64158
rect 12014 64082 12066 64094
rect 13022 64146 13074 64158
rect 39790 64146 39842 64158
rect 38434 64094 38446 64146
rect 38498 64094 38510 64146
rect 39330 64094 39342 64146
rect 39394 64094 39406 64146
rect 13022 64082 13074 64094
rect 39790 64082 39842 64094
rect 43038 64146 43090 64158
rect 43038 64082 43090 64094
rect 10782 64034 10834 64046
rect 10782 63970 10834 63982
rect 11790 64034 11842 64046
rect 11790 63970 11842 63982
rect 13918 64034 13970 64046
rect 13918 63970 13970 63982
rect 14142 64034 14194 64046
rect 14142 63970 14194 63982
rect 14590 64034 14642 64046
rect 26238 64034 26290 64046
rect 19618 63982 19630 64034
rect 19682 63982 19694 64034
rect 14590 63970 14642 63982
rect 26238 63970 26290 63982
rect 36654 64034 36706 64046
rect 36654 63970 36706 63982
rect 39902 64034 39954 64046
rect 39902 63970 39954 63982
rect 48190 64034 48242 64046
rect 48190 63970 48242 63982
rect 2270 63922 2322 63934
rect 1810 63870 1822 63922
rect 1874 63870 1886 63922
rect 2270 63858 2322 63870
rect 9774 63922 9826 63934
rect 9774 63858 9826 63870
rect 11342 63922 11394 63934
rect 11342 63858 11394 63870
rect 11678 63922 11730 63934
rect 11678 63858 11730 63870
rect 13470 63922 13522 63934
rect 23214 63922 23266 63934
rect 22754 63870 22766 63922
rect 22818 63870 22830 63922
rect 13470 63858 13522 63870
rect 23214 63858 23266 63870
rect 25454 63922 25506 63934
rect 25454 63858 25506 63870
rect 25678 63922 25730 63934
rect 25678 63858 25730 63870
rect 26014 63922 26066 63934
rect 37886 63922 37938 63934
rect 26674 63870 26686 63922
rect 26738 63870 26750 63922
rect 29586 63870 29598 63922
rect 29650 63870 29662 63922
rect 35634 63870 35646 63922
rect 35698 63870 35710 63922
rect 26014 63858 26066 63870
rect 37886 63858 37938 63870
rect 38782 63922 38834 63934
rect 44930 63870 44942 63922
rect 44994 63870 45006 63922
rect 45938 63870 45950 63922
rect 46002 63870 46014 63922
rect 38782 63858 38834 63870
rect 12574 63810 12626 63822
rect 25790 63810 25842 63822
rect 27694 63810 27746 63822
rect 13794 63758 13806 63810
rect 13858 63758 13870 63810
rect 26562 63758 26574 63810
rect 26626 63758 26638 63810
rect 12574 63746 12626 63758
rect 25790 63746 25842 63758
rect 27694 63746 27746 63758
rect 28926 63810 28978 63822
rect 28926 63746 28978 63758
rect 29262 63810 29314 63822
rect 29262 63746 29314 63758
rect 29374 63810 29426 63822
rect 29374 63746 29426 63758
rect 30046 63810 30098 63822
rect 30046 63746 30098 63758
rect 30270 63810 30322 63822
rect 30270 63746 30322 63758
rect 31502 63810 31554 63822
rect 31502 63746 31554 63758
rect 31950 63810 32002 63822
rect 36094 63810 36146 63822
rect 35186 63758 35198 63810
rect 35250 63758 35262 63810
rect 31950 63746 32002 63758
rect 36094 63746 36146 63758
rect 36430 63810 36482 63822
rect 39006 63810 39058 63822
rect 36754 63758 36766 63810
rect 36818 63758 36830 63810
rect 36430 63746 36482 63758
rect 39006 63746 39058 63758
rect 43150 63810 43202 63822
rect 45826 63758 45838 63810
rect 45890 63758 45902 63810
rect 43150 63746 43202 63758
rect 30494 63698 30546 63710
rect 30494 63634 30546 63646
rect 30942 63698 30994 63710
rect 30942 63634 30994 63646
rect 38110 63698 38162 63710
rect 38110 63634 38162 63646
rect 39678 63698 39730 63710
rect 44258 63646 44270 63698
rect 44322 63646 44334 63698
rect 39678 63634 39730 63646
rect 1344 63530 48608 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 48608 63530
rect 1344 63444 48608 63478
rect 17838 63362 17890 63374
rect 17838 63298 17890 63310
rect 18846 63362 18898 63374
rect 18846 63298 18898 63310
rect 19182 63362 19234 63374
rect 19182 63298 19234 63310
rect 19966 63362 20018 63374
rect 31950 63362 32002 63374
rect 35758 63362 35810 63374
rect 27010 63310 27022 63362
rect 27074 63310 27086 63362
rect 32274 63310 32286 63362
rect 32338 63310 32350 63362
rect 34402 63310 34414 63362
rect 34466 63310 34478 63362
rect 19966 63298 20018 63310
rect 31950 63298 32002 63310
rect 35758 63298 35810 63310
rect 42926 63362 42978 63374
rect 42926 63298 42978 63310
rect 1822 63250 1874 63262
rect 1822 63186 1874 63198
rect 6638 63250 6690 63262
rect 6638 63186 6690 63198
rect 17726 63250 17778 63262
rect 25678 63250 25730 63262
rect 20290 63198 20302 63250
rect 20354 63198 20366 63250
rect 17726 63186 17778 63198
rect 25678 63186 25730 63198
rect 29374 63250 29426 63262
rect 42254 63250 42306 63262
rect 34290 63198 34302 63250
rect 34354 63198 34366 63250
rect 29374 63186 29426 63198
rect 42254 63186 42306 63198
rect 43262 63250 43314 63262
rect 46846 63250 46898 63262
rect 44034 63198 44046 63250
rect 44098 63198 44110 63250
rect 43262 63186 43314 63198
rect 46846 63186 46898 63198
rect 17278 63138 17330 63150
rect 26574 63138 26626 63150
rect 17490 63086 17502 63138
rect 17554 63086 17566 63138
rect 18386 63086 18398 63138
rect 18450 63086 18462 63138
rect 18834 63086 18846 63138
rect 18898 63086 18910 63138
rect 26338 63086 26350 63138
rect 26402 63086 26414 63138
rect 17278 63074 17330 63086
rect 26574 63074 26626 63086
rect 27358 63138 27410 63150
rect 27358 63074 27410 63086
rect 27582 63138 27634 63150
rect 27582 63074 27634 63086
rect 31726 63138 31778 63150
rect 35422 63138 35474 63150
rect 45390 63138 45442 63150
rect 34178 63086 34190 63138
rect 34242 63086 34254 63138
rect 43922 63086 43934 63138
rect 43986 63086 43998 63138
rect 31726 63074 31778 63086
rect 35422 63074 35474 63086
rect 45390 63074 45442 63086
rect 45614 63138 45666 63150
rect 45614 63074 45666 63086
rect 46622 63138 46674 63150
rect 46622 63074 46674 63086
rect 14030 63026 14082 63038
rect 14030 62962 14082 62974
rect 14254 63026 14306 63038
rect 14254 62962 14306 62974
rect 14590 63026 14642 63038
rect 14590 62962 14642 62974
rect 18174 63026 18226 63038
rect 18174 62962 18226 62974
rect 25342 63026 25394 63038
rect 35198 63026 35250 63038
rect 29474 62974 29486 63026
rect 29538 62974 29550 63026
rect 31154 62974 31166 63026
rect 31218 62974 31230 63026
rect 25342 62962 25394 62974
rect 35198 62962 35250 62974
rect 6302 62914 6354 62926
rect 6302 62850 6354 62862
rect 16382 62914 16434 62926
rect 16382 62850 16434 62862
rect 16830 62914 16882 62926
rect 16830 62850 16882 62862
rect 19742 62914 19794 62926
rect 19742 62850 19794 62862
rect 20190 62914 20242 62926
rect 20190 62850 20242 62862
rect 28030 62914 28082 62926
rect 28030 62850 28082 62862
rect 28478 62914 28530 62926
rect 42702 62914 42754 62926
rect 31042 62862 31054 62914
rect 31106 62862 31118 62914
rect 28478 62850 28530 62862
rect 42702 62850 42754 62862
rect 42814 62914 42866 62926
rect 45938 62862 45950 62914
rect 46002 62862 46014 62914
rect 46274 62862 46286 62914
rect 46338 62862 46350 62914
rect 42814 62850 42866 62862
rect 1344 62746 48608 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 48608 62746
rect 1344 62660 48608 62694
rect 4622 62578 4674 62590
rect 4622 62514 4674 62526
rect 11118 62578 11170 62590
rect 11118 62514 11170 62526
rect 13134 62578 13186 62590
rect 13134 62514 13186 62526
rect 14702 62578 14754 62590
rect 15598 62578 15650 62590
rect 15250 62526 15262 62578
rect 15314 62526 15326 62578
rect 14702 62514 14754 62526
rect 15598 62514 15650 62526
rect 17502 62578 17554 62590
rect 17502 62514 17554 62526
rect 18174 62578 18226 62590
rect 18174 62514 18226 62526
rect 19406 62578 19458 62590
rect 19406 62514 19458 62526
rect 36766 62578 36818 62590
rect 36766 62514 36818 62526
rect 44046 62578 44098 62590
rect 45726 62578 45778 62590
rect 45266 62526 45278 62578
rect 45330 62526 45342 62578
rect 44046 62514 44098 62526
rect 45726 62514 45778 62526
rect 45950 62578 46002 62590
rect 45950 62514 46002 62526
rect 6414 62466 6466 62478
rect 16270 62466 16322 62478
rect 10658 62414 10670 62466
rect 10722 62414 10734 62466
rect 6414 62402 6466 62414
rect 16270 62402 16322 62414
rect 16606 62466 16658 62478
rect 16606 62402 16658 62414
rect 27022 62466 27074 62478
rect 27022 62402 27074 62414
rect 28030 62466 28082 62478
rect 28030 62402 28082 62414
rect 42478 62466 42530 62478
rect 42478 62402 42530 62414
rect 4958 62354 5010 62366
rect 6302 62354 6354 62366
rect 6974 62354 7026 62366
rect 5842 62302 5854 62354
rect 5906 62302 5918 62354
rect 6626 62302 6638 62354
rect 6690 62302 6702 62354
rect 4958 62290 5010 62302
rect 6302 62290 6354 62302
rect 6974 62290 7026 62302
rect 7758 62354 7810 62366
rect 7758 62290 7810 62302
rect 8430 62354 8482 62366
rect 14926 62354 14978 62366
rect 10434 62302 10446 62354
rect 10498 62302 10510 62354
rect 8430 62290 8482 62302
rect 14926 62290 14978 62302
rect 15934 62354 15986 62366
rect 15934 62290 15986 62302
rect 17278 62354 17330 62366
rect 17278 62290 17330 62302
rect 17614 62354 17666 62366
rect 17614 62290 17666 62302
rect 17950 62354 18002 62366
rect 17950 62290 18002 62302
rect 18286 62354 18338 62366
rect 33182 62354 33234 62366
rect 41582 62354 41634 62366
rect 21858 62302 21870 62354
rect 21922 62302 21934 62354
rect 29138 62302 29150 62354
rect 29202 62302 29214 62354
rect 30258 62302 30270 62354
rect 30322 62302 30334 62354
rect 31378 62302 31390 62354
rect 31442 62302 31454 62354
rect 36978 62302 36990 62354
rect 37042 62302 37054 62354
rect 18286 62290 18338 62302
rect 33182 62290 33234 62302
rect 41582 62290 41634 62302
rect 41694 62354 41746 62366
rect 41694 62290 41746 62302
rect 41806 62354 41858 62366
rect 41806 62290 41858 62302
rect 42254 62354 42306 62366
rect 43710 62354 43762 62366
rect 42914 62302 42926 62354
rect 42978 62302 42990 62354
rect 42254 62290 42306 62302
rect 43710 62290 43762 62302
rect 44046 62354 44098 62366
rect 44046 62290 44098 62302
rect 44270 62354 44322 62366
rect 44270 62290 44322 62302
rect 44942 62354 44994 62366
rect 46274 62302 46286 62354
rect 46338 62302 46350 62354
rect 44942 62290 44994 62302
rect 7310 62242 7362 62254
rect 5730 62190 5742 62242
rect 5794 62190 5806 62242
rect 7310 62178 7362 62190
rect 8990 62242 9042 62254
rect 8990 62178 9042 62190
rect 14254 62242 14306 62254
rect 14254 62178 14306 62190
rect 18846 62242 18898 62254
rect 26686 62242 26738 62254
rect 22530 62190 22542 62242
rect 22594 62190 22606 62242
rect 24658 62190 24670 62242
rect 24722 62190 24734 62242
rect 18846 62178 18898 62190
rect 26686 62178 26738 62190
rect 32174 62242 32226 62254
rect 44718 62242 44770 62254
rect 43362 62190 43374 62242
rect 43426 62190 43438 62242
rect 32174 62178 32226 62190
rect 44718 62178 44770 62190
rect 45838 62242 45890 62254
rect 45838 62178 45890 62190
rect 27246 62130 27298 62142
rect 27246 62066 27298 62078
rect 27582 62130 27634 62142
rect 36654 62130 36706 62142
rect 29362 62078 29374 62130
rect 29426 62078 29438 62130
rect 27582 62066 27634 62078
rect 36654 62066 36706 62078
rect 1344 61962 48608 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 48608 61962
rect 1344 61876 48608 61910
rect 22766 61794 22818 61806
rect 44830 61794 44882 61806
rect 29474 61742 29486 61794
rect 29538 61742 29550 61794
rect 37874 61742 37886 61794
rect 37938 61742 37950 61794
rect 40338 61742 40350 61794
rect 40402 61742 40414 61794
rect 22766 61730 22818 61742
rect 44830 61730 44882 61742
rect 21870 61682 21922 61694
rect 5058 61630 5070 61682
rect 5122 61630 5134 61682
rect 7298 61630 7310 61682
rect 7362 61630 7374 61682
rect 18274 61630 18286 61682
rect 18338 61630 18350 61682
rect 21870 61618 21922 61630
rect 27134 61682 27186 61694
rect 32734 61682 32786 61694
rect 29922 61630 29934 61682
rect 29986 61630 29998 61682
rect 42466 61630 42478 61682
rect 42530 61630 42542 61682
rect 27134 61618 27186 61630
rect 32734 61618 32786 61630
rect 6302 61570 6354 61582
rect 11230 61570 11282 61582
rect 2146 61518 2158 61570
rect 2210 61518 2222 61570
rect 10098 61518 10110 61570
rect 10162 61518 10174 61570
rect 6302 61506 6354 61518
rect 11230 61506 11282 61518
rect 12686 61570 12738 61582
rect 12686 61506 12738 61518
rect 13694 61570 13746 61582
rect 18958 61570 19010 61582
rect 15474 61518 15486 61570
rect 15538 61518 15550 61570
rect 13694 61506 13746 61518
rect 18958 61506 19010 61518
rect 20078 61570 20130 61582
rect 20078 61506 20130 61518
rect 21646 61570 21698 61582
rect 21646 61506 21698 61518
rect 22094 61570 22146 61582
rect 22094 61506 22146 61518
rect 27470 61570 27522 61582
rect 32846 61570 32898 61582
rect 29586 61518 29598 61570
rect 29650 61518 29662 61570
rect 27470 61506 27522 61518
rect 32846 61506 32898 61518
rect 37214 61570 37266 61582
rect 37214 61506 37266 61518
rect 37550 61570 37602 61582
rect 42814 61570 42866 61582
rect 38098 61518 38110 61570
rect 38162 61518 38174 61570
rect 38770 61518 38782 61570
rect 38834 61518 38846 61570
rect 41010 61518 41022 61570
rect 41074 61518 41086 61570
rect 42018 61518 42030 61570
rect 42082 61518 42094 61570
rect 37550 61506 37602 61518
rect 42814 61506 42866 61518
rect 43150 61570 43202 61582
rect 43150 61506 43202 61518
rect 5742 61458 5794 61470
rect 2930 61406 2942 61458
rect 2994 61406 3006 61458
rect 5742 61394 5794 61406
rect 5854 61458 5906 61470
rect 13022 61458 13074 61470
rect 9426 61406 9438 61458
rect 9490 61406 9502 61458
rect 11778 61406 11790 61458
rect 11842 61406 11854 61458
rect 5854 61394 5906 61406
rect 13022 61394 13074 61406
rect 13470 61458 13522 61470
rect 13470 61394 13522 61406
rect 14030 61458 14082 61470
rect 14030 61394 14082 61406
rect 14366 61458 14418 61470
rect 14366 61394 14418 61406
rect 14702 61458 14754 61470
rect 18622 61458 18674 61470
rect 16146 61406 16158 61458
rect 16210 61406 16222 61458
rect 14702 61394 14754 61406
rect 18622 61394 18674 61406
rect 19182 61458 19234 61470
rect 19182 61394 19234 61406
rect 19518 61458 19570 61470
rect 19518 61394 19570 61406
rect 19742 61458 19794 61470
rect 19742 61394 19794 61406
rect 19854 61458 19906 61470
rect 19854 61394 19906 61406
rect 20526 61458 20578 61470
rect 20526 61394 20578 61406
rect 22318 61458 22370 61470
rect 22318 61394 22370 61406
rect 22654 61458 22706 61470
rect 22654 61394 22706 61406
rect 31614 61458 31666 61470
rect 31614 61394 31666 61406
rect 31950 61458 32002 61470
rect 31950 61394 32002 61406
rect 32622 61458 32674 61470
rect 32622 61394 32674 61406
rect 33182 61458 33234 61470
rect 33182 61394 33234 61406
rect 33742 61458 33794 61470
rect 33742 61394 33794 61406
rect 37102 61458 37154 61470
rect 43038 61458 43090 61470
rect 37762 61406 37774 61458
rect 37826 61406 37838 61458
rect 37102 61394 37154 61406
rect 43038 61394 43090 61406
rect 44942 61458 44994 61470
rect 44942 61394 44994 61406
rect 6078 61346 6130 61358
rect 6078 61282 6130 61294
rect 6862 61346 6914 61358
rect 6862 61282 6914 61294
rect 10894 61346 10946 61358
rect 10894 61282 10946 61294
rect 11342 61346 11394 61358
rect 11342 61282 11394 61294
rect 11566 61346 11618 61358
rect 11566 61282 11618 61294
rect 12126 61346 12178 61358
rect 12126 61282 12178 61294
rect 12798 61346 12850 61358
rect 12798 61282 12850 61294
rect 13582 61346 13634 61358
rect 13582 61282 13634 61294
rect 18734 61346 18786 61358
rect 18734 61282 18786 61294
rect 19294 61346 19346 61358
rect 19294 61282 19346 61294
rect 20190 61346 20242 61358
rect 20190 61282 20242 61294
rect 20414 61346 20466 61358
rect 20414 61282 20466 61294
rect 22766 61346 22818 61358
rect 22766 61282 22818 61294
rect 24894 61346 24946 61358
rect 33406 61346 33458 61358
rect 27794 61294 27806 61346
rect 27858 61294 27870 61346
rect 24894 61282 24946 61294
rect 33406 61282 33458 61294
rect 33630 61346 33682 61358
rect 33630 61282 33682 61294
rect 34190 61346 34242 61358
rect 34190 61282 34242 61294
rect 48190 61346 48242 61358
rect 48190 61282 48242 61294
rect 1344 61178 48608 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 48608 61178
rect 1344 61092 48608 61126
rect 4062 61010 4114 61022
rect 4062 60946 4114 60958
rect 8654 61010 8706 61022
rect 8654 60946 8706 60958
rect 14814 61010 14866 61022
rect 31390 61010 31442 61022
rect 18050 60958 18062 61010
rect 18114 60958 18126 61010
rect 29810 60958 29822 61010
rect 29874 60958 29886 61010
rect 14814 60946 14866 60958
rect 31390 60946 31442 60958
rect 31502 61010 31554 61022
rect 37102 61010 37154 61022
rect 32498 60958 32510 61010
rect 32562 60958 32574 61010
rect 33394 60958 33406 61010
rect 33458 60958 33470 61010
rect 31502 60946 31554 60958
rect 37102 60946 37154 60958
rect 37214 61010 37266 61022
rect 41022 61010 41074 61022
rect 38434 60958 38446 61010
rect 38498 60958 38510 61010
rect 37214 60946 37266 60958
rect 41022 60946 41074 60958
rect 41918 61010 41970 61022
rect 41918 60946 41970 60958
rect 4398 60898 4450 60910
rect 16270 60898 16322 60910
rect 6626 60846 6638 60898
rect 6690 60846 6702 60898
rect 12002 60846 12014 60898
rect 12066 60846 12078 60898
rect 15922 60846 15934 60898
rect 15986 60846 15998 60898
rect 4398 60834 4450 60846
rect 16270 60834 16322 60846
rect 25230 60898 25282 60910
rect 25230 60834 25282 60846
rect 31950 60898 32002 60910
rect 31950 60834 32002 60846
rect 34862 60898 34914 60910
rect 34862 60834 34914 60846
rect 35758 60898 35810 60910
rect 35758 60834 35810 60846
rect 36318 60898 36370 60910
rect 36318 60834 36370 60846
rect 36766 60898 36818 60910
rect 41358 60898 41410 60910
rect 40002 60846 40014 60898
rect 40066 60846 40078 60898
rect 36766 60834 36818 60846
rect 41358 60834 41410 60846
rect 1710 60786 1762 60798
rect 1710 60722 1762 60734
rect 5518 60786 5570 60798
rect 5518 60722 5570 60734
rect 6414 60786 6466 60798
rect 9662 60786 9714 60798
rect 15598 60786 15650 60798
rect 6962 60734 6974 60786
rect 7026 60734 7038 60786
rect 7858 60734 7870 60786
rect 7922 60734 7934 60786
rect 8418 60734 8430 60786
rect 8482 60734 8494 60786
rect 11218 60734 11230 60786
rect 11282 60734 11294 60786
rect 6414 60722 6466 60734
rect 9662 60722 9714 60734
rect 15598 60722 15650 60734
rect 16606 60786 16658 60798
rect 16606 60722 16658 60734
rect 16942 60786 16994 60798
rect 25566 60786 25618 60798
rect 17826 60734 17838 60786
rect 17890 60734 17902 60786
rect 18498 60734 18510 60786
rect 18562 60734 18574 60786
rect 21746 60734 21758 60786
rect 21810 60734 21822 60786
rect 16942 60722 16994 60734
rect 25566 60722 25618 60734
rect 29486 60786 29538 60798
rect 29486 60722 29538 60734
rect 32958 60786 33010 60798
rect 33518 60786 33570 60798
rect 33282 60734 33294 60786
rect 33346 60734 33358 60786
rect 32958 60722 33010 60734
rect 33518 60722 33570 60734
rect 33966 60786 34018 60798
rect 33966 60722 34018 60734
rect 34750 60786 34802 60798
rect 34750 60722 34802 60734
rect 34974 60786 35026 60798
rect 35646 60786 35698 60798
rect 35298 60734 35310 60786
rect 35362 60734 35374 60786
rect 34974 60722 35026 60734
rect 35646 60722 35698 60734
rect 35982 60786 36034 60798
rect 35982 60722 36034 60734
rect 36206 60786 36258 60798
rect 36206 60722 36258 60734
rect 36990 60786 37042 60798
rect 36990 60722 37042 60734
rect 37326 60786 37378 60798
rect 40910 60786 40962 60798
rect 38658 60734 38670 60786
rect 38722 60734 38734 60786
rect 39442 60734 39454 60786
rect 39506 60734 39518 60786
rect 37326 60722 37378 60734
rect 40910 60722 40962 60734
rect 41134 60786 41186 60798
rect 41134 60722 41186 60734
rect 2270 60674 2322 60686
rect 2270 60610 2322 60622
rect 5294 60674 5346 60686
rect 15262 60674 15314 60686
rect 5954 60622 5966 60674
rect 6018 60622 6030 60674
rect 14130 60622 14142 60674
rect 14194 60622 14206 60674
rect 5294 60610 5346 60622
rect 15262 60610 15314 60622
rect 16718 60674 16770 60686
rect 28926 60674 28978 60686
rect 19170 60622 19182 60674
rect 19234 60622 19246 60674
rect 21298 60622 21310 60674
rect 21362 60622 21374 60674
rect 22418 60622 22430 60674
rect 22482 60622 22494 60674
rect 24546 60622 24558 60674
rect 24610 60622 24622 60674
rect 16718 60610 16770 60622
rect 28926 60610 28978 60622
rect 29262 60674 29314 60686
rect 29262 60610 29314 60622
rect 32174 60674 32226 60686
rect 32174 60610 32226 60622
rect 33742 60674 33794 60686
rect 33742 60610 33794 60622
rect 34526 60674 34578 60686
rect 41794 60622 41806 60674
rect 41858 60622 41870 60674
rect 34526 60610 34578 60622
rect 6302 60562 6354 60574
rect 6302 60498 6354 60510
rect 31614 60562 31666 60574
rect 36318 60562 36370 60574
rect 34178 60510 34190 60562
rect 34242 60559 34254 60562
rect 34514 60559 34526 60562
rect 34242 60513 34526 60559
rect 34242 60510 34254 60513
rect 34514 60510 34526 60513
rect 34578 60510 34590 60562
rect 31614 60498 31666 60510
rect 36318 60498 36370 60510
rect 42142 60562 42194 60574
rect 42142 60498 42194 60510
rect 1344 60394 48608 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 48608 60394
rect 1344 60308 48608 60342
rect 22766 60226 22818 60238
rect 22766 60162 22818 60174
rect 31614 60226 31666 60238
rect 31614 60162 31666 60174
rect 38222 60226 38274 60238
rect 38222 60162 38274 60174
rect 39790 60226 39842 60238
rect 40686 60226 40738 60238
rect 40114 60174 40126 60226
rect 40178 60174 40190 60226
rect 39790 60162 39842 60174
rect 40686 60162 40738 60174
rect 41022 60226 41074 60238
rect 41022 60162 41074 60174
rect 1822 60114 1874 60126
rect 17614 60114 17666 60126
rect 6738 60062 6750 60114
rect 6802 60062 6814 60114
rect 7858 60062 7870 60114
rect 7922 60062 7934 60114
rect 1822 60050 1874 60062
rect 17614 60050 17666 60062
rect 20078 60114 20130 60126
rect 20078 60050 20130 60062
rect 21870 60114 21922 60126
rect 21870 60050 21922 60062
rect 23326 60114 23378 60126
rect 32510 60114 32562 60126
rect 28578 60062 28590 60114
rect 28642 60062 28654 60114
rect 23326 60050 23378 60062
rect 32510 60050 32562 60062
rect 32846 60114 32898 60126
rect 32846 60050 32898 60062
rect 39566 60114 39618 60126
rect 39566 60050 39618 60062
rect 40462 60114 40514 60126
rect 40462 60050 40514 60062
rect 6414 60002 6466 60014
rect 19854 60002 19906 60014
rect 6850 59950 6862 60002
rect 6914 59950 6926 60002
rect 10658 59950 10670 60002
rect 10722 59950 10734 60002
rect 16930 59950 16942 60002
rect 16994 59950 17006 60002
rect 6414 59938 6466 59950
rect 19854 59938 19906 59950
rect 20190 60002 20242 60014
rect 20190 59938 20242 59950
rect 21646 60002 21698 60014
rect 21646 59938 21698 59950
rect 22094 60002 22146 60014
rect 22094 59938 22146 59950
rect 24670 60002 24722 60014
rect 24670 59938 24722 59950
rect 24894 60002 24946 60014
rect 24894 59938 24946 59950
rect 25342 60002 25394 60014
rect 33182 60002 33234 60014
rect 25666 59950 25678 60002
rect 25730 59950 25742 60002
rect 26450 59950 26462 60002
rect 26514 59950 26526 60002
rect 25342 59938 25394 59950
rect 33182 59938 33234 59950
rect 33406 60002 33458 60014
rect 33406 59938 33458 59950
rect 33630 60002 33682 60014
rect 33630 59938 33682 59950
rect 33854 60002 33906 60014
rect 33854 59938 33906 59950
rect 34862 60002 34914 60014
rect 38894 60002 38946 60014
rect 37426 59950 37438 60002
rect 37490 59950 37502 60002
rect 38322 59950 38334 60002
rect 38386 59950 38398 60002
rect 34862 59938 34914 59950
rect 38894 59938 38946 59950
rect 17166 59890 17218 59902
rect 9986 59838 9998 59890
rect 10050 59838 10062 59890
rect 17166 59826 17218 59838
rect 20526 59890 20578 59902
rect 20526 59826 20578 59838
rect 22318 59890 22370 59902
rect 22318 59826 22370 59838
rect 22654 59890 22706 59902
rect 22654 59826 22706 59838
rect 22766 59890 22818 59902
rect 22766 59826 22818 59838
rect 25118 59890 25170 59902
rect 25118 59826 25170 59838
rect 31726 59890 31778 59902
rect 31726 59826 31778 59838
rect 32174 59890 32226 59902
rect 32174 59826 32226 59838
rect 32958 59890 33010 59902
rect 32958 59826 33010 59838
rect 34190 59890 34242 59902
rect 37662 59890 37714 59902
rect 35186 59838 35198 59890
rect 35250 59838 35262 59890
rect 34190 59826 34242 59838
rect 37662 59826 37714 59838
rect 6190 59778 6242 59790
rect 6190 59714 6242 59726
rect 18286 59778 18338 59790
rect 18286 59714 18338 59726
rect 31278 59778 31330 59790
rect 31278 59714 31330 59726
rect 31614 59778 31666 59790
rect 31614 59714 31666 59726
rect 32398 59778 32450 59790
rect 32398 59714 32450 59726
rect 32622 59778 32674 59790
rect 32622 59714 32674 59726
rect 34078 59778 34130 59790
rect 36318 59778 36370 59790
rect 35970 59726 35982 59778
rect 36034 59726 36046 59778
rect 34078 59714 34130 59726
rect 36318 59714 36370 59726
rect 37102 59778 37154 59790
rect 37102 59714 37154 59726
rect 1344 59610 48608 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 48608 59610
rect 1344 59524 48608 59558
rect 7310 59442 7362 59454
rect 7310 59378 7362 59390
rect 8094 59442 8146 59454
rect 24222 59442 24274 59454
rect 21858 59390 21870 59442
rect 21922 59390 21934 59442
rect 8094 59378 8146 59390
rect 24222 59378 24274 59390
rect 25342 59442 25394 59454
rect 25342 59378 25394 59390
rect 25566 59442 25618 59454
rect 25566 59378 25618 59390
rect 37102 59442 37154 59454
rect 37762 59390 37774 59442
rect 37826 59390 37838 59442
rect 37102 59378 37154 59390
rect 23998 59330 24050 59342
rect 45838 59330 45890 59342
rect 18050 59278 18062 59330
rect 18114 59278 18126 59330
rect 31266 59278 31278 59330
rect 31330 59278 31342 59330
rect 23998 59266 24050 59278
rect 45838 59266 45890 59278
rect 9550 59218 9602 59230
rect 20638 59218 20690 59230
rect 23886 59218 23938 59230
rect 8306 59166 8318 59218
rect 8370 59166 8382 59218
rect 17938 59166 17950 59218
rect 18002 59166 18014 59218
rect 19618 59166 19630 59218
rect 19682 59166 19694 59218
rect 21410 59166 21422 59218
rect 21474 59166 21486 59218
rect 9550 59154 9602 59166
rect 20638 59154 20690 59166
rect 23886 59154 23938 59166
rect 24558 59218 24610 59230
rect 24558 59154 24610 59166
rect 25678 59218 25730 59230
rect 34078 59218 34130 59230
rect 27122 59166 27134 59218
rect 27186 59166 27198 59218
rect 31042 59166 31054 59218
rect 31106 59166 31118 59218
rect 33170 59166 33182 59218
rect 33234 59166 33246 59218
rect 25678 59154 25730 59166
rect 34078 59154 34130 59166
rect 35646 59218 35698 59230
rect 35646 59154 35698 59166
rect 36430 59218 36482 59230
rect 36430 59154 36482 59166
rect 36878 59218 36930 59230
rect 36878 59154 36930 59166
rect 36990 59218 37042 59230
rect 36990 59154 37042 59166
rect 37214 59218 37266 59230
rect 37214 59154 37266 59166
rect 37326 59218 37378 59230
rect 37326 59154 37378 59166
rect 38110 59218 38162 59230
rect 38110 59154 38162 59166
rect 38558 59218 38610 59230
rect 46274 59166 46286 59218
rect 46338 59166 46350 59218
rect 38558 59154 38610 59166
rect 5966 59106 6018 59118
rect 5966 59042 6018 59054
rect 6526 59106 6578 59118
rect 6526 59042 6578 59054
rect 6862 59106 6914 59118
rect 6862 59042 6914 59054
rect 7870 59106 7922 59118
rect 7870 59042 7922 59054
rect 9102 59106 9154 59118
rect 10558 59106 10610 59118
rect 9986 59054 9998 59106
rect 10050 59054 10062 59106
rect 9102 59042 9154 59054
rect 10558 59042 10610 59054
rect 17726 59106 17778 59118
rect 17726 59042 17778 59054
rect 23102 59106 23154 59118
rect 23102 59042 23154 59054
rect 23550 59106 23602 59118
rect 23550 59042 23602 59054
rect 26238 59106 26290 59118
rect 30606 59106 30658 59118
rect 39006 59106 39058 59118
rect 27794 59054 27806 59106
rect 27858 59054 27870 59106
rect 29922 59054 29934 59106
rect 29986 59054 29998 59106
rect 33506 59054 33518 59106
rect 33570 59054 33582 59106
rect 35970 59054 35982 59106
rect 36034 59054 36046 59106
rect 26238 59042 26290 59054
rect 30606 59042 30658 59054
rect 39006 59042 39058 59054
rect 39566 59106 39618 59118
rect 39566 59042 39618 59054
rect 39902 59106 39954 59118
rect 46162 59054 46174 59106
rect 46226 59054 46238 59106
rect 39902 59042 39954 59054
rect 5618 58942 5630 58994
rect 5682 58991 5694 58994
rect 5954 58991 5966 58994
rect 5682 58945 5966 58991
rect 5682 58942 5694 58945
rect 5954 58942 5966 58945
rect 6018 58991 6030 58994
rect 6738 58991 6750 58994
rect 6018 58945 6750 58991
rect 6018 58942 6030 58945
rect 6738 58942 6750 58945
rect 6802 58942 6814 58994
rect 1344 58826 48608 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 48608 58826
rect 1344 58740 48608 58774
rect 26910 58658 26962 58670
rect 17938 58655 17950 58658
rect 17505 58609 17950 58655
rect 6302 58546 6354 58558
rect 17505 58546 17551 58609
rect 17938 58606 17950 58609
rect 18002 58606 18014 58658
rect 22194 58606 22206 58658
rect 22258 58655 22270 58658
rect 22754 58655 22766 58658
rect 22258 58609 22766 58655
rect 22258 58606 22270 58609
rect 22754 58606 22766 58609
rect 22818 58606 22830 58658
rect 31938 58606 31950 58658
rect 32002 58606 32014 58658
rect 26910 58594 26962 58606
rect 17614 58546 17666 58558
rect 22206 58546 22258 58558
rect 43598 58546 43650 58558
rect 16370 58494 16382 58546
rect 16434 58494 16446 58546
rect 17490 58494 17502 58546
rect 17554 58494 17566 58546
rect 18834 58494 18846 58546
rect 18898 58494 18910 58546
rect 29810 58494 29822 58546
rect 29874 58494 29886 58546
rect 31378 58494 31390 58546
rect 31442 58494 31454 58546
rect 6302 58482 6354 58494
rect 17614 58482 17666 58494
rect 22206 58482 22258 58494
rect 43598 58482 43650 58494
rect 44830 58546 44882 58558
rect 45154 58494 45166 58546
rect 45218 58494 45230 58546
rect 44830 58482 44882 58494
rect 7422 58434 7474 58446
rect 6626 58382 6638 58434
rect 6690 58382 6702 58434
rect 6850 58382 6862 58434
rect 6914 58382 6926 58434
rect 7422 58370 7474 58382
rect 8766 58434 8818 58446
rect 8766 58370 8818 58382
rect 9102 58434 9154 58446
rect 18062 58434 18114 58446
rect 13458 58382 13470 58434
rect 13522 58382 13534 58434
rect 9102 58370 9154 58382
rect 18062 58370 18114 58382
rect 24110 58434 24162 58446
rect 24110 58370 24162 58382
rect 24670 58434 24722 58446
rect 24670 58370 24722 58382
rect 25790 58434 25842 58446
rect 25790 58370 25842 58382
rect 26238 58434 26290 58446
rect 26238 58370 26290 58382
rect 26350 58434 26402 58446
rect 30718 58434 30770 58446
rect 39790 58434 39842 58446
rect 43486 58434 43538 58446
rect 30146 58382 30158 58434
rect 30210 58382 30222 58434
rect 31266 58382 31278 58434
rect 31330 58382 31342 58434
rect 43138 58382 43150 58434
rect 43202 58382 43214 58434
rect 45266 58382 45278 58434
rect 45330 58382 45342 58434
rect 46946 58382 46958 58434
rect 47010 58382 47022 58434
rect 26350 58370 26402 58382
rect 30718 58370 30770 58382
rect 39790 58370 39842 58382
rect 43486 58370 43538 58382
rect 1710 58322 1762 58334
rect 1710 58258 1762 58270
rect 2494 58322 2546 58334
rect 2494 58258 2546 58270
rect 5966 58322 6018 58334
rect 5966 58258 6018 58270
rect 6078 58322 6130 58334
rect 6078 58258 6130 58270
rect 6414 58322 6466 58334
rect 6414 58258 6466 58270
rect 8318 58322 8370 58334
rect 8318 58258 8370 58270
rect 8430 58322 8482 58334
rect 8430 58258 8482 58270
rect 9438 58322 9490 58334
rect 9438 58258 9490 58270
rect 9550 58322 9602 58334
rect 18958 58322 19010 58334
rect 9550 58258 9602 58270
rect 10110 58266 10162 58278
rect 14242 58270 14254 58322
rect 14306 58270 14318 58322
rect 2046 58210 2098 58222
rect 2046 58146 2098 58158
rect 5742 58210 5794 58222
rect 5742 58146 5794 58158
rect 7534 58210 7586 58222
rect 7534 58146 7586 58158
rect 8094 58210 8146 58222
rect 8094 58146 8146 58158
rect 8878 58210 8930 58222
rect 8878 58146 8930 58158
rect 9214 58210 9266 58222
rect 9214 58146 9266 58158
rect 9774 58210 9826 58222
rect 9774 58146 9826 58158
rect 9998 58210 10050 58222
rect 18958 58258 19010 58270
rect 19182 58322 19234 58334
rect 19182 58258 19234 58270
rect 23102 58322 23154 58334
rect 23102 58258 23154 58270
rect 24222 58322 24274 58334
rect 24222 58258 24274 58270
rect 24446 58322 24498 58334
rect 24446 58258 24498 58270
rect 27022 58322 27074 58334
rect 27022 58258 27074 58270
rect 29262 58322 29314 58334
rect 29262 58258 29314 58270
rect 37886 58322 37938 58334
rect 40126 58322 40178 58334
rect 38882 58270 38894 58322
rect 38946 58270 38958 58322
rect 37886 58258 37938 58270
rect 40126 58258 40178 58270
rect 43934 58322 43986 58334
rect 43934 58258 43986 58270
rect 46398 58322 46450 58334
rect 46398 58258 46450 58270
rect 46510 58322 46562 58334
rect 48066 58270 48078 58322
rect 48130 58270 48142 58322
rect 46510 58258 46562 58270
rect 10110 58202 10162 58214
rect 10558 58210 10610 58222
rect 9998 58146 10050 58158
rect 10558 58146 10610 58158
rect 11006 58210 11058 58222
rect 11006 58146 11058 58158
rect 11454 58210 11506 58222
rect 11454 58146 11506 58158
rect 18622 58210 18674 58222
rect 18622 58146 18674 58158
rect 22654 58210 22706 58222
rect 22654 58146 22706 58158
rect 23886 58210 23938 58222
rect 23886 58146 23938 58158
rect 25006 58210 25058 58222
rect 25006 58146 25058 58158
rect 25566 58210 25618 58222
rect 25566 58146 25618 58158
rect 26126 58210 26178 58222
rect 26126 58146 26178 58158
rect 26910 58210 26962 58222
rect 26910 58146 26962 58158
rect 28590 58210 28642 58222
rect 28590 58146 28642 58158
rect 39230 58210 39282 58222
rect 39230 58146 39282 58158
rect 40014 58210 40066 58222
rect 40014 58146 40066 58158
rect 40574 58210 40626 58222
rect 40574 58146 40626 58158
rect 41134 58210 41186 58222
rect 41134 58146 41186 58158
rect 44046 58210 44098 58222
rect 44046 58146 44098 58158
rect 44270 58210 44322 58222
rect 44270 58146 44322 58158
rect 46734 58210 46786 58222
rect 46734 58146 46786 58158
rect 1344 58042 48608 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 48608 58042
rect 1344 57956 48608 57990
rect 7646 57874 7698 57886
rect 7646 57810 7698 57822
rect 9662 57874 9714 57886
rect 9662 57810 9714 57822
rect 14366 57874 14418 57886
rect 14366 57810 14418 57822
rect 18174 57874 18226 57886
rect 18174 57810 18226 57822
rect 18734 57874 18786 57886
rect 25566 57874 25618 57886
rect 24434 57822 24446 57874
rect 24498 57822 24510 57874
rect 18734 57810 18786 57822
rect 25566 57810 25618 57822
rect 25790 57874 25842 57886
rect 25790 57810 25842 57822
rect 33742 57874 33794 57886
rect 33742 57810 33794 57822
rect 38894 57874 38946 57886
rect 38894 57810 38946 57822
rect 45614 57874 45666 57886
rect 45614 57810 45666 57822
rect 45838 57874 45890 57886
rect 45838 57810 45890 57822
rect 46174 57874 46226 57886
rect 46174 57810 46226 57822
rect 3166 57762 3218 57774
rect 8766 57762 8818 57774
rect 5842 57710 5854 57762
rect 5906 57710 5918 57762
rect 3166 57698 3218 57710
rect 8766 57698 8818 57710
rect 9886 57762 9938 57774
rect 9886 57698 9938 57710
rect 10558 57762 10610 57774
rect 16718 57762 16770 57774
rect 15810 57710 15822 57762
rect 15874 57710 15886 57762
rect 10558 57698 10610 57710
rect 16718 57698 16770 57710
rect 17502 57762 17554 57774
rect 31278 57762 31330 57774
rect 20626 57710 20638 57762
rect 20690 57710 20702 57762
rect 23762 57710 23774 57762
rect 23826 57710 23838 57762
rect 28354 57710 28366 57762
rect 28418 57710 28430 57762
rect 17502 57698 17554 57710
rect 31278 57698 31330 57710
rect 33966 57762 34018 57774
rect 39118 57762 39170 57774
rect 38322 57710 38334 57762
rect 38386 57710 38398 57762
rect 33966 57698 34018 57710
rect 39118 57698 39170 57710
rect 43486 57762 43538 57774
rect 43486 57698 43538 57710
rect 45166 57762 45218 57774
rect 45166 57698 45218 57710
rect 46846 57762 46898 57774
rect 46846 57698 46898 57710
rect 3502 57650 3554 57662
rect 3502 57586 3554 57598
rect 3950 57650 4002 57662
rect 6414 57650 6466 57662
rect 4610 57598 4622 57650
rect 4674 57598 4686 57650
rect 3950 57586 4002 57598
rect 6414 57586 6466 57598
rect 6750 57650 6802 57662
rect 6750 57586 6802 57598
rect 7086 57650 7138 57662
rect 7086 57586 7138 57598
rect 9438 57650 9490 57662
rect 9438 57586 9490 57598
rect 10110 57650 10162 57662
rect 14142 57650 14194 57662
rect 10882 57598 10894 57650
rect 10946 57598 10958 57650
rect 10110 57586 10162 57598
rect 14142 57586 14194 57598
rect 14590 57650 14642 57662
rect 14590 57586 14642 57598
rect 14702 57650 14754 57662
rect 14702 57586 14754 57598
rect 15486 57650 15538 57662
rect 15486 57586 15538 57598
rect 16494 57650 16546 57662
rect 16494 57586 16546 57598
rect 16830 57650 16882 57662
rect 16830 57586 16882 57598
rect 17614 57650 17666 57662
rect 19966 57650 20018 57662
rect 25454 57650 25506 57662
rect 17938 57598 17950 57650
rect 18002 57598 18014 57650
rect 20178 57598 20190 57650
rect 20242 57598 20254 57650
rect 20514 57598 20526 57650
rect 20578 57598 20590 57650
rect 22194 57598 22206 57650
rect 22258 57598 22270 57650
rect 24546 57598 24558 57650
rect 24610 57598 24622 57650
rect 17614 57586 17666 57598
rect 19966 57586 20018 57598
rect 25454 57586 25506 57598
rect 26014 57650 26066 57662
rect 34078 57650 34130 57662
rect 26226 57598 26238 57650
rect 26290 57598 26302 57650
rect 28130 57598 28142 57650
rect 28194 57598 28206 57650
rect 29698 57598 29710 57650
rect 29762 57598 29774 57650
rect 30146 57598 30158 57650
rect 30210 57598 30222 57650
rect 26014 57586 26066 57598
rect 34078 57586 34130 57598
rect 38670 57650 38722 57662
rect 38670 57586 38722 57598
rect 39230 57650 39282 57662
rect 39230 57586 39282 57598
rect 39678 57650 39730 57662
rect 45502 57650 45554 57662
rect 42914 57598 42926 57650
rect 42978 57598 42990 57650
rect 44482 57598 44494 57650
rect 44546 57598 44558 57650
rect 39678 57586 39730 57598
rect 45502 57586 45554 57598
rect 46062 57650 46114 57662
rect 46062 57586 46114 57598
rect 6638 57538 6690 57550
rect 19406 57538 19458 57550
rect 6066 57486 6078 57538
rect 6130 57486 6142 57538
rect 8082 57486 8094 57538
rect 8146 57486 8158 57538
rect 8754 57486 8766 57538
rect 8818 57486 8830 57538
rect 11666 57486 11678 57538
rect 11730 57486 11742 57538
rect 13794 57486 13806 57538
rect 13858 57486 13870 57538
rect 6638 57474 6690 57486
rect 19406 57474 19458 57486
rect 28926 57538 28978 57550
rect 28926 57474 28978 57486
rect 29598 57538 29650 57550
rect 29598 57474 29650 57486
rect 31054 57538 31106 57550
rect 31054 57474 31106 57486
rect 33518 57538 33570 57550
rect 33518 57474 33570 57486
rect 40126 57538 40178 57550
rect 43026 57486 43038 57538
rect 43090 57486 43102 57538
rect 44258 57486 44270 57538
rect 44322 57486 44334 57538
rect 40126 57474 40178 57486
rect 8542 57426 8594 57438
rect 8542 57362 8594 57374
rect 17502 57426 17554 57438
rect 17502 57362 17554 57374
rect 18286 57426 18338 57438
rect 18286 57362 18338 57374
rect 18622 57426 18674 57438
rect 18622 57362 18674 57374
rect 18958 57426 19010 57438
rect 19854 57426 19906 57438
rect 19170 57374 19182 57426
rect 19234 57423 19246 57426
rect 19506 57423 19518 57426
rect 19234 57377 19518 57423
rect 19234 57374 19246 57377
rect 19506 57374 19518 57377
rect 19570 57374 19582 57426
rect 18958 57362 19010 57374
rect 19854 57362 19906 57374
rect 30718 57426 30770 57438
rect 30718 57362 30770 57374
rect 46174 57426 46226 57438
rect 46174 57362 46226 57374
rect 1344 57258 48608 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 48608 57258
rect 1344 57172 48608 57206
rect 15710 57090 15762 57102
rect 15710 57026 15762 57038
rect 21758 57090 21810 57102
rect 21758 57026 21810 57038
rect 22430 57090 22482 57102
rect 42130 57038 42142 57090
rect 42194 57038 42206 57090
rect 22430 57026 22482 57038
rect 12126 56978 12178 56990
rect 2706 56926 2718 56978
rect 2770 56926 2782 56978
rect 4834 56926 4846 56978
rect 4898 56926 4910 56978
rect 12126 56914 12178 56926
rect 15262 56978 15314 56990
rect 31278 56978 31330 56990
rect 22082 56926 22094 56978
rect 22146 56926 22158 56978
rect 15262 56914 15314 56926
rect 31278 56914 31330 56926
rect 36430 56978 36482 56990
rect 36430 56914 36482 56926
rect 7422 56866 7474 56878
rect 1922 56814 1934 56866
rect 1986 56814 1998 56866
rect 6178 56814 6190 56866
rect 6242 56814 6254 56866
rect 6626 56814 6638 56866
rect 6690 56814 6702 56866
rect 7422 56802 7474 56814
rect 7646 56866 7698 56878
rect 7646 56802 7698 56814
rect 7982 56866 8034 56878
rect 7982 56802 8034 56814
rect 8990 56866 9042 56878
rect 8990 56802 9042 56814
rect 9214 56866 9266 56878
rect 9214 56802 9266 56814
rect 9662 56866 9714 56878
rect 9662 56802 9714 56814
rect 9886 56866 9938 56878
rect 9886 56802 9938 56814
rect 12574 56866 12626 56878
rect 19294 56866 19346 56878
rect 28254 56866 28306 56878
rect 16818 56814 16830 56866
rect 16882 56814 16894 56866
rect 18834 56814 18846 56866
rect 18898 56814 18910 56866
rect 20066 56814 20078 56866
rect 20130 56814 20142 56866
rect 22754 56814 22766 56866
rect 22818 56814 22830 56866
rect 23874 56814 23886 56866
rect 23938 56814 23950 56866
rect 25442 56814 25454 56866
rect 25506 56814 25518 56866
rect 27346 56814 27358 56866
rect 27410 56814 27422 56866
rect 12574 56802 12626 56814
rect 19294 56802 19346 56814
rect 28254 56802 28306 56814
rect 29262 56866 29314 56878
rect 29262 56802 29314 56814
rect 30382 56866 30434 56878
rect 30382 56802 30434 56814
rect 30942 56866 30994 56878
rect 36318 56866 36370 56878
rect 40798 56866 40850 56878
rect 43374 56866 43426 56878
rect 35746 56814 35758 56866
rect 35810 56814 35822 56866
rect 40450 56814 40462 56866
rect 40514 56814 40526 56866
rect 41458 56814 41470 56866
rect 41522 56814 41534 56866
rect 30942 56802 30994 56814
rect 36318 56802 36370 56814
rect 40798 56802 40850 56814
rect 43374 56802 43426 56814
rect 43598 56866 43650 56878
rect 43598 56802 43650 56814
rect 43934 56866 43986 56878
rect 43934 56802 43986 56814
rect 44830 56866 44882 56878
rect 44830 56802 44882 56814
rect 45166 56866 45218 56878
rect 45166 56802 45218 56814
rect 7870 56754 7922 56766
rect 5954 56702 5966 56754
rect 6018 56702 6030 56754
rect 7870 56690 7922 56702
rect 11454 56754 11506 56766
rect 11454 56690 11506 56702
rect 11790 56754 11842 56766
rect 11790 56690 11842 56702
rect 12014 56754 12066 56766
rect 12014 56690 12066 56702
rect 12350 56754 12402 56766
rect 12350 56690 12402 56702
rect 13358 56754 13410 56766
rect 13358 56690 13410 56702
rect 13582 56754 13634 56766
rect 13582 56690 13634 56702
rect 13694 56754 13746 56766
rect 13694 56690 13746 56702
rect 15710 56754 15762 56766
rect 15710 56690 15762 56702
rect 15822 56754 15874 56766
rect 21982 56754 22034 56766
rect 28142 56754 28194 56766
rect 17490 56702 17502 56754
rect 17554 56702 17566 56754
rect 24098 56702 24110 56754
rect 24162 56702 24174 56754
rect 27570 56702 27582 56754
rect 27634 56702 27646 56754
rect 15822 56690 15874 56702
rect 21982 56690 22034 56702
rect 28142 56690 28194 56702
rect 30046 56754 30098 56766
rect 30046 56690 30098 56702
rect 30158 56754 30210 56766
rect 30158 56690 30210 56702
rect 30606 56754 30658 56766
rect 30606 56690 30658 56702
rect 36990 56754 37042 56766
rect 36990 56690 37042 56702
rect 43038 56754 43090 56766
rect 43038 56690 43090 56702
rect 43710 56754 43762 56766
rect 43710 56690 43762 56702
rect 9550 56642 9602 56654
rect 6626 56590 6638 56642
rect 6690 56590 6702 56642
rect 8418 56590 8430 56642
rect 8482 56590 8494 56642
rect 9550 56578 9602 56590
rect 10334 56642 10386 56654
rect 10334 56578 10386 56590
rect 11118 56642 11170 56654
rect 11118 56578 11170 56590
rect 11566 56642 11618 56654
rect 11566 56578 11618 56590
rect 19182 56642 19234 56654
rect 19182 56578 19234 56590
rect 21422 56642 21474 56654
rect 21422 56578 21474 56590
rect 22542 56642 22594 56654
rect 22542 56578 22594 56590
rect 23214 56642 23266 56654
rect 23214 56578 23266 56590
rect 26126 56642 26178 56654
rect 26126 56578 26178 56590
rect 27918 56642 27970 56654
rect 27918 56578 27970 56590
rect 29710 56642 29762 56654
rect 29710 56578 29762 56590
rect 30718 56642 30770 56654
rect 30718 56578 30770 56590
rect 31726 56642 31778 56654
rect 31726 56578 31778 56590
rect 32846 56642 32898 56654
rect 32846 56578 32898 56590
rect 33070 56642 33122 56654
rect 37102 56642 37154 56654
rect 33394 56590 33406 56642
rect 33458 56590 33470 56642
rect 33070 56578 33122 56590
rect 37102 56578 37154 56590
rect 37326 56642 37378 56654
rect 37326 56578 37378 56590
rect 38894 56642 38946 56654
rect 38894 56578 38946 56590
rect 43150 56642 43202 56654
rect 43150 56578 43202 56590
rect 44942 56642 44994 56654
rect 44942 56578 44994 56590
rect 1344 56474 48608 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 48608 56474
rect 1344 56388 48608 56422
rect 7086 56306 7138 56318
rect 7086 56242 7138 56254
rect 10446 56306 10498 56318
rect 10446 56242 10498 56254
rect 14142 56306 14194 56318
rect 14142 56242 14194 56254
rect 16942 56306 16994 56318
rect 16942 56242 16994 56254
rect 18958 56306 19010 56318
rect 25342 56306 25394 56318
rect 37102 56306 37154 56318
rect 24434 56254 24446 56306
rect 24498 56254 24510 56306
rect 28466 56254 28478 56306
rect 28530 56254 28542 56306
rect 34962 56254 34974 56306
rect 35026 56254 35038 56306
rect 18958 56242 19010 56254
rect 25342 56242 25394 56254
rect 37102 56242 37154 56254
rect 41246 56306 41298 56318
rect 41246 56242 41298 56254
rect 2046 56194 2098 56206
rect 11566 56194 11618 56206
rect 7746 56142 7758 56194
rect 7810 56142 7822 56194
rect 2046 56130 2098 56142
rect 11566 56130 11618 56142
rect 12126 56194 12178 56206
rect 12126 56130 12178 56142
rect 13470 56194 13522 56206
rect 13470 56130 13522 56142
rect 13918 56194 13970 56206
rect 13918 56130 13970 56142
rect 17502 56194 17554 56206
rect 25230 56194 25282 56206
rect 36654 56194 36706 56206
rect 20626 56142 20638 56194
rect 20690 56142 20702 56194
rect 24658 56142 24670 56194
rect 24722 56142 24734 56194
rect 26450 56142 26462 56194
rect 26514 56142 26526 56194
rect 28690 56142 28702 56194
rect 28754 56142 28766 56194
rect 33506 56142 33518 56194
rect 33570 56142 33582 56194
rect 17502 56130 17554 56142
rect 25230 56130 25282 56142
rect 36654 56130 36706 56142
rect 37214 56194 37266 56206
rect 37214 56130 37266 56142
rect 41022 56194 41074 56206
rect 41022 56130 41074 56142
rect 42030 56194 42082 56206
rect 42030 56130 42082 56142
rect 1710 56082 1762 56094
rect 11454 56082 11506 56094
rect 10658 56030 10670 56082
rect 10722 56030 10734 56082
rect 1710 56018 1762 56030
rect 11454 56018 11506 56030
rect 11790 56082 11842 56094
rect 11790 56018 11842 56030
rect 13806 56082 13858 56094
rect 13806 56018 13858 56030
rect 17614 56082 17666 56094
rect 17614 56018 17666 56030
rect 20190 56082 20242 56094
rect 25566 56082 25618 56094
rect 40910 56082 40962 56094
rect 20514 56030 20526 56082
rect 20578 56030 20590 56082
rect 22194 56030 22206 56082
rect 22258 56030 22270 56082
rect 24546 56030 24558 56082
rect 24610 56030 24622 56082
rect 27682 56030 27694 56082
rect 27746 56030 27758 56082
rect 29026 56030 29038 56082
rect 29090 56030 29102 56082
rect 34626 56030 34638 56082
rect 34690 56030 34702 56082
rect 36194 56030 36206 56082
rect 36258 56030 36270 56082
rect 37986 56030 37998 56082
rect 38050 56030 38062 56082
rect 47058 56030 47070 56082
rect 47122 56030 47134 56082
rect 20190 56018 20242 56030
rect 25566 56018 25618 56030
rect 40910 56018 40962 56030
rect 2494 55970 2546 55982
rect 2494 55906 2546 55918
rect 5070 55970 5122 55982
rect 5070 55906 5122 55918
rect 6190 55970 6242 55982
rect 6190 55906 6242 55918
rect 6526 55970 6578 55982
rect 6526 55906 6578 55918
rect 9662 55970 9714 55982
rect 9662 55906 9714 55918
rect 18398 55970 18450 55982
rect 26126 55970 26178 55982
rect 19618 55918 19630 55970
rect 19682 55918 19694 55970
rect 18398 55906 18450 55918
rect 26126 55906 26178 55918
rect 30158 55970 30210 55982
rect 30158 55906 30210 55918
rect 30606 55970 30658 55982
rect 30606 55906 30658 55918
rect 33294 55970 33346 55982
rect 38670 55970 38722 55982
rect 35858 55918 35870 55970
rect 35922 55918 35934 55970
rect 38210 55918 38222 55970
rect 38274 55918 38286 55970
rect 33294 55906 33346 55918
rect 38670 55906 38722 55918
rect 41582 55970 41634 55982
rect 41582 55906 41634 55918
rect 46734 55970 46786 55982
rect 48066 55918 48078 55970
rect 48130 55918 48142 55970
rect 46734 55906 46786 55918
rect 8318 55858 8370 55870
rect 8318 55794 8370 55806
rect 17502 55858 17554 55870
rect 17502 55794 17554 55806
rect 18734 55858 18786 55870
rect 18734 55794 18786 55806
rect 19070 55858 19122 55870
rect 19070 55794 19122 55806
rect 37102 55858 37154 55870
rect 37102 55794 37154 55806
rect 1344 55690 48608 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 48608 55690
rect 1344 55604 48608 55638
rect 13582 55522 13634 55534
rect 13582 55458 13634 55470
rect 35758 55522 35810 55534
rect 35758 55458 35810 55470
rect 26014 55410 26066 55422
rect 6066 55358 6078 55410
rect 6130 55358 6142 55410
rect 12898 55358 12910 55410
rect 12962 55358 12974 55410
rect 21522 55358 21534 55410
rect 21586 55358 21598 55410
rect 26014 55346 26066 55358
rect 28030 55410 28082 55422
rect 28030 55346 28082 55358
rect 39342 55410 39394 55422
rect 39342 55346 39394 55358
rect 45614 55410 45666 55422
rect 45614 55346 45666 55358
rect 13694 55298 13746 55310
rect 7746 55246 7758 55298
rect 7810 55246 7822 55298
rect 10098 55246 10110 55298
rect 10162 55246 10174 55298
rect 13694 55234 13746 55246
rect 16046 55298 16098 55310
rect 19294 55298 19346 55310
rect 23102 55298 23154 55310
rect 33294 55298 33346 55310
rect 16930 55246 16942 55298
rect 16994 55246 17006 55298
rect 18610 55246 18622 55298
rect 18674 55246 18686 55298
rect 20066 55246 20078 55298
rect 20130 55246 20142 55298
rect 22306 55246 22318 55298
rect 22370 55246 22382 55298
rect 23538 55246 23550 55298
rect 23602 55246 23614 55298
rect 25442 55246 25454 55298
rect 25506 55246 25518 55298
rect 27346 55246 27358 55298
rect 27410 55246 27422 55298
rect 16046 55234 16098 55246
rect 19294 55234 19346 55246
rect 23102 55234 23154 55246
rect 33294 55234 33346 55246
rect 33518 55298 33570 55310
rect 33518 55234 33570 55246
rect 34414 55298 34466 55310
rect 40798 55298 40850 55310
rect 37986 55246 37998 55298
rect 38050 55246 38062 55298
rect 34414 55234 34466 55246
rect 40798 55234 40850 55246
rect 45838 55298 45890 55310
rect 45838 55234 45890 55246
rect 46846 55298 46898 55310
rect 46846 55234 46898 55246
rect 47070 55298 47122 55310
rect 47070 55234 47122 55246
rect 15934 55186 15986 55198
rect 34190 55186 34242 55198
rect 10770 55134 10782 55186
rect 10834 55134 10846 55186
rect 17490 55134 17502 55186
rect 17554 55134 17566 55186
rect 24098 55134 24110 55186
rect 24162 55134 24174 55186
rect 27570 55134 27582 55186
rect 27634 55134 27646 55186
rect 15934 55122 15986 55134
rect 34190 55122 34242 55134
rect 35870 55186 35922 55198
rect 43934 55186 43986 55198
rect 37426 55134 37438 55186
rect 37490 55134 37502 55186
rect 39106 55134 39118 55186
rect 39170 55134 39182 55186
rect 35870 55122 35922 55134
rect 43934 55122 43986 55134
rect 13582 55074 13634 55086
rect 13582 55010 13634 55022
rect 15710 55074 15762 55086
rect 15710 55010 15762 55022
rect 19182 55074 19234 55086
rect 19182 55010 19234 55022
rect 22766 55074 22818 55086
rect 22766 55010 22818 55022
rect 22990 55074 23042 55086
rect 35758 55074 35810 55086
rect 33842 55022 33854 55074
rect 33906 55022 33918 55074
rect 34738 55022 34750 55074
rect 34802 55022 34814 55074
rect 22990 55010 23042 55022
rect 35758 55010 35810 55022
rect 40574 55074 40626 55086
rect 40574 55010 40626 55022
rect 40686 55074 40738 55086
rect 40686 55010 40738 55022
rect 41022 55074 41074 55086
rect 41022 55010 41074 55022
rect 44046 55074 44098 55086
rect 44046 55010 44098 55022
rect 44158 55074 44210 55086
rect 46162 55022 46174 55074
rect 46226 55022 46238 55074
rect 46498 55022 46510 55074
rect 46562 55022 46574 55074
rect 44158 55010 44210 55022
rect 1344 54906 48608 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 48608 54906
rect 1344 54820 48608 54854
rect 8542 54738 8594 54750
rect 8542 54674 8594 54686
rect 11902 54738 11954 54750
rect 11902 54674 11954 54686
rect 13022 54738 13074 54750
rect 13022 54674 13074 54686
rect 13470 54738 13522 54750
rect 13470 54674 13522 54686
rect 17950 54738 18002 54750
rect 17950 54674 18002 54686
rect 18174 54738 18226 54750
rect 27582 54738 27634 54750
rect 22418 54686 22430 54738
rect 22482 54686 22494 54738
rect 23314 54686 23326 54738
rect 23378 54686 23390 54738
rect 18174 54674 18226 54686
rect 27582 54674 27634 54686
rect 33518 54738 33570 54750
rect 33518 54674 33570 54686
rect 33742 54738 33794 54750
rect 33742 54674 33794 54686
rect 33966 54738 34018 54750
rect 33966 54674 34018 54686
rect 34078 54738 34130 54750
rect 34078 54674 34130 54686
rect 34190 54738 34242 54750
rect 34190 54674 34242 54686
rect 40798 54738 40850 54750
rect 44146 54686 44158 54738
rect 44210 54686 44222 54738
rect 40798 54674 40850 54686
rect 1710 54626 1762 54638
rect 10334 54626 10386 54638
rect 6178 54574 6190 54626
rect 6242 54574 6254 54626
rect 1710 54562 1762 54574
rect 10334 54562 10386 54574
rect 11790 54626 11842 54638
rect 11790 54562 11842 54574
rect 12126 54626 12178 54638
rect 12126 54562 12178 54574
rect 12350 54626 12402 54638
rect 12350 54562 12402 54574
rect 13582 54626 13634 54638
rect 13582 54562 13634 54574
rect 17614 54626 17666 54638
rect 26238 54626 26290 54638
rect 18610 54574 18622 54626
rect 18674 54574 18686 54626
rect 24322 54574 24334 54626
rect 24386 54574 24398 54626
rect 17614 54562 17666 54574
rect 26238 54562 26290 54574
rect 27134 54626 27186 54638
rect 27134 54562 27186 54574
rect 38782 54626 38834 54638
rect 41022 54626 41074 54638
rect 39218 54574 39230 54626
rect 39282 54574 39294 54626
rect 38782 54562 38834 54574
rect 41022 54562 41074 54574
rect 43262 54626 43314 54638
rect 43262 54562 43314 54574
rect 43598 54626 43650 54638
rect 46834 54574 46846 54626
rect 46898 54574 46910 54626
rect 43598 54562 43650 54574
rect 5854 54514 5906 54526
rect 8094 54514 8146 54526
rect 1922 54462 1934 54514
rect 1986 54462 1998 54514
rect 6066 54462 6078 54514
rect 6130 54462 6142 54514
rect 5854 54450 5906 54462
rect 8094 54450 8146 54462
rect 13246 54514 13298 54526
rect 17838 54514 17890 54526
rect 21198 54514 21250 54526
rect 22990 54514 23042 54526
rect 13906 54462 13918 54514
rect 13970 54462 13982 54514
rect 18498 54462 18510 54514
rect 18562 54462 18574 54514
rect 20178 54462 20190 54514
rect 20242 54462 20254 54514
rect 21970 54462 21982 54514
rect 22034 54462 22046 54514
rect 13246 54450 13298 54462
rect 17838 54450 17890 54462
rect 21198 54450 21250 54462
rect 22990 54450 23042 54462
rect 23998 54514 24050 54526
rect 23998 54450 24050 54462
rect 25566 54514 25618 54526
rect 25566 54450 25618 54462
rect 25790 54514 25842 54526
rect 25790 54450 25842 54462
rect 26014 54514 26066 54526
rect 26014 54450 26066 54462
rect 26574 54514 26626 54526
rect 26574 54450 26626 54462
rect 26910 54514 26962 54526
rect 26910 54450 26962 54462
rect 27470 54514 27522 54526
rect 33406 54514 33458 54526
rect 28466 54462 28478 54514
rect 28530 54462 28542 54514
rect 27470 54450 27522 54462
rect 33406 54450 33458 54462
rect 34638 54514 34690 54526
rect 41134 54514 41186 54526
rect 43150 54514 43202 54526
rect 45614 54514 45666 54526
rect 38322 54462 38334 54514
rect 38386 54462 38398 54514
rect 39442 54462 39454 54514
rect 39506 54462 39518 54514
rect 40002 54462 40014 54514
rect 40066 54462 40078 54514
rect 42802 54462 42814 54514
rect 42866 54462 42878 54514
rect 45266 54462 45278 54514
rect 45330 54462 45342 54514
rect 46274 54462 46286 54514
rect 46338 54462 46350 54514
rect 34638 54450 34690 54462
rect 41134 54450 41186 54462
rect 43150 54450 43202 54462
rect 45614 54450 45666 54462
rect 2494 54402 2546 54414
rect 25342 54402 25394 54414
rect 14690 54350 14702 54402
rect 14754 54350 14766 54402
rect 16818 54350 16830 54402
rect 16882 54350 16894 54402
rect 2494 54338 2546 54350
rect 25342 54338 25394 54350
rect 27022 54402 27074 54414
rect 27022 54338 27074 54350
rect 28142 54402 28194 54414
rect 32286 54402 32338 54414
rect 43822 54402 43874 54414
rect 29250 54350 29262 54402
rect 29314 54350 29326 54402
rect 31378 54350 31390 54402
rect 31442 54350 31454 54402
rect 37986 54350 37998 54402
rect 38050 54350 38062 54402
rect 39218 54350 39230 54402
rect 39282 54350 39294 54402
rect 28142 54338 28194 54350
rect 32286 54338 32338 54350
rect 43822 54338 43874 54350
rect 7086 54290 7138 54302
rect 7086 54226 7138 54238
rect 27582 54290 27634 54302
rect 32274 54238 32286 54290
rect 32338 54287 32350 54290
rect 32610 54287 32622 54290
rect 32338 54241 32622 54287
rect 32338 54238 32350 54241
rect 32610 54238 32622 54241
rect 32674 54238 32686 54290
rect 27582 54226 27634 54238
rect 1344 54122 48608 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 48608 54122
rect 1344 54036 48608 54070
rect 18622 53954 18674 53966
rect 18622 53890 18674 53902
rect 33406 53954 33458 53966
rect 38658 53902 38670 53954
rect 38722 53902 38734 53954
rect 41122 53951 41134 53954
rect 40689 53905 41134 53951
rect 33406 53890 33458 53902
rect 15038 53842 15090 53854
rect 38334 53842 38386 53854
rect 40689 53842 40735 53905
rect 41122 53902 41134 53905
rect 41186 53902 41198 53954
rect 44270 53842 44322 53854
rect 4610 53790 4622 53842
rect 4674 53790 4686 53842
rect 32050 53790 32062 53842
rect 32114 53790 32126 53842
rect 40674 53790 40686 53842
rect 40738 53790 40750 53842
rect 45938 53790 45950 53842
rect 46002 53790 46014 53842
rect 15038 53778 15090 53790
rect 38334 53778 38386 53790
rect 44270 53778 44322 53790
rect 14814 53730 14866 53742
rect 1810 53678 1822 53730
rect 1874 53678 1886 53730
rect 11218 53678 11230 53730
rect 11282 53678 11294 53730
rect 14814 53666 14866 53678
rect 15262 53730 15314 53742
rect 25902 53730 25954 53742
rect 21522 53678 21534 53730
rect 21586 53678 21598 53730
rect 23090 53678 23102 53730
rect 23154 53678 23166 53730
rect 24882 53678 24894 53730
rect 24946 53678 24958 53730
rect 15262 53666 15314 53678
rect 25902 53666 25954 53678
rect 26238 53730 26290 53742
rect 26238 53666 26290 53678
rect 26574 53730 26626 53742
rect 26574 53666 26626 53678
rect 27022 53730 27074 53742
rect 33518 53730 33570 53742
rect 29138 53678 29150 53730
rect 29202 53678 29214 53730
rect 29922 53678 29934 53730
rect 29986 53678 29998 53730
rect 27022 53666 27074 53678
rect 33518 53666 33570 53678
rect 38110 53730 38162 53742
rect 38110 53666 38162 53678
rect 41358 53730 41410 53742
rect 41358 53666 41410 53678
rect 41694 53730 41746 53742
rect 41694 53666 41746 53678
rect 41918 53730 41970 53742
rect 41918 53666 41970 53678
rect 42254 53730 42306 53742
rect 43374 53730 43426 53742
rect 42690 53678 42702 53730
rect 42754 53678 42766 53730
rect 43810 53678 43822 53730
rect 43874 53678 43886 53730
rect 46050 53678 46062 53730
rect 46114 53678 46126 53730
rect 46498 53678 46510 53730
rect 46562 53678 46574 53730
rect 46946 53678 46958 53730
rect 47010 53678 47022 53730
rect 42254 53666 42306 53678
rect 43374 53666 43426 53678
rect 15486 53618 15538 53630
rect 2482 53566 2494 53618
rect 2546 53566 2558 53618
rect 6066 53566 6078 53618
rect 6130 53566 6142 53618
rect 6850 53566 6862 53618
rect 6914 53566 6926 53618
rect 10546 53566 10558 53618
rect 10610 53566 10622 53618
rect 15486 53554 15538 53566
rect 16270 53618 16322 53630
rect 16270 53554 16322 53566
rect 18734 53618 18786 53630
rect 27582 53618 27634 53630
rect 21410 53566 21422 53618
rect 21474 53566 21486 53618
rect 24658 53566 24670 53618
rect 24722 53566 24734 53618
rect 18734 53554 18786 53566
rect 27582 53554 27634 53566
rect 27918 53618 27970 53630
rect 32946 53566 32958 53618
rect 33010 53566 33022 53618
rect 27918 53554 27970 53566
rect 41470 53562 41522 53574
rect 42914 53566 42926 53618
rect 42978 53566 42990 53618
rect 45490 53566 45502 53618
rect 45554 53566 45566 53618
rect 48066 53566 48078 53618
rect 48130 53566 48142 53618
rect 5070 53506 5122 53518
rect 16718 53506 16770 53518
rect 8306 53454 8318 53506
rect 8370 53454 8382 53506
rect 5070 53442 5122 53454
rect 16718 53442 16770 53454
rect 18622 53506 18674 53518
rect 26238 53506 26290 53518
rect 25330 53454 25342 53506
rect 25394 53454 25406 53506
rect 18622 53442 18674 53454
rect 26238 53442 26290 53454
rect 28366 53506 28418 53518
rect 28366 53442 28418 53454
rect 32622 53506 32674 53518
rect 32622 53442 32674 53454
rect 33406 53506 33458 53518
rect 33406 53442 33458 53454
rect 33966 53506 34018 53518
rect 33966 53442 34018 53454
rect 41134 53506 41186 53518
rect 41470 53498 41522 53510
rect 42030 53506 42082 53518
rect 41134 53442 41186 53454
rect 42030 53442 42082 53454
rect 1344 53338 48608 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 48608 53338
rect 1344 53252 48608 53286
rect 7534 53170 7586 53182
rect 7534 53106 7586 53118
rect 8878 53170 8930 53182
rect 8878 53106 8930 53118
rect 9774 53170 9826 53182
rect 9774 53106 9826 53118
rect 11566 53170 11618 53182
rect 11566 53106 11618 53118
rect 12014 53170 12066 53182
rect 12014 53106 12066 53118
rect 12574 53170 12626 53182
rect 12574 53106 12626 53118
rect 13806 53170 13858 53182
rect 13806 53106 13858 53118
rect 14254 53170 14306 53182
rect 14254 53106 14306 53118
rect 15598 53170 15650 53182
rect 15598 53106 15650 53118
rect 16382 53170 16434 53182
rect 16382 53106 16434 53118
rect 18286 53170 18338 53182
rect 20750 53170 20802 53182
rect 19282 53118 19294 53170
rect 19346 53118 19358 53170
rect 18286 53106 18338 53118
rect 20750 53106 20802 53118
rect 20974 53170 21026 53182
rect 20974 53106 21026 53118
rect 24782 53170 24834 53182
rect 24782 53106 24834 53118
rect 32510 53170 32562 53182
rect 32510 53106 32562 53118
rect 33966 53170 34018 53182
rect 33966 53106 34018 53118
rect 40462 53170 40514 53182
rect 40462 53106 40514 53118
rect 41918 53170 41970 53182
rect 41918 53106 41970 53118
rect 42478 53170 42530 53182
rect 42478 53106 42530 53118
rect 46734 53170 46786 53182
rect 46734 53106 46786 53118
rect 9102 53058 9154 53070
rect 9102 52994 9154 53006
rect 9550 53058 9602 53070
rect 9550 52994 9602 53006
rect 10110 53058 10162 53070
rect 10110 52994 10162 53006
rect 10558 53058 10610 53070
rect 10558 52994 10610 53006
rect 11230 53058 11282 53070
rect 11230 52994 11282 53006
rect 16270 53058 16322 53070
rect 16270 52994 16322 53006
rect 21870 53058 21922 53070
rect 23214 53058 23266 53070
rect 22642 53006 22654 53058
rect 22706 53006 22718 53058
rect 21870 52994 21922 53006
rect 23214 52994 23266 53006
rect 24446 53058 24498 53070
rect 24446 52994 24498 53006
rect 24558 53058 24610 53070
rect 24558 52994 24610 53006
rect 25678 53058 25730 53070
rect 25678 52994 25730 53006
rect 25790 53058 25842 53070
rect 25790 52994 25842 53006
rect 26014 53058 26066 53070
rect 31390 53058 31442 53070
rect 28130 53006 28142 53058
rect 28194 53006 28206 53058
rect 26014 52994 26066 53006
rect 31390 52994 31442 53006
rect 32286 53058 32338 53070
rect 32286 52994 32338 53006
rect 33742 53058 33794 53070
rect 33742 52994 33794 53006
rect 35870 53058 35922 53070
rect 35870 52994 35922 53006
rect 37438 53058 37490 53070
rect 37438 52994 37490 53006
rect 40238 53058 40290 53070
rect 41806 53058 41858 53070
rect 41234 53006 41246 53058
rect 41298 53006 41310 53058
rect 40238 52994 40290 53006
rect 41806 52994 41858 53006
rect 8766 52946 8818 52958
rect 1698 52894 1710 52946
rect 1762 52894 1774 52946
rect 4946 52894 4958 52946
rect 5010 52894 5022 52946
rect 5954 52894 5966 52946
rect 6018 52894 6030 52946
rect 6178 52894 6190 52946
rect 6242 52894 6254 52946
rect 8766 52882 8818 52894
rect 9886 52946 9938 52958
rect 9886 52882 9938 52894
rect 10334 52946 10386 52958
rect 10334 52882 10386 52894
rect 10670 52946 10722 52958
rect 10670 52882 10722 52894
rect 11902 52946 11954 52958
rect 11902 52882 11954 52894
rect 12238 52946 12290 52958
rect 12238 52882 12290 52894
rect 14142 52946 14194 52958
rect 14142 52882 14194 52894
rect 14478 52946 14530 52958
rect 14478 52882 14530 52894
rect 15262 52946 15314 52958
rect 15262 52882 15314 52894
rect 15710 52946 15762 52958
rect 15710 52882 15762 52894
rect 15822 52946 15874 52958
rect 15822 52882 15874 52894
rect 16606 52946 16658 52958
rect 18958 52946 19010 52958
rect 18498 52894 18510 52946
rect 18562 52894 18574 52946
rect 16606 52882 16658 52894
rect 18958 52882 19010 52894
rect 20638 52946 20690 52958
rect 20638 52882 20690 52894
rect 21982 52946 22034 52958
rect 31054 52946 31106 52958
rect 22418 52894 22430 52946
rect 22482 52894 22494 52946
rect 23538 52894 23550 52946
rect 23602 52894 23614 52946
rect 26898 52894 26910 52946
rect 26962 52894 26974 52946
rect 27458 52894 27470 52946
rect 27522 52894 27534 52946
rect 21982 52882 22034 52894
rect 31054 52882 31106 52894
rect 32174 52946 32226 52958
rect 32174 52882 32226 52894
rect 33630 52946 33682 52958
rect 40126 52946 40178 52958
rect 42142 52946 42194 52958
rect 36306 52894 36318 52946
rect 36370 52894 36382 52946
rect 41010 52894 41022 52946
rect 41074 52894 41086 52946
rect 33630 52882 33682 52894
rect 40126 52882 40178 52894
rect 42142 52882 42194 52894
rect 6750 52834 6802 52846
rect 2482 52782 2494 52834
rect 2546 52782 2558 52834
rect 4610 52782 4622 52834
rect 4674 52782 4686 52834
rect 6750 52770 6802 52782
rect 8094 52834 8146 52846
rect 8094 52770 8146 52782
rect 8430 52834 8482 52846
rect 8430 52770 8482 52782
rect 21422 52834 21474 52846
rect 21422 52770 21474 52782
rect 23998 52834 24050 52846
rect 23998 52770 24050 52782
rect 25454 52834 25506 52846
rect 30718 52834 30770 52846
rect 30258 52782 30270 52834
rect 30322 52782 30334 52834
rect 25454 52770 25506 52782
rect 30718 52770 30770 52782
rect 34302 52834 34354 52846
rect 42926 52834 42978 52846
rect 36754 52782 36766 52834
rect 36818 52782 36830 52834
rect 37538 52782 37550 52834
rect 37602 52782 37614 52834
rect 34302 52770 34354 52782
rect 42926 52770 42978 52782
rect 43374 52834 43426 52846
rect 43374 52770 43426 52782
rect 5406 52722 5458 52734
rect 5406 52658 5458 52670
rect 21870 52722 21922 52734
rect 21870 52658 21922 52670
rect 26238 52722 26290 52734
rect 26238 52658 26290 52670
rect 37214 52722 37266 52734
rect 37214 52658 37266 52670
rect 1344 52554 48608 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 48608 52554
rect 1344 52468 48608 52502
rect 4958 52386 5010 52398
rect 4958 52322 5010 52334
rect 18846 52386 18898 52398
rect 34974 52386 35026 52398
rect 41694 52386 41746 52398
rect 21970 52334 21982 52386
rect 22034 52334 22046 52386
rect 36082 52334 36094 52386
rect 36146 52334 36158 52386
rect 18846 52322 18898 52334
rect 34974 52322 35026 52334
rect 41694 52322 41746 52334
rect 6190 52274 6242 52286
rect 6190 52210 6242 52222
rect 6638 52274 6690 52286
rect 21646 52274 21698 52286
rect 9202 52222 9214 52274
rect 9266 52222 9278 52274
rect 10994 52222 11006 52274
rect 11058 52222 11070 52274
rect 15586 52222 15598 52274
rect 15650 52222 15662 52274
rect 17714 52222 17726 52274
rect 17778 52222 17790 52274
rect 6638 52210 6690 52222
rect 21646 52210 21698 52222
rect 22878 52274 22930 52286
rect 22878 52210 22930 52222
rect 23438 52274 23490 52286
rect 23438 52210 23490 52222
rect 32286 52274 32338 52286
rect 37986 52222 37998 52274
rect 38050 52222 38062 52274
rect 39554 52222 39566 52274
rect 39618 52222 39630 52274
rect 40338 52222 40350 52274
rect 40402 52222 40414 52274
rect 32286 52210 32338 52222
rect 4174 52162 4226 52174
rect 4174 52098 4226 52110
rect 5630 52162 5682 52174
rect 12238 52162 12290 52174
rect 7186 52110 7198 52162
rect 7250 52110 7262 52162
rect 8306 52110 8318 52162
rect 8370 52110 8382 52162
rect 9090 52110 9102 52162
rect 9154 52110 9166 52162
rect 10210 52110 10222 52162
rect 10274 52110 10286 52162
rect 5630 52098 5682 52110
rect 12238 52098 12290 52110
rect 12574 52162 12626 52174
rect 12574 52098 12626 52110
rect 12686 52162 12738 52174
rect 12686 52098 12738 52110
rect 13358 52162 13410 52174
rect 13358 52098 13410 52110
rect 13694 52162 13746 52174
rect 19182 52162 19234 52174
rect 14802 52110 14814 52162
rect 14866 52110 14878 52162
rect 13694 52098 13746 52110
rect 19182 52098 19234 52110
rect 19854 52162 19906 52174
rect 19854 52098 19906 52110
rect 21422 52162 21474 52174
rect 21422 52098 21474 52110
rect 22318 52162 22370 52174
rect 29262 52162 29314 52174
rect 23650 52110 23662 52162
rect 23714 52110 23726 52162
rect 24994 52110 25006 52162
rect 25058 52110 25070 52162
rect 25330 52110 25342 52162
rect 25394 52110 25406 52162
rect 26674 52110 26686 52162
rect 26738 52110 26750 52162
rect 28466 52110 28478 52162
rect 28530 52110 28542 52162
rect 22318 52098 22370 52110
rect 29262 52098 29314 52110
rect 31726 52162 31778 52174
rect 35086 52162 35138 52174
rect 32834 52110 32846 52162
rect 32898 52110 32910 52162
rect 31726 52098 31778 52110
rect 35086 52098 35138 52110
rect 35534 52162 35586 52174
rect 35534 52098 35586 52110
rect 35758 52162 35810 52174
rect 39118 52162 39170 52174
rect 37650 52110 37662 52162
rect 37714 52110 37726 52162
rect 37874 52110 37886 52162
rect 37938 52110 37950 52162
rect 41010 52110 41022 52162
rect 41074 52110 41086 52162
rect 35758 52098 35810 52110
rect 39118 52098 39170 52110
rect 2382 52050 2434 52062
rect 2382 51986 2434 51998
rect 2718 52050 2770 52062
rect 2718 51986 2770 51998
rect 3614 52050 3666 52062
rect 3614 51986 3666 51998
rect 4846 52050 4898 52062
rect 4846 51986 4898 51998
rect 4958 52050 5010 52062
rect 4958 51986 5010 51998
rect 6526 52050 6578 52062
rect 6526 51986 6578 51998
rect 6750 52050 6802 52062
rect 6750 51986 6802 51998
rect 13582 52050 13634 52062
rect 13582 51986 13634 51998
rect 18846 52050 18898 52062
rect 18846 51986 18898 51998
rect 18958 52050 19010 52062
rect 18958 51986 19010 51998
rect 19518 52050 19570 52062
rect 19518 51986 19570 51998
rect 20414 52050 20466 52062
rect 41806 52050 41858 52062
rect 27122 51998 27134 52050
rect 27186 51998 27198 52050
rect 32610 51998 32622 52050
rect 32674 51998 32686 52050
rect 20414 51986 20466 51998
rect 41806 51986 41858 51998
rect 42142 52050 42194 52062
rect 42142 51986 42194 51998
rect 4062 51938 4114 51950
rect 4062 51874 4114 51886
rect 12350 51938 12402 51950
rect 12350 51874 12402 51886
rect 19406 51938 19458 51950
rect 34638 51938 34690 51950
rect 26898 51886 26910 51938
rect 26962 51886 26974 51938
rect 19406 51874 19458 51886
rect 34638 51874 34690 51886
rect 34974 51938 35026 51950
rect 41694 51938 41746 51950
rect 37650 51886 37662 51938
rect 37714 51886 37726 51938
rect 34974 51874 35026 51886
rect 41694 51874 41746 51886
rect 42254 51938 42306 51950
rect 42254 51874 42306 51886
rect 42478 51938 42530 51950
rect 42478 51874 42530 51886
rect 42814 51938 42866 51950
rect 42814 51874 42866 51886
rect 1344 51770 48608 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 48608 51770
rect 1344 51684 48608 51718
rect 9774 51602 9826 51614
rect 9774 51538 9826 51550
rect 20862 51602 20914 51614
rect 20862 51538 20914 51550
rect 22318 51602 22370 51614
rect 22318 51538 22370 51550
rect 22542 51602 22594 51614
rect 22542 51538 22594 51550
rect 22766 51602 22818 51614
rect 22766 51538 22818 51550
rect 23886 51602 23938 51614
rect 35534 51602 35586 51614
rect 40910 51602 40962 51614
rect 24210 51550 24222 51602
rect 24274 51550 24286 51602
rect 38882 51550 38894 51602
rect 38946 51550 38958 51602
rect 23886 51538 23938 51550
rect 35534 51538 35586 51550
rect 40910 51538 40962 51550
rect 46622 51602 46674 51614
rect 46622 51538 46674 51550
rect 4174 51490 4226 51502
rect 20526 51490 20578 51502
rect 7298 51438 7310 51490
rect 7362 51438 7374 51490
rect 11778 51438 11790 51490
rect 11842 51438 11854 51490
rect 4174 51426 4226 51438
rect 20526 51426 20578 51438
rect 20638 51490 20690 51502
rect 43822 51490 43874 51502
rect 41234 51438 41246 51490
rect 41298 51438 41310 51490
rect 20638 51426 20690 51438
rect 43822 51426 43874 51438
rect 44046 51490 44098 51502
rect 44046 51426 44098 51438
rect 5630 51378 5682 51390
rect 8318 51378 8370 51390
rect 4722 51326 4734 51378
rect 4786 51326 4798 51378
rect 6290 51326 6302 51378
rect 6354 51326 6366 51378
rect 5630 51314 5682 51326
rect 8318 51314 8370 51326
rect 8766 51378 8818 51390
rect 22206 51378 22258 51390
rect 30718 51378 30770 51390
rect 10994 51326 11006 51378
rect 11058 51326 11070 51378
rect 25778 51326 25790 51378
rect 25842 51326 25854 51378
rect 26898 51326 26910 51378
rect 26962 51326 26974 51378
rect 28018 51326 28030 51378
rect 28082 51326 28094 51378
rect 28242 51326 28254 51378
rect 28306 51326 28318 51378
rect 29026 51326 29038 51378
rect 29090 51326 29102 51378
rect 8766 51314 8818 51326
rect 22206 51314 22258 51326
rect 30718 51314 30770 51326
rect 35422 51378 35474 51390
rect 39106 51326 39118 51378
rect 39170 51326 39182 51378
rect 42578 51326 42590 51378
rect 42642 51326 42654 51378
rect 46946 51326 46958 51378
rect 47010 51326 47022 51378
rect 35422 51314 35474 51326
rect 2382 51266 2434 51278
rect 2382 51202 2434 51214
rect 3166 51266 3218 51278
rect 3166 51202 3218 51214
rect 8430 51266 8482 51278
rect 8430 51202 8482 51214
rect 10334 51266 10386 51278
rect 18958 51266 19010 51278
rect 33630 51266 33682 51278
rect 13906 51214 13918 51266
rect 13970 51214 13982 51266
rect 23202 51214 23214 51266
rect 23266 51214 23278 51266
rect 28914 51214 28926 51266
rect 28978 51214 28990 51266
rect 30258 51214 30270 51266
rect 30322 51214 30334 51266
rect 10334 51202 10386 51214
rect 18958 51202 19010 51214
rect 33630 51202 33682 51214
rect 36318 51266 36370 51278
rect 36318 51202 36370 51214
rect 41694 51266 41746 51278
rect 43934 51266 43986 51278
rect 42690 51214 42702 51266
rect 42754 51214 42766 51266
rect 48066 51214 48078 51266
rect 48130 51214 48142 51266
rect 41694 51202 41746 51214
rect 43934 51202 43986 51214
rect 8878 51154 8930 51166
rect 28814 51154 28866 51166
rect 26786 51102 26798 51154
rect 26850 51102 26862 51154
rect 8878 51090 8930 51102
rect 28814 51090 28866 51102
rect 35534 51154 35586 51166
rect 42914 51102 42926 51154
rect 42978 51102 42990 51154
rect 35534 51090 35586 51102
rect 1344 50986 48608 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 48608 50986
rect 1344 50900 48608 50934
rect 21310 50818 21362 50830
rect 21310 50754 21362 50766
rect 33294 50818 33346 50830
rect 35970 50766 35982 50818
rect 36034 50766 36046 50818
rect 33294 50754 33346 50766
rect 3726 50706 3778 50718
rect 15374 50706 15426 50718
rect 23438 50706 23490 50718
rect 6514 50654 6526 50706
rect 6578 50654 6590 50706
rect 18162 50654 18174 50706
rect 18226 50654 18238 50706
rect 20066 50654 20078 50706
rect 20130 50654 20142 50706
rect 3726 50642 3778 50654
rect 15374 50642 15426 50654
rect 23438 50642 23490 50654
rect 29822 50706 29874 50718
rect 43038 50706 43090 50718
rect 33954 50654 33966 50706
rect 34018 50654 34030 50706
rect 35298 50654 35310 50706
rect 35362 50654 35374 50706
rect 46050 50654 46062 50706
rect 46114 50654 46126 50706
rect 47618 50654 47630 50706
rect 47682 50654 47694 50706
rect 29822 50642 29874 50654
rect 43038 50642 43090 50654
rect 2494 50594 2546 50606
rect 22206 50594 22258 50606
rect 29374 50594 29426 50606
rect 4498 50542 4510 50594
rect 4562 50542 4574 50594
rect 5618 50542 5630 50594
rect 5682 50542 5694 50594
rect 7522 50542 7534 50594
rect 7586 50542 7598 50594
rect 9762 50542 9774 50594
rect 9826 50542 9838 50594
rect 19058 50542 19070 50594
rect 19122 50542 19134 50594
rect 23650 50542 23662 50594
rect 23714 50542 23726 50594
rect 24994 50542 25006 50594
rect 25058 50542 25070 50594
rect 25330 50542 25342 50594
rect 25394 50542 25406 50594
rect 26674 50542 26686 50594
rect 26738 50542 26750 50594
rect 28354 50542 28366 50594
rect 28418 50542 28430 50594
rect 2494 50530 2546 50542
rect 22206 50530 22258 50542
rect 29374 50530 29426 50542
rect 30270 50594 30322 50606
rect 38334 50594 38386 50606
rect 43486 50594 43538 50606
rect 32498 50542 32510 50594
rect 32562 50542 32574 50594
rect 34290 50542 34302 50594
rect 34354 50542 34366 50594
rect 35746 50542 35758 50594
rect 35810 50542 35822 50594
rect 37874 50542 37886 50594
rect 37938 50542 37950 50594
rect 42802 50542 42814 50594
rect 42866 50542 42878 50594
rect 30270 50530 30322 50542
rect 38334 50530 38386 50542
rect 43486 50530 43538 50542
rect 43934 50594 43986 50606
rect 45938 50542 45950 50594
rect 46002 50542 46014 50594
rect 47394 50542 47406 50594
rect 47458 50542 47470 50594
rect 43934 50530 43986 50542
rect 2158 50482 2210 50494
rect 2158 50418 2210 50430
rect 2830 50482 2882 50494
rect 4958 50482 5010 50494
rect 10222 50482 10274 50494
rect 4274 50430 4286 50482
rect 4338 50430 4350 50482
rect 7634 50430 7646 50482
rect 7698 50430 7710 50482
rect 2830 50418 2882 50430
rect 4958 50418 5010 50430
rect 10222 50418 10274 50430
rect 21422 50482 21474 50494
rect 21422 50418 21474 50430
rect 21646 50482 21698 50494
rect 29038 50482 29090 50494
rect 27122 50430 27134 50482
rect 27186 50430 27198 50482
rect 21646 50418 21698 50430
rect 29038 50418 29090 50430
rect 29262 50482 29314 50494
rect 32734 50482 32786 50494
rect 31042 50430 31054 50482
rect 31106 50430 31118 50482
rect 29262 50418 29314 50430
rect 32734 50418 32786 50430
rect 33294 50482 33346 50494
rect 33294 50418 33346 50430
rect 33406 50482 33458 50494
rect 33406 50418 33458 50430
rect 34750 50482 34802 50494
rect 34750 50418 34802 50430
rect 43150 50482 43202 50494
rect 43150 50418 43202 50430
rect 44270 50482 44322 50494
rect 44270 50418 44322 50430
rect 1934 50370 1986 50382
rect 1934 50306 1986 50318
rect 2046 50370 2098 50382
rect 18622 50370 18674 50382
rect 11106 50318 11118 50370
rect 11170 50318 11182 50370
rect 2046 50306 2098 50318
rect 18622 50306 18674 50318
rect 20750 50370 20802 50382
rect 31390 50370 31442 50382
rect 28578 50318 28590 50370
rect 28642 50318 28654 50370
rect 20750 50306 20802 50318
rect 31390 50306 31442 50318
rect 1344 50202 48608 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 48608 50202
rect 1344 50116 48608 50150
rect 3838 50034 3890 50046
rect 12238 50034 12290 50046
rect 17838 50034 17890 50046
rect 2594 49982 2606 50034
rect 2658 49982 2670 50034
rect 7858 49982 7870 50034
rect 7922 49982 7934 50034
rect 13458 49982 13470 50034
rect 13522 49982 13534 50034
rect 15810 49982 15822 50034
rect 15874 49982 15886 50034
rect 3838 49970 3890 49982
rect 12238 49970 12290 49982
rect 16382 49978 16434 49990
rect 11006 49922 11058 49934
rect 6850 49870 6862 49922
rect 6914 49870 6926 49922
rect 8530 49870 8542 49922
rect 8594 49870 8606 49922
rect 11006 49858 11058 49870
rect 12350 49922 12402 49934
rect 12350 49858 12402 49870
rect 16270 49922 16322 49934
rect 17838 49970 17890 49982
rect 17950 50034 18002 50046
rect 18846 50034 18898 50046
rect 18498 49982 18510 50034
rect 18562 49982 18574 50034
rect 17950 49970 18002 49982
rect 18846 49970 18898 49982
rect 19406 50034 19458 50046
rect 26238 50034 26290 50046
rect 25554 49982 25566 50034
rect 25618 49982 25630 50034
rect 35758 50034 35810 50046
rect 41582 50034 41634 50046
rect 19406 49970 19458 49982
rect 26238 49970 26290 49982
rect 33182 49978 33234 49990
rect 16382 49914 16434 49926
rect 19630 49922 19682 49934
rect 25230 49922 25282 49934
rect 16270 49858 16322 49870
rect 21858 49870 21870 49922
rect 21922 49870 21934 49922
rect 19630 49858 19682 49870
rect 25230 49858 25282 49870
rect 25902 49922 25954 49934
rect 25902 49858 25954 49870
rect 26014 49922 26066 49934
rect 26014 49858 26066 49870
rect 26574 49922 26626 49934
rect 39890 49982 39902 50034
rect 39954 49982 39966 50034
rect 35758 49970 35810 49982
rect 41582 49970 41634 49982
rect 33182 49914 33234 49926
rect 33406 49922 33458 49934
rect 26574 49858 26626 49870
rect 33406 49858 33458 49870
rect 34302 49922 34354 49934
rect 34302 49858 34354 49870
rect 35982 49922 36034 49934
rect 35982 49858 36034 49870
rect 39566 49922 39618 49934
rect 39566 49858 39618 49870
rect 40910 49922 40962 49934
rect 40910 49858 40962 49870
rect 41022 49922 41074 49934
rect 47730 49870 47742 49922
rect 47794 49870 47806 49922
rect 41022 49858 41074 49870
rect 2158 49810 2210 49822
rect 2606 49810 2658 49822
rect 11118 49810 11170 49822
rect 2370 49758 2382 49810
rect 2434 49758 2446 49810
rect 2930 49758 2942 49810
rect 2994 49758 3006 49810
rect 6626 49758 6638 49810
rect 6690 49758 6702 49810
rect 7746 49758 7758 49810
rect 7810 49758 7822 49810
rect 2158 49746 2210 49758
rect 2606 49746 2658 49758
rect 11118 49746 11170 49758
rect 13806 49810 13858 49822
rect 13806 49746 13858 49758
rect 15150 49810 15202 49822
rect 19742 49810 19794 49822
rect 15586 49758 15598 49810
rect 15650 49758 15662 49810
rect 19170 49758 19182 49810
rect 19234 49758 19246 49810
rect 15150 49746 15202 49758
rect 19742 49746 19794 49758
rect 20750 49810 20802 49822
rect 20750 49746 20802 49758
rect 21198 49810 21250 49822
rect 23438 49810 23490 49822
rect 22194 49758 22206 49810
rect 22258 49758 22270 49810
rect 21198 49746 21250 49758
rect 23438 49746 23490 49758
rect 26462 49810 26514 49822
rect 26462 49746 26514 49758
rect 26798 49810 26850 49822
rect 26798 49746 26850 49758
rect 27134 49810 27186 49822
rect 31614 49810 31666 49822
rect 27794 49758 27806 49810
rect 27858 49758 27870 49810
rect 27134 49746 27186 49758
rect 31614 49746 31666 49758
rect 33070 49810 33122 49822
rect 33070 49746 33122 49758
rect 33742 49810 33794 49822
rect 33742 49746 33794 49758
rect 34526 49810 34578 49822
rect 34526 49746 34578 49758
rect 36094 49810 36146 49822
rect 43262 49810 43314 49822
rect 40114 49758 40126 49810
rect 40178 49758 40190 49810
rect 43698 49758 43710 49810
rect 43762 49758 43774 49810
rect 46162 49758 46174 49810
rect 46226 49758 46238 49810
rect 47506 49758 47518 49810
rect 47570 49758 47582 49810
rect 36094 49746 36146 49758
rect 43262 49746 43314 49758
rect 1934 49698 1986 49710
rect 4510 49698 4562 49710
rect 3378 49646 3390 49698
rect 3442 49646 3454 49698
rect 1934 49634 1986 49646
rect 4510 49634 4562 49646
rect 4958 49698 5010 49710
rect 4958 49634 5010 49646
rect 5518 49698 5570 49710
rect 5518 49634 5570 49646
rect 10558 49698 10610 49710
rect 10558 49634 10610 49646
rect 14254 49698 14306 49710
rect 14254 49634 14306 49646
rect 14814 49698 14866 49710
rect 23774 49698 23826 49710
rect 20290 49646 20302 49698
rect 20354 49646 20366 49698
rect 14814 49634 14866 49646
rect 23774 49634 23826 49646
rect 24670 49698 24722 49710
rect 31390 49698 31442 49710
rect 28578 49646 28590 49698
rect 28642 49646 28654 49698
rect 30706 49646 30718 49698
rect 30770 49646 30782 49698
rect 24670 49634 24722 49646
rect 31390 49634 31442 49646
rect 36542 49698 36594 49710
rect 36542 49634 36594 49646
rect 44158 49698 44210 49710
rect 45938 49646 45950 49698
rect 46002 49646 46014 49698
rect 44158 49634 44210 49646
rect 11006 49586 11058 49598
rect 11006 49522 11058 49534
rect 12238 49586 12290 49598
rect 16270 49586 16322 49598
rect 14802 49534 14814 49586
rect 14866 49583 14878 49586
rect 15138 49583 15150 49586
rect 14866 49537 15150 49583
rect 14866 49534 14878 49537
rect 15138 49534 15150 49537
rect 15202 49534 15214 49586
rect 12238 49522 12290 49534
rect 16270 49522 16322 49534
rect 18062 49586 18114 49598
rect 18062 49522 18114 49534
rect 31950 49586 32002 49598
rect 31950 49522 32002 49534
rect 34862 49586 34914 49598
rect 34862 49522 34914 49534
rect 41022 49586 41074 49598
rect 41022 49522 41074 49534
rect 1344 49418 48608 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 48608 49418
rect 1344 49332 48608 49366
rect 46050 49198 46062 49250
rect 46114 49198 46126 49250
rect 18398 49138 18450 49150
rect 35870 49138 35922 49150
rect 12674 49086 12686 49138
rect 12738 49086 12750 49138
rect 21746 49086 21758 49138
rect 21810 49086 21822 49138
rect 22642 49086 22654 49138
rect 22706 49086 22718 49138
rect 32050 49086 32062 49138
rect 32114 49086 32126 49138
rect 18398 49074 18450 49086
rect 35870 49074 35922 49086
rect 38894 49138 38946 49150
rect 40798 49138 40850 49150
rect 40450 49086 40462 49138
rect 40514 49086 40526 49138
rect 38894 49074 38946 49086
rect 40798 49074 40850 49086
rect 44270 49138 44322 49150
rect 46386 49086 46398 49138
rect 46450 49086 46462 49138
rect 44270 49074 44322 49086
rect 14142 49026 14194 49038
rect 1698 48974 1710 49026
rect 1762 48974 1774 49026
rect 7186 48974 7198 49026
rect 7250 48974 7262 49026
rect 7634 48974 7646 49026
rect 7698 48974 7710 49026
rect 8978 48974 8990 49026
rect 9042 48974 9054 49026
rect 9874 48974 9886 49026
rect 9938 48974 9950 49026
rect 10546 48974 10558 49026
rect 10610 48974 10622 49026
rect 13570 48974 13582 49026
rect 13634 48974 13646 49026
rect 14142 48962 14194 48974
rect 15038 49026 15090 49038
rect 15038 48962 15090 48974
rect 15710 49026 15762 49038
rect 20750 49026 20802 49038
rect 22206 49026 22258 49038
rect 36094 49026 36146 49038
rect 16146 48974 16158 49026
rect 16210 48974 16222 49026
rect 17042 48974 17054 49026
rect 17106 48974 17118 49026
rect 17714 48974 17726 49026
rect 17778 48974 17790 49026
rect 18610 48974 18622 49026
rect 18674 48974 18686 49026
rect 19058 48974 19070 49026
rect 19122 48974 19134 49026
rect 21410 48974 21422 49026
rect 21474 48974 21486 49026
rect 23314 48974 23326 49026
rect 23378 48974 23390 49026
rect 25218 48974 25230 49026
rect 25282 48974 25294 49026
rect 26898 48974 26910 49026
rect 26962 48974 26974 49026
rect 29138 48974 29150 49026
rect 29202 48974 29214 49026
rect 35074 48974 35086 49026
rect 35138 48974 35150 49026
rect 15710 48962 15762 48974
rect 20750 48962 20802 48974
rect 22206 48962 22258 48974
rect 36094 48962 36146 48974
rect 39230 49026 39282 49038
rect 39230 48962 39282 48974
rect 40014 49026 40066 49038
rect 44158 49026 44210 49038
rect 46958 49026 47010 49038
rect 43810 48974 43822 49026
rect 43874 48974 43886 49026
rect 46162 48974 46174 49026
rect 46226 48974 46238 49026
rect 40014 48962 40066 48974
rect 44158 48962 44210 48974
rect 46958 48962 47010 48974
rect 14478 48914 14530 48926
rect 2482 48862 2494 48914
rect 2546 48862 2558 48914
rect 7522 48862 7534 48914
rect 7586 48862 7598 48914
rect 13794 48862 13806 48914
rect 13858 48862 13870 48914
rect 14478 48850 14530 48862
rect 14702 48914 14754 48926
rect 14702 48850 14754 48862
rect 15262 48914 15314 48926
rect 15262 48850 15314 48862
rect 19518 48914 19570 48926
rect 32398 48914 32450 48926
rect 23202 48862 23214 48914
rect 23266 48862 23278 48914
rect 27346 48862 27358 48914
rect 27410 48862 27422 48914
rect 29922 48862 29934 48914
rect 29986 48862 29998 48914
rect 19518 48850 19570 48862
rect 32398 48850 32450 48862
rect 32958 48914 33010 48926
rect 35534 48914 35586 48926
rect 33618 48862 33630 48914
rect 33682 48862 33694 48914
rect 32958 48850 33010 48862
rect 35534 48850 35586 48862
rect 35646 48914 35698 48926
rect 35646 48850 35698 48862
rect 37998 48914 38050 48926
rect 37998 48850 38050 48862
rect 39566 48914 39618 48926
rect 39566 48850 39618 48862
rect 40126 48914 40178 48926
rect 40126 48850 40178 48862
rect 40910 48914 40962 48926
rect 40910 48850 40962 48862
rect 41582 48914 41634 48926
rect 41582 48850 41634 48862
rect 14254 48802 14306 48814
rect 4722 48750 4734 48802
rect 4786 48750 4798 48802
rect 14254 48738 14306 48750
rect 14814 48802 14866 48814
rect 14814 48738 14866 48750
rect 20190 48802 20242 48814
rect 20190 48738 20242 48750
rect 25790 48802 25842 48814
rect 25790 48738 25842 48750
rect 27806 48802 27858 48814
rect 27806 48738 27858 48750
rect 33294 48802 33346 48814
rect 33294 48738 33346 48750
rect 34862 48802 34914 48814
rect 34862 48738 34914 48750
rect 35310 48802 35362 48814
rect 37662 48802 37714 48814
rect 36418 48750 36430 48802
rect 36482 48750 36494 48802
rect 35310 48738 35362 48750
rect 37662 48738 37714 48750
rect 37886 48802 37938 48814
rect 37886 48738 37938 48750
rect 40350 48802 40402 48814
rect 40350 48738 40402 48750
rect 40462 48802 40514 48814
rect 40462 48738 40514 48750
rect 41134 48802 41186 48814
rect 41134 48738 41186 48750
rect 41358 48802 41410 48814
rect 41358 48738 41410 48750
rect 47742 48802 47794 48814
rect 47742 48738 47794 48750
rect 1344 48634 48608 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 48608 48634
rect 1344 48548 48608 48582
rect 4846 48466 4898 48478
rect 2482 48414 2494 48466
rect 2546 48414 2558 48466
rect 4846 48402 4898 48414
rect 6078 48466 6130 48478
rect 6078 48402 6130 48414
rect 8990 48466 9042 48478
rect 8990 48402 9042 48414
rect 9550 48466 9602 48478
rect 9550 48402 9602 48414
rect 10782 48466 10834 48478
rect 24334 48466 24386 48478
rect 12226 48414 12238 48466
rect 12290 48414 12302 48466
rect 10782 48402 10834 48414
rect 24334 48402 24386 48414
rect 25342 48466 25394 48478
rect 34414 48466 34466 48478
rect 28466 48414 28478 48466
rect 28530 48414 28542 48466
rect 31826 48414 31838 48466
rect 31890 48414 31902 48466
rect 25342 48402 25394 48414
rect 34414 48402 34466 48414
rect 41022 48466 41074 48478
rect 41022 48402 41074 48414
rect 41246 48466 41298 48478
rect 46734 48466 46786 48478
rect 46162 48414 46174 48466
rect 46226 48414 46238 48466
rect 41246 48402 41298 48414
rect 46734 48402 46786 48414
rect 47182 48466 47234 48478
rect 47182 48402 47234 48414
rect 2158 48354 2210 48366
rect 4398 48354 4450 48366
rect 11006 48354 11058 48366
rect 3602 48302 3614 48354
rect 3666 48302 3678 48354
rect 6402 48302 6414 48354
rect 6466 48302 6478 48354
rect 2158 48290 2210 48302
rect 4398 48290 4450 48302
rect 11006 48290 11058 48302
rect 12574 48354 12626 48366
rect 17838 48354 17890 48366
rect 14130 48302 14142 48354
rect 14194 48302 14206 48354
rect 12574 48290 12626 48302
rect 17838 48290 17890 48302
rect 17950 48354 18002 48366
rect 37886 48354 37938 48366
rect 26450 48302 26462 48354
rect 26514 48302 26526 48354
rect 17950 48290 18002 48302
rect 37886 48290 37938 48302
rect 38222 48354 38274 48366
rect 38222 48290 38274 48302
rect 43038 48354 43090 48366
rect 43038 48290 43090 48302
rect 44382 48354 44434 48366
rect 44382 48290 44434 48302
rect 44494 48354 44546 48366
rect 44494 48290 44546 48302
rect 47406 48354 47458 48366
rect 47406 48290 47458 48302
rect 47742 48354 47794 48366
rect 47742 48290 47794 48302
rect 2494 48242 2546 48254
rect 4286 48242 4338 48254
rect 8206 48242 8258 48254
rect 2706 48190 2718 48242
rect 2770 48190 2782 48242
rect 3378 48190 3390 48242
rect 3442 48190 3454 48242
rect 6626 48190 6638 48242
rect 6690 48190 6702 48242
rect 2494 48178 2546 48190
rect 4286 48178 4338 48190
rect 8206 48178 8258 48190
rect 10670 48242 10722 48254
rect 10670 48178 10722 48190
rect 11230 48242 11282 48254
rect 23998 48242 24050 48254
rect 13458 48190 13470 48242
rect 13522 48190 13534 48242
rect 23650 48190 23662 48242
rect 23714 48190 23726 48242
rect 11230 48178 11282 48190
rect 23998 48178 24050 48190
rect 24334 48242 24386 48254
rect 24334 48178 24386 48190
rect 24558 48242 24610 48254
rect 24558 48178 24610 48190
rect 25230 48242 25282 48254
rect 25230 48178 25282 48190
rect 25454 48242 25506 48254
rect 25454 48178 25506 48190
rect 25790 48242 25842 48254
rect 31502 48242 31554 48254
rect 26786 48190 26798 48242
rect 26850 48190 26862 48242
rect 28242 48190 28254 48242
rect 28306 48190 28318 48242
rect 28578 48190 28590 48242
rect 28642 48190 28654 48242
rect 25790 48178 25842 48190
rect 31502 48178 31554 48190
rect 34526 48242 34578 48254
rect 39566 48242 39618 48254
rect 35186 48190 35198 48242
rect 35250 48190 35262 48242
rect 37202 48190 37214 48242
rect 37266 48190 37278 48242
rect 38658 48190 38670 48242
rect 38722 48190 38734 48242
rect 34526 48178 34578 48190
rect 39566 48178 39618 48190
rect 40910 48242 40962 48254
rect 40910 48178 40962 48190
rect 42590 48242 42642 48254
rect 42590 48178 42642 48190
rect 42814 48242 42866 48254
rect 42814 48178 42866 48190
rect 44718 48242 44770 48254
rect 44718 48178 44770 48190
rect 11678 48130 11730 48142
rect 35870 48130 35922 48142
rect 40126 48130 40178 48142
rect 9986 48078 9998 48130
rect 10050 48078 10062 48130
rect 11330 48078 11342 48130
rect 11394 48078 11406 48130
rect 16258 48078 16270 48130
rect 16322 48078 16334 48130
rect 18610 48078 18622 48130
rect 18674 48078 18686 48130
rect 34962 48078 34974 48130
rect 35026 48078 35038 48130
rect 37090 48078 37102 48130
rect 37154 48078 37166 48130
rect 38546 48078 38558 48130
rect 38610 48078 38622 48130
rect 2606 48018 2658 48030
rect 11345 48015 11391 48078
rect 11678 48066 11730 48078
rect 35870 48066 35922 48078
rect 40126 48066 40178 48078
rect 42702 48130 42754 48142
rect 42702 48066 42754 48078
rect 45390 48130 45442 48142
rect 45390 48066 45442 48078
rect 45614 48130 45666 48142
rect 45614 48066 45666 48078
rect 18062 48018 18114 48030
rect 11666 48015 11678 48018
rect 11345 47969 11678 48015
rect 11666 47966 11678 47969
rect 11730 47966 11742 48018
rect 2606 47954 2658 47966
rect 18062 47954 18114 47966
rect 34414 48018 34466 48030
rect 34414 47954 34466 47966
rect 45838 48018 45890 48030
rect 45838 47954 45890 47966
rect 1344 47850 48608 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 48608 47850
rect 1344 47764 48608 47798
rect 2158 47682 2210 47694
rect 2158 47618 2210 47630
rect 2494 47682 2546 47694
rect 2494 47618 2546 47630
rect 20302 47682 20354 47694
rect 20302 47618 20354 47630
rect 32958 47682 33010 47694
rect 43474 47630 43486 47682
rect 43538 47630 43550 47682
rect 32958 47618 33010 47630
rect 3838 47570 3890 47582
rect 3838 47506 3890 47518
rect 19742 47570 19794 47582
rect 19742 47506 19794 47518
rect 23774 47570 23826 47582
rect 23774 47506 23826 47518
rect 25678 47570 25730 47582
rect 25678 47506 25730 47518
rect 26574 47570 26626 47582
rect 34414 47570 34466 47582
rect 33618 47518 33630 47570
rect 33682 47518 33694 47570
rect 41906 47518 41918 47570
rect 41970 47518 41982 47570
rect 26574 47506 26626 47518
rect 34414 47506 34466 47518
rect 2942 47458 2994 47470
rect 2482 47406 2494 47458
rect 2546 47406 2558 47458
rect 2942 47394 2994 47406
rect 4846 47458 4898 47470
rect 20414 47458 20466 47470
rect 24334 47458 24386 47470
rect 7634 47406 7646 47458
rect 7698 47406 7710 47458
rect 10546 47406 10558 47458
rect 10610 47406 10622 47458
rect 10994 47406 11006 47458
rect 11058 47406 11070 47458
rect 14578 47406 14590 47458
rect 14642 47406 14654 47458
rect 15138 47406 15150 47458
rect 15202 47406 15214 47458
rect 21298 47406 21310 47458
rect 21362 47406 21374 47458
rect 4846 47394 4898 47406
rect 20414 47394 20466 47406
rect 22990 47402 23042 47414
rect 4174 47346 4226 47358
rect 4174 47282 4226 47294
rect 4398 47346 4450 47358
rect 4398 47282 4450 47294
rect 4958 47346 5010 47358
rect 24334 47394 24386 47406
rect 24670 47458 24722 47470
rect 24670 47394 24722 47406
rect 25342 47458 25394 47470
rect 34750 47458 34802 47470
rect 33842 47406 33854 47458
rect 33906 47406 33918 47458
rect 25342 47394 25394 47406
rect 34750 47394 34802 47406
rect 34974 47458 35026 47470
rect 34974 47394 35026 47406
rect 37214 47458 37266 47470
rect 37214 47394 37266 47406
rect 37438 47458 37490 47470
rect 37438 47394 37490 47406
rect 40238 47458 40290 47470
rect 41794 47406 41806 47458
rect 41858 47406 41870 47458
rect 42802 47406 42814 47458
rect 42866 47406 42878 47458
rect 40238 47394 40290 47406
rect 7970 47294 7982 47346
rect 8034 47294 8046 47346
rect 14354 47294 14366 47346
rect 14418 47294 14430 47346
rect 15362 47294 15374 47346
rect 15426 47294 15438 47346
rect 22418 47294 22430 47346
rect 22482 47294 22494 47346
rect 22990 47338 23042 47350
rect 23102 47346 23154 47358
rect 4958 47282 5010 47294
rect 23102 47282 23154 47294
rect 25006 47346 25058 47358
rect 25006 47282 25058 47294
rect 25118 47346 25170 47358
rect 25118 47282 25170 47294
rect 32958 47346 33010 47358
rect 32958 47282 33010 47294
rect 33070 47346 33122 47358
rect 33070 47282 33122 47294
rect 37662 47346 37714 47358
rect 37662 47282 37714 47294
rect 39902 47346 39954 47358
rect 39902 47282 39954 47294
rect 40014 47346 40066 47358
rect 40014 47282 40066 47294
rect 40462 47346 40514 47358
rect 40462 47282 40514 47294
rect 4286 47234 4338 47246
rect 4286 47170 4338 47182
rect 5182 47234 5234 47246
rect 20302 47234 20354 47246
rect 7634 47182 7646 47234
rect 7698 47182 7710 47234
rect 5182 47170 5234 47182
rect 20302 47170 20354 47182
rect 23326 47234 23378 47246
rect 23326 47170 23378 47182
rect 24222 47234 24274 47246
rect 24222 47170 24274 47182
rect 24558 47234 24610 47246
rect 24558 47170 24610 47182
rect 26126 47234 26178 47246
rect 26126 47170 26178 47182
rect 34862 47234 34914 47246
rect 34862 47170 34914 47182
rect 35198 47234 35250 47246
rect 35198 47170 35250 47182
rect 37326 47234 37378 47246
rect 37326 47170 37378 47182
rect 38446 47234 38498 47246
rect 39678 47234 39730 47246
rect 38770 47182 38782 47234
rect 38834 47182 38846 47234
rect 38446 47170 38498 47182
rect 39678 47170 39730 47182
rect 40574 47234 40626 47246
rect 40574 47170 40626 47182
rect 40798 47234 40850 47246
rect 40798 47170 40850 47182
rect 1344 47066 48608 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 48608 47066
rect 1344 46980 48608 47014
rect 7534 46898 7586 46910
rect 7534 46834 7586 46846
rect 8318 46898 8370 46910
rect 8318 46834 8370 46846
rect 9886 46898 9938 46910
rect 9886 46834 9938 46846
rect 11678 46898 11730 46910
rect 11678 46834 11730 46846
rect 13470 46898 13522 46910
rect 17502 46898 17554 46910
rect 20638 46898 20690 46910
rect 14130 46846 14142 46898
rect 14194 46846 14206 46898
rect 18050 46846 18062 46898
rect 18114 46846 18126 46898
rect 13470 46834 13522 46846
rect 17502 46834 17554 46846
rect 20638 46834 20690 46846
rect 23326 46898 23378 46910
rect 26238 46898 26290 46910
rect 23874 46846 23886 46898
rect 23938 46846 23950 46898
rect 23326 46834 23378 46846
rect 26238 46834 26290 46846
rect 34974 46898 35026 46910
rect 34974 46834 35026 46846
rect 35086 46898 35138 46910
rect 46622 46898 46674 46910
rect 42578 46846 42590 46898
rect 42642 46846 42654 46898
rect 35086 46834 35138 46846
rect 46622 46834 46674 46846
rect 5406 46786 5458 46798
rect 3490 46734 3502 46786
rect 3554 46734 3566 46786
rect 5406 46722 5458 46734
rect 5742 46786 5794 46798
rect 5742 46722 5794 46734
rect 6078 46786 6130 46798
rect 6078 46722 6130 46734
rect 8878 46786 8930 46798
rect 11230 46786 11282 46798
rect 9538 46734 9550 46786
rect 9602 46734 9614 46786
rect 10546 46734 10558 46786
rect 10610 46734 10622 46786
rect 8878 46722 8930 46734
rect 11230 46722 11282 46734
rect 13806 46786 13858 46798
rect 13806 46722 13858 46734
rect 22990 46786 23042 46798
rect 22990 46722 23042 46734
rect 23102 46786 23154 46798
rect 23102 46722 23154 46734
rect 24222 46786 24274 46798
rect 24222 46722 24274 46734
rect 24334 46786 24386 46798
rect 24334 46722 24386 46734
rect 30718 46786 30770 46798
rect 30718 46722 30770 46734
rect 33742 46786 33794 46798
rect 33742 46722 33794 46734
rect 33854 46786 33906 46798
rect 33854 46722 33906 46734
rect 44494 46786 44546 46798
rect 44494 46722 44546 46734
rect 10222 46674 10274 46686
rect 3826 46622 3838 46674
rect 3890 46622 3902 46674
rect 4834 46622 4846 46674
rect 4898 46622 4910 46674
rect 10222 46610 10274 46622
rect 17390 46674 17442 46686
rect 20750 46674 20802 46686
rect 18274 46622 18286 46674
rect 18338 46622 18350 46674
rect 17390 46610 17442 46622
rect 20750 46610 20802 46622
rect 23550 46674 23602 46686
rect 23550 46610 23602 46622
rect 24558 46674 24610 46686
rect 24558 46610 24610 46622
rect 25118 46674 25170 46686
rect 25118 46610 25170 46622
rect 25566 46674 25618 46686
rect 25566 46610 25618 46622
rect 25678 46674 25730 46686
rect 25678 46610 25730 46622
rect 26126 46674 26178 46686
rect 34414 46674 34466 46686
rect 42254 46674 42306 46686
rect 26786 46622 26798 46674
rect 26850 46622 26862 46674
rect 34738 46622 34750 46674
rect 34802 46622 34814 46674
rect 43810 46622 43822 46674
rect 43874 46622 43886 46674
rect 46946 46622 46958 46674
rect 47010 46622 47022 46674
rect 26126 46610 26178 46622
rect 34414 46610 34466 46622
rect 42254 46610 42306 46622
rect 7982 46562 8034 46574
rect 7982 46498 8034 46510
rect 18958 46562 19010 46574
rect 18958 46498 19010 46510
rect 21198 46562 21250 46574
rect 21198 46498 21250 46510
rect 22206 46562 22258 46574
rect 22206 46498 22258 46510
rect 22654 46562 22706 46574
rect 22654 46498 22706 46510
rect 25342 46562 25394 46574
rect 31278 46562 31330 46574
rect 27458 46510 27470 46562
rect 27522 46510 27534 46562
rect 29586 46510 29598 46562
rect 29650 46510 29662 46562
rect 25342 46498 25394 46510
rect 31278 46498 31330 46510
rect 38110 46562 38162 46574
rect 38110 46498 38162 46510
rect 40126 46562 40178 46574
rect 40126 46498 40178 46510
rect 42030 46562 42082 46574
rect 44034 46510 44046 46562
rect 44098 46510 44110 46562
rect 48066 46510 48078 46562
rect 48130 46510 48142 46562
rect 42030 46498 42082 46510
rect 17502 46450 17554 46462
rect 11218 46398 11230 46450
rect 11282 46447 11294 46450
rect 11666 46447 11678 46450
rect 11282 46401 11678 46447
rect 11282 46398 11294 46401
rect 11666 46398 11678 46401
rect 11730 46398 11742 46450
rect 17502 46386 17554 46398
rect 26238 46450 26290 46462
rect 26238 46386 26290 46398
rect 30606 46450 30658 46462
rect 30606 46386 30658 46398
rect 33742 46450 33794 46462
rect 33742 46386 33794 46398
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 17502 46114 17554 46126
rect 42478 46114 42530 46126
rect 18498 46062 18510 46114
rect 18562 46062 18574 46114
rect 17502 46050 17554 46062
rect 42478 46050 42530 46062
rect 42814 46114 42866 46126
rect 42814 46050 42866 46062
rect 13582 46002 13634 46014
rect 6402 45950 6414 46002
rect 6466 45950 6478 46002
rect 8530 45950 8542 46002
rect 8594 45950 8606 46002
rect 11554 45950 11566 46002
rect 11618 45950 11630 46002
rect 13582 45938 13634 45950
rect 17166 46002 17218 46014
rect 17166 45938 17218 45950
rect 24894 46002 24946 46014
rect 24894 45938 24946 45950
rect 39902 46002 39954 46014
rect 39902 45938 39954 45950
rect 43710 46002 43762 46014
rect 43710 45938 43762 45950
rect 45166 46002 45218 46014
rect 45166 45938 45218 45950
rect 4398 45890 4450 45902
rect 4398 45826 4450 45838
rect 4734 45890 4786 45902
rect 4734 45826 4786 45838
rect 4958 45890 5010 45902
rect 14142 45890 14194 45902
rect 5730 45838 5742 45890
rect 5794 45838 5806 45890
rect 4958 45826 5010 45838
rect 14142 45826 14194 45838
rect 14814 45890 14866 45902
rect 14814 45826 14866 45838
rect 15374 45890 15426 45902
rect 15374 45826 15426 45838
rect 15822 45890 15874 45902
rect 15822 45826 15874 45838
rect 15934 45890 15986 45902
rect 17838 45890 17890 45902
rect 16594 45838 16606 45890
rect 16658 45838 16670 45890
rect 15934 45826 15986 45838
rect 17838 45826 17890 45838
rect 18622 45890 18674 45902
rect 22318 45890 22370 45902
rect 18946 45838 18958 45890
rect 19010 45838 19022 45890
rect 20626 45838 20638 45890
rect 20690 45838 20702 45890
rect 18622 45826 18674 45838
rect 22318 45826 22370 45838
rect 22878 45890 22930 45902
rect 22878 45826 22930 45838
rect 23886 45890 23938 45902
rect 23886 45826 23938 45838
rect 24446 45890 24498 45902
rect 24446 45826 24498 45838
rect 26910 45890 26962 45902
rect 40798 45890 40850 45902
rect 31378 45838 31390 45890
rect 31442 45838 31454 45890
rect 26910 45826 26962 45838
rect 40798 45826 40850 45838
rect 42254 45890 42306 45902
rect 42254 45826 42306 45838
rect 44046 45890 44098 45902
rect 44046 45826 44098 45838
rect 9550 45778 9602 45790
rect 9550 45714 9602 45726
rect 9886 45778 9938 45790
rect 9886 45714 9938 45726
rect 10222 45778 10274 45790
rect 11006 45778 11058 45790
rect 10546 45726 10558 45778
rect 10610 45726 10622 45778
rect 10222 45714 10274 45726
rect 11006 45714 11058 45726
rect 11230 45778 11282 45790
rect 11230 45714 11282 45726
rect 11678 45778 11730 45790
rect 11678 45714 11730 45726
rect 11902 45778 11954 45790
rect 11902 45714 11954 45726
rect 14478 45778 14530 45790
rect 14478 45714 14530 45726
rect 18062 45778 18114 45790
rect 23214 45778 23266 45790
rect 20738 45726 20750 45778
rect 20802 45726 20814 45778
rect 21522 45726 21534 45778
rect 21586 45726 21598 45778
rect 21858 45726 21870 45778
rect 21922 45726 21934 45778
rect 18062 45714 18114 45726
rect 23214 45714 23266 45726
rect 23438 45778 23490 45790
rect 23438 45714 23490 45726
rect 26238 45778 26290 45790
rect 26238 45714 26290 45726
rect 26574 45778 26626 45790
rect 30830 45778 30882 45790
rect 30258 45726 30270 45778
rect 30322 45726 30334 45778
rect 26574 45714 26626 45726
rect 30830 45714 30882 45726
rect 31054 45778 31106 45790
rect 40462 45778 40514 45790
rect 31490 45726 31502 45778
rect 31554 45726 31566 45778
rect 32050 45726 32062 45778
rect 32114 45726 32126 45778
rect 31054 45714 31106 45726
rect 40462 45714 40514 45726
rect 40574 45778 40626 45790
rect 40574 45714 40626 45726
rect 44158 45778 44210 45790
rect 45602 45726 45614 45778
rect 45666 45726 45678 45778
rect 46946 45726 46958 45778
rect 47010 45726 47022 45778
rect 44158 45714 44210 45726
rect 4846 45666 4898 45678
rect 4846 45602 4898 45614
rect 9326 45666 9378 45678
rect 9326 45602 9378 45614
rect 11118 45666 11170 45678
rect 11118 45602 11170 45614
rect 12350 45666 12402 45678
rect 15598 45666 15650 45678
rect 19630 45666 19682 45678
rect 23326 45666 23378 45678
rect 15138 45614 15150 45666
rect 15202 45614 15214 45666
rect 16370 45614 16382 45666
rect 16434 45614 16446 45666
rect 20178 45614 20190 45666
rect 20242 45614 20254 45666
rect 21970 45614 21982 45666
rect 22034 45614 22046 45666
rect 12350 45602 12402 45614
rect 15598 45602 15650 45614
rect 19630 45602 19682 45614
rect 23326 45602 23378 45614
rect 29598 45666 29650 45678
rect 29598 45602 29650 45614
rect 29934 45666 29986 45678
rect 29934 45602 29986 45614
rect 30942 45666 30994 45678
rect 30942 45602 30994 45614
rect 41246 45666 41298 45678
rect 41246 45602 41298 45614
rect 44382 45666 44434 45678
rect 46834 45614 46846 45666
rect 46898 45614 46910 45666
rect 44382 45602 44434 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 1934 45330 1986 45342
rect 14590 45330 14642 45342
rect 2146 45278 2158 45330
rect 2210 45278 2222 45330
rect 1934 45266 1986 45278
rect 14590 45266 14642 45278
rect 15262 45330 15314 45342
rect 15262 45266 15314 45278
rect 15374 45330 15426 45342
rect 15374 45266 15426 45278
rect 15598 45330 15650 45342
rect 15598 45266 15650 45278
rect 18622 45330 18674 45342
rect 18622 45266 18674 45278
rect 29934 45330 29986 45342
rect 29934 45266 29986 45278
rect 41022 45330 41074 45342
rect 41022 45266 41074 45278
rect 41470 45330 41522 45342
rect 41470 45266 41522 45278
rect 3166 45218 3218 45230
rect 13694 45218 13746 45230
rect 20414 45218 20466 45230
rect 12226 45166 12238 45218
rect 12290 45166 12302 45218
rect 18946 45166 18958 45218
rect 19010 45166 19022 45218
rect 3166 45154 3218 45166
rect 13694 45154 13746 45166
rect 20414 45154 20466 45166
rect 20750 45218 20802 45230
rect 25902 45218 25954 45230
rect 32062 45218 32114 45230
rect 23650 45166 23662 45218
rect 23714 45166 23726 45218
rect 27122 45166 27134 45218
rect 27186 45166 27198 45218
rect 20750 45154 20802 45166
rect 25902 45154 25954 45166
rect 32062 45154 32114 45166
rect 35198 45218 35250 45230
rect 35198 45154 35250 45166
rect 35646 45218 35698 45230
rect 35646 45154 35698 45166
rect 35870 45218 35922 45230
rect 35870 45154 35922 45166
rect 36206 45218 36258 45230
rect 36206 45154 36258 45166
rect 36318 45218 36370 45230
rect 36318 45154 36370 45166
rect 36766 45218 36818 45230
rect 39902 45218 39954 45230
rect 36766 45154 36818 45166
rect 36878 45162 36930 45174
rect 38322 45166 38334 45218
rect 38386 45166 38398 45218
rect 2494 45106 2546 45118
rect 7870 45106 7922 45118
rect 2818 45054 2830 45106
rect 2882 45054 2894 45106
rect 2494 45042 2546 45054
rect 7870 45042 7922 45054
rect 8318 45106 8370 45118
rect 15710 45106 15762 45118
rect 13010 45054 13022 45106
rect 13074 45054 13086 45106
rect 13346 45054 13358 45106
rect 13410 45054 13422 45106
rect 8318 45042 8370 45054
rect 15710 45042 15762 45054
rect 17502 45106 17554 45118
rect 17502 45042 17554 45054
rect 17838 45106 17890 45118
rect 23326 45106 23378 45118
rect 26014 45106 26066 45118
rect 29822 45106 29874 45118
rect 21186 45054 21198 45106
rect 21250 45054 21262 45106
rect 25218 45054 25230 45106
rect 25282 45054 25294 45106
rect 25778 45054 25790 45106
rect 25842 45054 25854 45106
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 17838 45042 17890 45054
rect 23326 45042 23378 45054
rect 26014 45042 26066 45054
rect 29822 45042 29874 45054
rect 30158 45106 30210 45118
rect 31838 45106 31890 45118
rect 35534 45106 35586 45118
rect 30818 45054 30830 45106
rect 30882 45054 30894 45106
rect 34738 45054 34750 45106
rect 34802 45054 34814 45106
rect 30158 45042 30210 45054
rect 31838 45042 31890 45054
rect 35534 45042 35586 45054
rect 36542 45106 36594 45118
rect 39902 45154 39954 45166
rect 40238 45218 40290 45230
rect 40238 45154 40290 45166
rect 42030 45218 42082 45230
rect 42030 45154 42082 45166
rect 44718 45218 44770 45230
rect 44718 45154 44770 45166
rect 44830 45218 44882 45230
rect 44830 45154 44882 45166
rect 36878 45098 36930 45110
rect 38670 45106 38722 45118
rect 36542 45042 36594 45054
rect 38670 45042 38722 45054
rect 41358 45106 41410 45118
rect 41358 45042 41410 45054
rect 45054 45106 45106 45118
rect 45054 45042 45106 45054
rect 3614 44994 3666 45006
rect 3614 44930 3666 44942
rect 7534 44994 7586 45006
rect 7534 44930 7586 44942
rect 8990 44994 9042 45006
rect 8990 44930 9042 44942
rect 9662 44994 9714 45006
rect 14142 44994 14194 45006
rect 10098 44942 10110 44994
rect 10162 44942 10174 44994
rect 9662 44930 9714 44942
rect 14142 44930 14194 44942
rect 17726 44994 17778 45006
rect 19630 44994 19682 45006
rect 19170 44942 19182 44994
rect 19234 44942 19246 44994
rect 17726 44930 17778 44942
rect 2830 44882 2882 44894
rect 2830 44818 2882 44830
rect 13358 44882 13410 44894
rect 19185 44879 19231 44942
rect 19630 44930 19682 44942
rect 21758 44994 21810 45006
rect 21758 44930 21810 44942
rect 22206 44994 22258 45006
rect 22206 44930 22258 44942
rect 24670 44994 24722 45006
rect 31950 44994 32002 45006
rect 37998 44994 38050 45006
rect 29250 44942 29262 44994
rect 29314 44942 29326 44994
rect 30706 44942 30718 44994
rect 30770 44942 30782 44994
rect 34290 44942 34302 44994
rect 34354 44942 34366 44994
rect 24670 44930 24722 44942
rect 31950 44930 32002 44942
rect 37998 44930 38050 44942
rect 39566 44994 39618 45006
rect 39566 44930 39618 44942
rect 45726 44994 45778 45006
rect 45726 44930 45778 44942
rect 19854 44882 19906 44894
rect 19506 44879 19518 44882
rect 19185 44833 19518 44879
rect 19506 44830 19518 44833
rect 19570 44830 19582 44882
rect 13358 44818 13410 44830
rect 19854 44818 19906 44830
rect 20190 44882 20242 44894
rect 36206 44882 36258 44894
rect 24434 44830 24446 44882
rect 24498 44879 24510 44882
rect 24658 44879 24670 44882
rect 24498 44833 24670 44879
rect 24498 44830 24510 44833
rect 24658 44830 24670 44833
rect 24722 44830 24734 44882
rect 25442 44830 25454 44882
rect 25506 44830 25518 44882
rect 31042 44830 31054 44882
rect 31106 44830 31118 44882
rect 20190 44818 20242 44830
rect 36206 44818 36258 44830
rect 41470 44882 41522 44894
rect 41470 44818 41522 44830
rect 45838 44882 45890 44894
rect 45838 44818 45890 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 13694 44546 13746 44558
rect 2706 44494 2718 44546
rect 2770 44494 2782 44546
rect 13694 44482 13746 44494
rect 20078 44546 20130 44558
rect 20078 44482 20130 44494
rect 23102 44546 23154 44558
rect 46622 44546 46674 44558
rect 25106 44494 25118 44546
rect 25170 44494 25182 44546
rect 43250 44494 43262 44546
rect 43314 44494 43326 44546
rect 23102 44482 23154 44494
rect 46622 44482 46674 44494
rect 5742 44434 5794 44446
rect 5742 44370 5794 44382
rect 6302 44434 6354 44446
rect 15934 44434 15986 44446
rect 14018 44382 14030 44434
rect 14082 44382 14094 44434
rect 6302 44370 6354 44382
rect 15934 44370 15986 44382
rect 18062 44434 18114 44446
rect 23550 44434 23602 44446
rect 20402 44382 20414 44434
rect 20466 44382 20478 44434
rect 18062 44370 18114 44382
rect 23550 44370 23602 44382
rect 24670 44434 24722 44446
rect 32398 44434 32450 44446
rect 45950 44434 46002 44446
rect 31490 44382 31502 44434
rect 31554 44382 31566 44434
rect 34066 44382 34078 44434
rect 34130 44382 34142 44434
rect 42690 44382 42702 44434
rect 42754 44382 42766 44434
rect 24670 44370 24722 44382
rect 32398 44370 32450 44382
rect 45950 44370 46002 44382
rect 2158 44322 2210 44334
rect 16382 44322 16434 44334
rect 17838 44322 17890 44334
rect 2930 44270 2942 44322
rect 2994 44270 3006 44322
rect 12898 44270 12910 44322
rect 12962 44270 12974 44322
rect 14578 44270 14590 44322
rect 14642 44270 14654 44322
rect 16818 44270 16830 44322
rect 16882 44270 16894 44322
rect 2158 44258 2210 44270
rect 16382 44258 16434 44270
rect 17838 44258 17890 44270
rect 22094 44322 22146 44334
rect 22094 44258 22146 44270
rect 23886 44322 23938 44334
rect 25342 44322 25394 44334
rect 24882 44270 24894 44322
rect 24946 44270 24958 44322
rect 23886 44258 23938 44270
rect 25342 44258 25394 44270
rect 30046 44322 30098 44334
rect 30046 44258 30098 44270
rect 30718 44322 30770 44334
rect 34974 44322 35026 44334
rect 30930 44270 30942 44322
rect 30994 44270 31006 44322
rect 31826 44270 31838 44322
rect 31890 44270 31902 44322
rect 34402 44270 34414 44322
rect 34466 44270 34478 44322
rect 30718 44258 30770 44270
rect 34974 44258 35026 44270
rect 37102 44322 37154 44334
rect 37998 44322 38050 44334
rect 37314 44270 37326 44322
rect 37378 44270 37390 44322
rect 37102 44258 37154 44270
rect 37998 44258 38050 44270
rect 38446 44322 38498 44334
rect 39678 44322 39730 44334
rect 38658 44270 38670 44322
rect 38722 44270 38734 44322
rect 42578 44270 42590 44322
rect 42642 44270 42654 44322
rect 47058 44270 47070 44322
rect 47122 44270 47134 44322
rect 38446 44258 38498 44270
rect 39678 44258 39730 44270
rect 3950 44210 4002 44222
rect 2370 44158 2382 44210
rect 2434 44158 2446 44210
rect 3266 44158 3278 44210
rect 3330 44158 3342 44210
rect 3950 44146 4002 44158
rect 4174 44210 4226 44222
rect 4174 44146 4226 44158
rect 6526 44210 6578 44222
rect 6526 44146 6578 44158
rect 7198 44210 7250 44222
rect 13918 44210 13970 44222
rect 7858 44158 7870 44210
rect 7922 44158 7934 44210
rect 7198 44146 7250 44158
rect 13918 44146 13970 44158
rect 14366 44210 14418 44222
rect 14366 44146 14418 44158
rect 16270 44210 16322 44222
rect 22766 44210 22818 44222
rect 17042 44158 17054 44210
rect 17106 44158 17118 44210
rect 22418 44158 22430 44210
rect 22482 44158 22494 44210
rect 16270 44146 16322 44158
rect 22766 44146 22818 44158
rect 23998 44210 24050 44222
rect 23998 44146 24050 44158
rect 25678 44210 25730 44222
rect 25678 44146 25730 44158
rect 29710 44210 29762 44222
rect 29710 44146 29762 44158
rect 31054 44210 31106 44222
rect 31054 44146 31106 44158
rect 39342 44210 39394 44222
rect 41022 44210 41074 44222
rect 40002 44158 40014 44210
rect 40066 44158 40078 44210
rect 40674 44158 40686 44210
rect 40738 44158 40750 44210
rect 39342 44146 39394 44158
rect 41022 44146 41074 44158
rect 41134 44210 41186 44222
rect 41134 44146 41186 44158
rect 41582 44210 41634 44222
rect 41582 44146 41634 44158
rect 41694 44210 41746 44222
rect 41694 44146 41746 44158
rect 46286 44210 46338 44222
rect 46286 44146 46338 44158
rect 46510 44210 46562 44222
rect 46510 44146 46562 44158
rect 3614 44098 3666 44110
rect 2482 44046 2494 44098
rect 2546 44046 2558 44098
rect 3614 44034 3666 44046
rect 4062 44098 4114 44110
rect 4062 44034 4114 44046
rect 4734 44098 4786 44110
rect 4734 44034 4786 44046
rect 6638 44098 6690 44110
rect 6638 44034 6690 44046
rect 6862 44098 6914 44110
rect 6862 44034 6914 44046
rect 7086 44098 7138 44110
rect 7086 44034 7138 44046
rect 15262 44098 15314 44110
rect 15262 44034 15314 44046
rect 16046 44098 16098 44110
rect 20302 44098 20354 44110
rect 17490 44046 17502 44098
rect 17554 44046 17566 44098
rect 16046 44034 16098 44046
rect 20302 44034 20354 44046
rect 21758 44098 21810 44110
rect 21758 44034 21810 44046
rect 22990 44098 23042 44110
rect 22990 44034 23042 44046
rect 24222 44098 24274 44110
rect 24222 44034 24274 44046
rect 25566 44098 25618 44110
rect 25566 44034 25618 44046
rect 26238 44098 26290 44110
rect 26238 44034 26290 44046
rect 29374 44098 29426 44110
rect 29374 44034 29426 44046
rect 29822 44098 29874 44110
rect 29822 44034 29874 44046
rect 40350 44098 40402 44110
rect 40350 44034 40402 44046
rect 41358 44098 41410 44110
rect 41358 44034 41410 44046
rect 41918 44098 41970 44110
rect 41918 44034 41970 44046
rect 47742 44098 47794 44110
rect 47742 44034 47794 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 3726 43762 3778 43774
rect 3726 43698 3778 43710
rect 10894 43762 10946 43774
rect 14478 43762 14530 43774
rect 12450 43710 12462 43762
rect 12514 43710 12526 43762
rect 10894 43698 10946 43710
rect 14478 43698 14530 43710
rect 18286 43762 18338 43774
rect 39342 43762 39394 43774
rect 41022 43762 41074 43774
rect 19506 43710 19518 43762
rect 19570 43710 19582 43762
rect 20290 43710 20302 43762
rect 20354 43710 20366 43762
rect 39890 43710 39902 43762
rect 39954 43710 39966 43762
rect 18286 43698 18338 43710
rect 39342 43698 39394 43710
rect 41022 43698 41074 43710
rect 2158 43650 2210 43662
rect 2158 43586 2210 43598
rect 5294 43650 5346 43662
rect 5294 43586 5346 43598
rect 5406 43650 5458 43662
rect 6638 43650 6690 43662
rect 5842 43598 5854 43650
rect 5906 43598 5918 43650
rect 5406 43586 5458 43598
rect 6638 43586 6690 43598
rect 6862 43650 6914 43662
rect 15374 43650 15426 43662
rect 8866 43598 8878 43650
rect 8930 43598 8942 43650
rect 10210 43598 10222 43650
rect 10274 43598 10286 43650
rect 11442 43598 11454 43650
rect 11506 43598 11518 43650
rect 6862 43586 6914 43598
rect 15374 43586 15426 43598
rect 15598 43650 15650 43662
rect 15598 43586 15650 43598
rect 16382 43650 16434 43662
rect 16382 43586 16434 43598
rect 16606 43650 16658 43662
rect 16606 43586 16658 43598
rect 16718 43650 16770 43662
rect 16718 43586 16770 43598
rect 18510 43650 18562 43662
rect 20862 43650 20914 43662
rect 23774 43650 23826 43662
rect 20178 43598 20190 43650
rect 20242 43598 20254 43650
rect 22082 43598 22094 43650
rect 22146 43598 22158 43650
rect 18510 43586 18562 43598
rect 20862 43586 20914 43598
rect 23774 43586 23826 43598
rect 23998 43650 24050 43662
rect 23998 43586 24050 43598
rect 24110 43650 24162 43662
rect 24110 43586 24162 43598
rect 42478 43650 42530 43662
rect 42478 43586 42530 43598
rect 42814 43650 42866 43662
rect 42814 43586 42866 43598
rect 2606 43538 2658 43550
rect 4510 43538 4562 43550
rect 2370 43486 2382 43538
rect 2434 43486 2446 43538
rect 2930 43486 2942 43538
rect 2994 43486 3006 43538
rect 2606 43474 2658 43486
rect 4510 43474 4562 43486
rect 4622 43538 4674 43550
rect 4622 43474 4674 43486
rect 4958 43538 5010 43550
rect 4958 43474 5010 43486
rect 5630 43538 5682 43550
rect 5630 43474 5682 43486
rect 6190 43538 6242 43550
rect 6190 43474 6242 43486
rect 7086 43538 7138 43550
rect 7086 43474 7138 43486
rect 7646 43538 7698 43550
rect 7646 43474 7698 43486
rect 9550 43538 9602 43550
rect 10558 43538 10610 43550
rect 11230 43538 11282 43550
rect 9874 43486 9886 43538
rect 9938 43486 9950 43538
rect 10994 43486 11006 43538
rect 11058 43486 11070 43538
rect 9550 43474 9602 43486
rect 10558 43474 10610 43486
rect 11230 43474 11282 43486
rect 11678 43538 11730 43550
rect 12350 43538 12402 43550
rect 12798 43538 12850 43550
rect 12002 43486 12014 43538
rect 12066 43486 12078 43538
rect 12562 43486 12574 43538
rect 12626 43486 12638 43538
rect 11678 43474 11730 43486
rect 12350 43474 12402 43486
rect 12798 43474 12850 43486
rect 13694 43538 13746 43550
rect 13694 43474 13746 43486
rect 14030 43538 14082 43550
rect 14030 43474 14082 43486
rect 14142 43538 14194 43550
rect 15934 43538 15986 43550
rect 14242 43486 14254 43538
rect 14306 43486 14318 43538
rect 14142 43474 14194 43486
rect 15934 43474 15986 43486
rect 16270 43538 16322 43550
rect 16270 43474 16322 43486
rect 18622 43538 18674 43550
rect 24334 43538 24386 43550
rect 19842 43486 19854 43538
rect 19906 43486 19918 43538
rect 21298 43486 21310 43538
rect 21362 43486 21374 43538
rect 21858 43486 21870 43538
rect 21922 43486 21934 43538
rect 18622 43474 18674 43486
rect 24334 43474 24386 43486
rect 25230 43538 25282 43550
rect 25230 43474 25282 43486
rect 25566 43538 25618 43550
rect 25566 43474 25618 43486
rect 25790 43538 25842 43550
rect 37886 43538 37938 43550
rect 26450 43486 26462 43538
rect 26514 43486 26526 43538
rect 25790 43474 25842 43486
rect 37886 43474 37938 43486
rect 38110 43538 38162 43550
rect 41582 43538 41634 43550
rect 43038 43538 43090 43550
rect 46510 43538 46562 43550
rect 40114 43486 40126 43538
rect 40178 43486 40190 43538
rect 42018 43486 42030 43538
rect 42082 43486 42094 43538
rect 45938 43486 45950 43538
rect 46002 43486 46014 43538
rect 38110 43474 38162 43486
rect 41582 43474 41634 43486
rect 43038 43474 43090 43486
rect 46510 43474 46562 43486
rect 46622 43538 46674 43550
rect 46622 43474 46674 43486
rect 46846 43538 46898 43550
rect 46846 43474 46898 43486
rect 47182 43538 47234 43550
rect 47182 43474 47234 43486
rect 47406 43538 47458 43550
rect 47406 43474 47458 43486
rect 2270 43426 2322 43438
rect 2270 43362 2322 43374
rect 4846 43426 4898 43438
rect 4846 43362 4898 43374
rect 6750 43426 6802 43438
rect 6750 43362 6802 43374
rect 7534 43426 7586 43438
rect 13246 43426 13298 43438
rect 8530 43374 8542 43426
rect 8594 43374 8606 43426
rect 7534 43362 7586 43374
rect 13246 43362 13298 43374
rect 16046 43426 16098 43438
rect 16046 43362 16098 43374
rect 18174 43426 18226 43438
rect 18174 43362 18226 43374
rect 18958 43426 19010 43438
rect 18958 43362 19010 43374
rect 25342 43426 25394 43438
rect 45278 43426 45330 43438
rect 27234 43374 27246 43426
rect 27298 43374 27310 43426
rect 29362 43374 29374 43426
rect 29426 43374 29438 43426
rect 25342 43362 25394 43374
rect 45278 43362 45330 43374
rect 47070 43426 47122 43438
rect 47070 43362 47122 43374
rect 9886 43314 9938 43326
rect 9886 43250 9938 43262
rect 19182 43314 19234 43326
rect 43374 43314 43426 43326
rect 38434 43262 38446 43314
rect 38498 43262 38510 43314
rect 19182 43250 19234 43262
rect 43374 43250 43426 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 6638 42978 6690 42990
rect 6638 42914 6690 42926
rect 7086 42978 7138 42990
rect 9886 42978 9938 42990
rect 8642 42926 8654 42978
rect 8706 42926 8718 42978
rect 7086 42914 7138 42926
rect 9886 42914 9938 42926
rect 11006 42978 11058 42990
rect 27022 42978 27074 42990
rect 12562 42926 12574 42978
rect 12626 42975 12638 42978
rect 13010 42975 13022 42978
rect 12626 42929 13022 42975
rect 12626 42926 12638 42929
rect 13010 42926 13022 42929
rect 13074 42926 13086 42978
rect 11006 42914 11058 42926
rect 27022 42914 27074 42926
rect 33070 42978 33122 42990
rect 33070 42914 33122 42926
rect 42590 42978 42642 42990
rect 42590 42914 42642 42926
rect 12798 42866 12850 42878
rect 8754 42814 8766 42866
rect 8818 42814 8830 42866
rect 12798 42802 12850 42814
rect 15038 42866 15090 42878
rect 15038 42802 15090 42814
rect 16382 42866 16434 42878
rect 16382 42802 16434 42814
rect 34414 42866 34466 42878
rect 41246 42866 41298 42878
rect 37538 42814 37550 42866
rect 37602 42814 37614 42866
rect 38098 42814 38110 42866
rect 38162 42814 38174 42866
rect 34414 42802 34466 42814
rect 41246 42802 41298 42814
rect 41918 42866 41970 42878
rect 41918 42802 41970 42814
rect 43038 42866 43090 42878
rect 46846 42866 46898 42878
rect 46386 42814 46398 42866
rect 46450 42814 46462 42866
rect 43038 42802 43090 42814
rect 46846 42802 46898 42814
rect 5630 42754 5682 42766
rect 3714 42702 3726 42754
rect 3778 42702 3790 42754
rect 4386 42702 4398 42754
rect 4450 42702 4462 42754
rect 5630 42690 5682 42702
rect 7310 42754 7362 42766
rect 10334 42754 10386 42766
rect 11454 42754 11506 42766
rect 9538 42702 9550 42754
rect 9602 42702 9614 42754
rect 10882 42702 10894 42754
rect 10946 42702 10958 42754
rect 11218 42702 11230 42754
rect 11282 42702 11294 42754
rect 7310 42690 7362 42702
rect 10334 42690 10386 42702
rect 11454 42690 11506 42702
rect 13806 42754 13858 42766
rect 13806 42690 13858 42702
rect 20414 42754 20466 42766
rect 26910 42754 26962 42766
rect 22418 42702 22430 42754
rect 22482 42702 22494 42754
rect 24098 42702 24110 42754
rect 24162 42702 24174 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 20414 42690 20466 42702
rect 26910 42690 26962 42702
rect 27694 42754 27746 42766
rect 27694 42690 27746 42702
rect 33294 42754 33346 42766
rect 43262 42754 43314 42766
rect 37426 42702 37438 42754
rect 37490 42702 37502 42754
rect 38434 42702 38446 42754
rect 38498 42702 38510 42754
rect 46162 42702 46174 42754
rect 46226 42702 46238 42754
rect 33294 42690 33346 42702
rect 43262 42690 43314 42702
rect 6526 42642 6578 42654
rect 3154 42590 3166 42642
rect 3218 42590 3230 42642
rect 6526 42578 6578 42590
rect 6974 42642 7026 42654
rect 6974 42578 7026 42590
rect 7758 42642 7810 42654
rect 13470 42642 13522 42654
rect 9090 42590 9102 42642
rect 9154 42590 9166 42642
rect 10098 42590 10110 42642
rect 10162 42590 10174 42642
rect 7758 42578 7810 42590
rect 13470 42578 13522 42590
rect 20078 42642 20130 42654
rect 20078 42578 20130 42590
rect 20302 42642 20354 42654
rect 27022 42642 27074 42654
rect 23202 42590 23214 42642
rect 23266 42590 23278 42642
rect 25666 42590 25678 42642
rect 25730 42590 25742 42642
rect 20302 42578 20354 42590
rect 27022 42578 27074 42590
rect 33966 42642 34018 42654
rect 42702 42642 42754 42654
rect 37202 42590 37214 42642
rect 37266 42590 37278 42642
rect 33966 42578 34018 42590
rect 42702 42578 42754 42590
rect 5742 42530 5794 42542
rect 4946 42478 4958 42530
rect 5010 42478 5022 42530
rect 5742 42466 5794 42478
rect 5854 42530 5906 42542
rect 5854 42466 5906 42478
rect 9550 42530 9602 42542
rect 9550 42466 9602 42478
rect 11342 42530 11394 42542
rect 11342 42466 11394 42478
rect 11902 42530 11954 42542
rect 11902 42466 11954 42478
rect 12350 42530 12402 42542
rect 12350 42466 12402 42478
rect 19742 42530 19794 42542
rect 19742 42466 19794 42478
rect 21422 42530 21474 42542
rect 21422 42466 21474 42478
rect 22094 42530 22146 42542
rect 22094 42466 22146 42478
rect 25006 42530 25058 42542
rect 25006 42466 25058 42478
rect 28030 42530 28082 42542
rect 36318 42530 36370 42542
rect 32722 42478 32734 42530
rect 32786 42478 32798 42530
rect 28030 42466 28082 42478
rect 36318 42466 36370 42478
rect 39006 42530 39058 42542
rect 39006 42466 39058 42478
rect 40686 42530 40738 42542
rect 40686 42466 40738 42478
rect 42254 42530 42306 42542
rect 42254 42466 42306 42478
rect 42478 42530 42530 42542
rect 43586 42478 43598 42530
rect 43650 42478 43662 42530
rect 42478 42466 42530 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 10222 42194 10274 42206
rect 10222 42130 10274 42142
rect 10894 42194 10946 42206
rect 10894 42130 10946 42142
rect 16494 42194 16546 42206
rect 33294 42194 33346 42206
rect 20626 42142 20638 42194
rect 20690 42142 20702 42194
rect 20962 42142 20974 42194
rect 21026 42142 21038 42194
rect 16494 42130 16546 42142
rect 33294 42130 33346 42142
rect 36654 42194 36706 42206
rect 36654 42130 36706 42142
rect 4734 42082 4786 42094
rect 4734 42018 4786 42030
rect 16382 42082 16434 42094
rect 33406 42082 33458 42094
rect 24210 42030 24222 42082
rect 24274 42030 24286 42082
rect 16382 42018 16434 42030
rect 33406 42018 33458 42030
rect 33742 42082 33794 42094
rect 33742 42018 33794 42030
rect 33854 42082 33906 42094
rect 33854 42018 33906 42030
rect 34302 42082 34354 42094
rect 34302 42018 34354 42030
rect 34414 42082 34466 42094
rect 34414 42018 34466 42030
rect 36766 42082 36818 42094
rect 36766 42018 36818 42030
rect 38110 42082 38162 42094
rect 45726 42082 45778 42094
rect 41234 42030 41246 42082
rect 41298 42030 41310 42082
rect 38110 42018 38162 42030
rect 45726 42018 45778 42030
rect 9662 41970 9714 41982
rect 5058 41918 5070 41970
rect 5122 41918 5134 41970
rect 9662 41906 9714 41918
rect 16718 41970 16770 41982
rect 20302 41970 20354 41982
rect 19618 41918 19630 41970
rect 19682 41918 19694 41970
rect 16718 41906 16770 41918
rect 20302 41906 20354 41918
rect 21534 41970 21586 41982
rect 25118 41970 25170 41982
rect 23202 41918 23214 41970
rect 23266 41918 23278 41970
rect 23650 41918 23662 41970
rect 23714 41918 23726 41970
rect 21534 41906 21586 41918
rect 25118 41906 25170 41918
rect 25454 41970 25506 41982
rect 25454 41906 25506 41918
rect 25790 41970 25842 41982
rect 31502 41970 31554 41982
rect 33070 41970 33122 41982
rect 26674 41918 26686 41970
rect 26738 41918 26750 41970
rect 31938 41918 31950 41970
rect 32002 41918 32014 41970
rect 25790 41906 25842 41918
rect 31502 41906 31554 41918
rect 33070 41906 33122 41918
rect 34078 41970 34130 41982
rect 36094 41970 36146 41982
rect 40014 41970 40066 41982
rect 35410 41918 35422 41970
rect 35474 41918 35486 41970
rect 37426 41918 37438 41970
rect 37490 41918 37502 41970
rect 34078 41906 34130 41918
rect 36094 41906 36146 41918
rect 40014 41906 40066 41918
rect 40910 41970 40962 41982
rect 40910 41906 40962 41918
rect 45838 41970 45890 41982
rect 45838 41906 45890 41918
rect 5518 41858 5570 41870
rect 5518 41794 5570 41806
rect 6190 41858 6242 41870
rect 6190 41794 6242 41806
rect 8990 41858 9042 41870
rect 8990 41794 9042 41806
rect 11342 41858 11394 41870
rect 11342 41794 11394 41806
rect 11790 41858 11842 41870
rect 11790 41794 11842 41806
rect 16046 41858 16098 41870
rect 16046 41794 16098 41806
rect 17502 41858 17554 41870
rect 17502 41794 17554 41806
rect 18958 41858 19010 41870
rect 18958 41794 19010 41806
rect 19182 41858 19234 41870
rect 19182 41794 19234 41806
rect 20078 41858 20130 41870
rect 20078 41794 20130 41806
rect 22318 41858 22370 41870
rect 22318 41794 22370 41806
rect 22766 41858 22818 41870
rect 24670 41858 24722 41870
rect 24098 41806 24110 41858
rect 24162 41806 24174 41858
rect 22766 41794 22818 41806
rect 24670 41794 24722 41806
rect 25342 41858 25394 41870
rect 32398 41858 32450 41870
rect 27458 41806 27470 41858
rect 27522 41806 27534 41858
rect 29586 41806 29598 41858
rect 29650 41806 29662 41858
rect 31042 41806 31054 41858
rect 31106 41806 31118 41858
rect 35634 41806 35646 41858
rect 35698 41806 35710 41858
rect 37202 41806 37214 41858
rect 37266 41806 37278 41858
rect 25342 41794 25394 41806
rect 32398 41794 32450 41806
rect 5070 41746 5122 41758
rect 21310 41746 21362 41758
rect 10994 41694 11006 41746
rect 11058 41743 11070 41746
rect 11330 41743 11342 41746
rect 11058 41697 11342 41743
rect 11058 41694 11070 41697
rect 11330 41694 11342 41697
rect 11394 41743 11406 41746
rect 11778 41743 11790 41746
rect 11394 41697 11790 41743
rect 11394 41694 11406 41697
rect 11778 41694 11790 41697
rect 11842 41694 11854 41746
rect 5070 41682 5122 41694
rect 21310 41682 21362 41694
rect 34414 41746 34466 41758
rect 34414 41682 34466 41694
rect 36654 41746 36706 41758
rect 36654 41682 36706 41694
rect 45726 41746 45778 41758
rect 45726 41682 45778 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 35422 41410 35474 41422
rect 18946 41358 18958 41410
rect 19010 41407 19022 41410
rect 19282 41407 19294 41410
rect 19010 41361 19294 41407
rect 19010 41358 19022 41361
rect 19282 41358 19294 41361
rect 19346 41358 19358 41410
rect 21298 41358 21310 41410
rect 21362 41407 21374 41410
rect 21746 41407 21758 41410
rect 21362 41361 21758 41407
rect 21362 41358 21374 41361
rect 21746 41358 21758 41361
rect 21810 41407 21822 41410
rect 22418 41407 22430 41410
rect 21810 41361 22430 41407
rect 21810 41358 21822 41361
rect 22418 41358 22430 41361
rect 22482 41358 22494 41410
rect 35422 41346 35474 41358
rect 37214 41410 37266 41422
rect 37214 41346 37266 41358
rect 45054 41410 45106 41422
rect 45054 41346 45106 41358
rect 15038 41298 15090 41310
rect 6738 41246 6750 41298
rect 6802 41246 6814 41298
rect 15038 41234 15090 41246
rect 17838 41298 17890 41310
rect 17838 41234 17890 41246
rect 21982 41298 22034 41310
rect 41582 41298 41634 41310
rect 33058 41246 33070 41298
rect 33122 41246 33134 41298
rect 38210 41246 38222 41298
rect 38274 41246 38286 41298
rect 21982 41234 22034 41246
rect 41582 41234 41634 41246
rect 15374 41186 15426 41198
rect 15374 41122 15426 41134
rect 16382 41186 16434 41198
rect 16382 41122 16434 41134
rect 16718 41186 16770 41198
rect 16718 41122 16770 41134
rect 17054 41186 17106 41198
rect 17054 41122 17106 41134
rect 17278 41186 17330 41198
rect 17278 41122 17330 41134
rect 19630 41186 19682 41198
rect 19630 41122 19682 41134
rect 24446 41186 24498 41198
rect 24446 41122 24498 41134
rect 24782 41186 24834 41198
rect 24782 41122 24834 41134
rect 30382 41186 30434 41198
rect 34414 41186 34466 41198
rect 39342 41186 39394 41198
rect 30930 41134 30942 41186
rect 30994 41134 31006 41186
rect 31826 41134 31838 41186
rect 31890 41134 31902 41186
rect 32946 41134 32958 41186
rect 33010 41134 33022 41186
rect 33954 41134 33966 41186
rect 34018 41134 34030 41186
rect 35746 41134 35758 41186
rect 35810 41134 35822 41186
rect 38546 41134 38558 41186
rect 38610 41134 38622 41186
rect 30382 41122 30434 41134
rect 34414 41122 34466 41134
rect 39342 41122 39394 41134
rect 39790 41186 39842 41198
rect 39790 41122 39842 41134
rect 40014 41186 40066 41198
rect 40014 41122 40066 41134
rect 40462 41186 40514 41198
rect 40462 41122 40514 41134
rect 40574 41186 40626 41198
rect 40574 41122 40626 41134
rect 45390 41186 45442 41198
rect 45390 41122 45442 41134
rect 45838 41186 45890 41198
rect 47170 41134 47182 41186
rect 47234 41134 47246 41186
rect 45838 41122 45890 41134
rect 2158 41074 2210 41086
rect 2158 41010 2210 41022
rect 3166 41074 3218 41086
rect 3166 41010 3218 41022
rect 3726 41074 3778 41086
rect 3726 41010 3778 41022
rect 8094 41074 8146 41086
rect 8094 41010 8146 41022
rect 15710 41074 15762 41086
rect 15710 41010 15762 41022
rect 15934 41074 15986 41086
rect 15934 41010 15986 41022
rect 16270 41074 16322 41086
rect 16270 41010 16322 41022
rect 19518 41074 19570 41086
rect 22430 41074 22482 41086
rect 33406 41074 33458 41086
rect 34526 41074 34578 41086
rect 20178 41022 20190 41074
rect 20242 41022 20254 41074
rect 20402 41022 20414 41074
rect 20466 41022 20478 41074
rect 31378 41022 31390 41074
rect 31442 41022 31454 41074
rect 33730 41022 33742 41074
rect 33794 41022 33806 41074
rect 19518 41010 19570 41022
rect 22430 41010 22482 41022
rect 33406 41010 33458 41022
rect 34526 41010 34578 41022
rect 36318 41074 36370 41086
rect 36318 41010 36370 41022
rect 37438 41074 37490 41086
rect 37438 41010 37490 41022
rect 40686 41074 40738 41086
rect 40686 41010 40738 41022
rect 45614 41074 45666 41086
rect 45614 41010 45666 41022
rect 46062 41074 46114 41086
rect 46062 41010 46114 41022
rect 46174 41074 46226 41086
rect 48066 41022 48078 41074
rect 48130 41022 48142 41074
rect 46174 41010 46226 41022
rect 2494 40962 2546 40974
rect 2494 40898 2546 40910
rect 2830 40962 2882 40974
rect 2830 40898 2882 40910
rect 7198 40962 7250 40974
rect 7198 40898 7250 40910
rect 8206 40962 8258 40974
rect 8206 40898 8258 40910
rect 8430 40962 8482 40974
rect 8430 40898 8482 40910
rect 15486 40962 15538 40974
rect 15486 40898 15538 40910
rect 16046 40962 16098 40974
rect 16046 40898 16098 40910
rect 17054 40962 17106 40974
rect 17054 40898 17106 40910
rect 19294 40962 19346 40974
rect 19294 40898 19346 40910
rect 21422 40962 21474 40974
rect 21422 40898 21474 40910
rect 22878 40962 22930 40974
rect 22878 40898 22930 40910
rect 24558 40962 24610 40974
rect 24558 40898 24610 40910
rect 30158 40962 30210 40974
rect 30158 40898 30210 40910
rect 30494 40962 30546 40974
rect 30494 40898 30546 40910
rect 30606 40962 30658 40974
rect 34750 40962 34802 40974
rect 31602 40910 31614 40962
rect 31666 40910 31678 40962
rect 30606 40898 30658 40910
rect 34750 40898 34802 40910
rect 35534 40962 35586 40974
rect 35534 40898 35586 40910
rect 35982 40962 36034 40974
rect 35982 40898 36034 40910
rect 36206 40962 36258 40974
rect 36206 40898 36258 40910
rect 37326 40962 37378 40974
rect 37326 40898 37378 40910
rect 39118 40962 39170 40974
rect 39118 40898 39170 40910
rect 39902 40962 39954 40974
rect 41122 40910 41134 40962
rect 41186 40910 41198 40962
rect 39902 40898 39954 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 5518 40626 5570 40638
rect 4722 40574 4734 40626
rect 4786 40574 4798 40626
rect 5518 40562 5570 40574
rect 9662 40626 9714 40638
rect 9662 40562 9714 40574
rect 16382 40626 16434 40638
rect 16382 40562 16434 40574
rect 16942 40626 16994 40638
rect 16942 40562 16994 40574
rect 21646 40626 21698 40638
rect 21646 40562 21698 40574
rect 23102 40626 23154 40638
rect 23102 40562 23154 40574
rect 23662 40626 23714 40638
rect 23662 40562 23714 40574
rect 24222 40626 24274 40638
rect 32398 40626 32450 40638
rect 31938 40574 31950 40626
rect 32002 40574 32014 40626
rect 24222 40562 24274 40574
rect 32398 40562 32450 40574
rect 34078 40626 34130 40638
rect 34078 40562 34130 40574
rect 34862 40626 34914 40638
rect 34862 40562 34914 40574
rect 38670 40626 38722 40638
rect 41134 40626 41186 40638
rect 39106 40574 39118 40626
rect 39170 40574 39182 40626
rect 38670 40562 38722 40574
rect 41134 40562 41186 40574
rect 41694 40626 41746 40638
rect 41694 40562 41746 40574
rect 42254 40626 42306 40638
rect 42254 40562 42306 40574
rect 42702 40626 42754 40638
rect 42702 40562 42754 40574
rect 11678 40514 11730 40526
rect 16718 40514 16770 40526
rect 21534 40514 21586 40526
rect 2482 40462 2494 40514
rect 2546 40462 2558 40514
rect 7186 40462 7198 40514
rect 7250 40462 7262 40514
rect 8418 40462 8430 40514
rect 8482 40462 8494 40514
rect 12898 40462 12910 40514
rect 12962 40462 12974 40514
rect 18162 40462 18174 40514
rect 18226 40462 18238 40514
rect 11678 40450 11730 40462
rect 16718 40450 16770 40462
rect 21534 40450 21586 40462
rect 22094 40514 22146 40526
rect 22094 40450 22146 40462
rect 22990 40514 23042 40526
rect 22990 40450 23042 40462
rect 23326 40514 23378 40526
rect 23326 40450 23378 40462
rect 23550 40514 23602 40526
rect 23550 40450 23602 40462
rect 33070 40514 33122 40526
rect 33070 40450 33122 40462
rect 33182 40514 33234 40526
rect 33182 40450 33234 40462
rect 34638 40514 34690 40526
rect 41582 40514 41634 40526
rect 40226 40462 40238 40514
rect 40290 40462 40302 40514
rect 34638 40450 34690 40462
rect 41582 40450 41634 40462
rect 44494 40514 44546 40526
rect 44494 40450 44546 40462
rect 45950 40514 46002 40526
rect 45950 40450 46002 40462
rect 16606 40402 16658 40414
rect 20974 40402 21026 40414
rect 1810 40350 1822 40402
rect 1874 40350 1886 40402
rect 5730 40350 5742 40402
rect 5794 40350 5806 40402
rect 8306 40350 8318 40402
rect 8370 40350 8382 40402
rect 11218 40350 11230 40402
rect 11282 40350 11294 40402
rect 12114 40350 12126 40402
rect 12178 40350 12190 40402
rect 17490 40350 17502 40402
rect 17554 40350 17566 40402
rect 16606 40338 16658 40350
rect 20974 40338 21026 40350
rect 22430 40402 22482 40414
rect 22430 40338 22482 40350
rect 22654 40402 22706 40414
rect 30830 40402 30882 40414
rect 25778 40350 25790 40402
rect 25842 40350 25854 40402
rect 26562 40350 26574 40402
rect 26626 40350 26638 40402
rect 30370 40350 30382 40402
rect 30434 40350 30446 40402
rect 22654 40338 22706 40350
rect 30830 40338 30882 40350
rect 31390 40402 31442 40414
rect 31390 40338 31442 40350
rect 31614 40402 31666 40414
rect 38558 40402 38610 40414
rect 34402 40350 34414 40402
rect 34466 40350 34478 40402
rect 35410 40350 35422 40402
rect 35474 40350 35486 40402
rect 35858 40350 35870 40402
rect 35922 40350 35934 40402
rect 37426 40350 37438 40402
rect 37490 40350 37502 40402
rect 31614 40338 31666 40350
rect 38558 40338 38610 40350
rect 38894 40402 38946 40414
rect 39902 40402 39954 40414
rect 39330 40350 39342 40402
rect 39394 40350 39406 40402
rect 38894 40338 38946 40350
rect 39902 40338 39954 40350
rect 41918 40402 41970 40414
rect 43698 40350 43710 40402
rect 43762 40350 43774 40402
rect 45266 40350 45278 40402
rect 45330 40350 45342 40402
rect 41918 40338 41970 40350
rect 10110 40290 10162 40302
rect 22542 40290 22594 40302
rect 15026 40238 15038 40290
rect 15090 40238 15102 40290
rect 20290 40238 20302 40290
rect 20354 40238 20366 40290
rect 10110 40226 10162 40238
rect 22542 40226 22594 40238
rect 24782 40290 24834 40302
rect 34974 40290 35026 40302
rect 28690 40238 28702 40290
rect 28754 40238 28766 40290
rect 35970 40238 35982 40290
rect 36034 40238 36046 40290
rect 37314 40238 37326 40290
rect 37378 40238 37390 40290
rect 43586 40238 43598 40290
rect 43650 40238 43662 40290
rect 45042 40238 45054 40290
rect 45106 40238 45118 40290
rect 24782 40226 24834 40238
rect 34974 40226 35026 40238
rect 6750 40178 6802 40190
rect 6750 40114 6802 40126
rect 21646 40178 21698 40190
rect 21646 40114 21698 40126
rect 23662 40178 23714 40190
rect 33182 40178 33234 40190
rect 23986 40126 23998 40178
rect 24050 40175 24062 40178
rect 24770 40175 24782 40178
rect 24050 40129 24782 40175
rect 24050 40126 24062 40129
rect 24770 40126 24782 40129
rect 24834 40126 24846 40178
rect 36194 40126 36206 40178
rect 36258 40126 36270 40178
rect 37874 40126 37886 40178
rect 37938 40126 37950 40178
rect 42018 40126 42030 40178
rect 42082 40175 42094 40178
rect 42578 40175 42590 40178
rect 42082 40129 42590 40175
rect 42082 40126 42094 40129
rect 42578 40126 42590 40129
rect 42642 40126 42654 40178
rect 23662 40114 23714 40126
rect 33182 40114 33234 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 6862 39842 6914 39854
rect 6862 39778 6914 39790
rect 23102 39842 23154 39854
rect 44158 39842 44210 39854
rect 38882 39790 38894 39842
rect 38946 39839 38958 39842
rect 39330 39839 39342 39842
rect 38946 39793 39342 39839
rect 38946 39790 38958 39793
rect 39330 39790 39342 39793
rect 39394 39790 39406 39842
rect 23102 39778 23154 39790
rect 44158 39778 44210 39790
rect 11902 39730 11954 39742
rect 32062 39730 32114 39742
rect 36318 39730 36370 39742
rect 2482 39678 2494 39730
rect 2546 39678 2558 39730
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 9202 39678 9214 39730
rect 9266 39678 9278 39730
rect 14242 39678 14254 39730
rect 14306 39678 14318 39730
rect 16370 39678 16382 39730
rect 16434 39678 16446 39730
rect 21746 39678 21758 39730
rect 21810 39678 21822 39730
rect 33618 39678 33630 39730
rect 33682 39678 33694 39730
rect 35970 39678 35982 39730
rect 36034 39678 36046 39730
rect 11902 39666 11954 39678
rect 32062 39666 32114 39678
rect 36318 39666 36370 39678
rect 38446 39730 38498 39742
rect 38446 39666 38498 39678
rect 38894 39730 38946 39742
rect 43026 39678 43038 39730
rect 43090 39678 43102 39730
rect 38894 39666 38946 39678
rect 7086 39618 7138 39630
rect 10558 39618 10610 39630
rect 16942 39618 16994 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 7410 39566 7422 39618
rect 7474 39566 7486 39618
rect 13458 39566 13470 39618
rect 13522 39566 13534 39618
rect 7086 39554 7138 39566
rect 10558 39554 10610 39566
rect 16942 39554 16994 39566
rect 17278 39618 17330 39630
rect 17278 39554 17330 39566
rect 22430 39618 22482 39630
rect 22430 39554 22482 39566
rect 23214 39618 23266 39630
rect 23214 39554 23266 39566
rect 23550 39618 23602 39630
rect 23550 39554 23602 39566
rect 23886 39618 23938 39630
rect 32286 39618 32338 39630
rect 24210 39566 24222 39618
rect 24274 39566 24286 39618
rect 25330 39566 25342 39618
rect 25394 39566 25406 39618
rect 25890 39566 25902 39618
rect 25954 39566 25966 39618
rect 23886 39554 23938 39566
rect 32286 39554 32338 39566
rect 32622 39618 32674 39630
rect 35086 39618 35138 39630
rect 40238 39618 40290 39630
rect 33170 39566 33182 39618
rect 33234 39566 33246 39618
rect 33506 39566 33518 39618
rect 33570 39566 33582 39618
rect 35858 39566 35870 39618
rect 35922 39566 35934 39618
rect 32622 39554 32674 39566
rect 35086 39554 35138 39566
rect 40238 39554 40290 39566
rect 40910 39618 40962 39630
rect 40910 39554 40962 39566
rect 41582 39618 41634 39630
rect 41582 39554 41634 39566
rect 41918 39618 41970 39630
rect 43486 39618 43538 39630
rect 42578 39566 42590 39618
rect 42642 39566 42654 39618
rect 41918 39554 41970 39566
rect 43486 39554 43538 39566
rect 45054 39618 45106 39630
rect 45054 39554 45106 39566
rect 45502 39618 45554 39630
rect 45502 39554 45554 39566
rect 5966 39506 6018 39518
rect 23662 39506 23714 39518
rect 34750 39506 34802 39518
rect 7970 39454 7982 39506
rect 8034 39454 8046 39506
rect 9202 39454 9214 39506
rect 9266 39454 9278 39506
rect 20738 39454 20750 39506
rect 20802 39454 20814 39506
rect 26002 39454 26014 39506
rect 26066 39454 26078 39506
rect 33954 39454 33966 39506
rect 34018 39454 34030 39506
rect 5966 39442 6018 39454
rect 23662 39442 23714 39454
rect 34750 39442 34802 39454
rect 34862 39506 34914 39518
rect 34862 39442 34914 39454
rect 39342 39506 39394 39518
rect 39342 39442 39394 39454
rect 39678 39506 39730 39518
rect 41694 39506 41746 39518
rect 41234 39454 41246 39506
rect 41298 39454 41310 39506
rect 39678 39442 39730 39454
rect 41694 39442 41746 39454
rect 43934 39506 43986 39518
rect 43934 39442 43986 39454
rect 5630 39394 5682 39406
rect 11118 39394 11170 39406
rect 6514 39342 6526 39394
rect 6578 39342 6590 39394
rect 5630 39330 5682 39342
rect 11118 39330 11170 39342
rect 17166 39394 17218 39406
rect 17166 39330 17218 39342
rect 17838 39394 17890 39406
rect 17838 39330 17890 39342
rect 20414 39394 20466 39406
rect 20414 39330 20466 39342
rect 21310 39394 21362 39406
rect 21310 39330 21362 39342
rect 22542 39394 22594 39406
rect 22542 39330 22594 39342
rect 22766 39394 22818 39406
rect 22766 39330 22818 39342
rect 23102 39394 23154 39406
rect 23102 39330 23154 39342
rect 32398 39394 32450 39406
rect 32398 39330 32450 39342
rect 37998 39394 38050 39406
rect 37998 39330 38050 39342
rect 44046 39394 44098 39406
rect 44046 39330 44098 39342
rect 44830 39394 44882 39406
rect 44830 39330 44882 39342
rect 44942 39394 44994 39406
rect 44942 39330 44994 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 2606 39058 2658 39070
rect 2606 38994 2658 39006
rect 3950 39058 4002 39070
rect 3950 38994 4002 39006
rect 16494 39058 16546 39070
rect 16494 38994 16546 39006
rect 21310 39058 21362 39070
rect 21310 38994 21362 39006
rect 21870 39058 21922 39070
rect 21870 38994 21922 39006
rect 22318 39058 22370 39070
rect 22318 38994 22370 39006
rect 23214 39058 23266 39070
rect 23214 38994 23266 39006
rect 28814 39058 28866 39070
rect 28814 38994 28866 39006
rect 34638 39058 34690 39070
rect 34638 38994 34690 39006
rect 41470 39058 41522 39070
rect 42254 39058 42306 39070
rect 41794 39006 41806 39058
rect 41858 39006 41870 39058
rect 41470 38994 41522 39006
rect 42254 38994 42306 39006
rect 42926 39058 42978 39070
rect 42926 38994 42978 39006
rect 5406 38946 5458 38958
rect 15486 38946 15538 38958
rect 7186 38894 7198 38946
rect 7250 38894 7262 38946
rect 8082 38894 8094 38946
rect 8146 38894 8158 38946
rect 11666 38894 11678 38946
rect 11730 38894 11742 38946
rect 5406 38882 5458 38894
rect 15486 38882 15538 38894
rect 15822 38946 15874 38958
rect 25230 38946 25282 38958
rect 23986 38894 23998 38946
rect 24050 38894 24062 38946
rect 15822 38882 15874 38894
rect 25230 38882 25282 38894
rect 25566 38946 25618 38958
rect 25566 38882 25618 38894
rect 25790 38946 25842 38958
rect 25790 38882 25842 38894
rect 26238 38946 26290 38958
rect 26238 38882 26290 38894
rect 26798 38946 26850 38958
rect 30942 38946 30994 38958
rect 29586 38894 29598 38946
rect 29650 38894 29662 38946
rect 29810 38894 29822 38946
rect 29874 38894 29886 38946
rect 26798 38882 26850 38894
rect 30942 38882 30994 38894
rect 42702 38946 42754 38958
rect 42702 38882 42754 38894
rect 43710 38946 43762 38958
rect 43710 38882 43762 38894
rect 48190 38946 48242 38958
rect 48190 38882 48242 38894
rect 1710 38834 1762 38846
rect 1710 38770 1762 38782
rect 2942 38834 2994 38846
rect 2942 38770 2994 38782
rect 3390 38834 3442 38846
rect 26126 38834 26178 38846
rect 7298 38782 7310 38834
rect 7362 38782 7374 38834
rect 8306 38782 8318 38834
rect 8370 38782 8382 38834
rect 12338 38782 12350 38834
rect 12402 38782 12414 38834
rect 16258 38782 16270 38834
rect 16322 38782 16334 38834
rect 23538 38782 23550 38834
rect 23602 38782 23614 38834
rect 24658 38782 24670 38834
rect 24722 38782 24734 38834
rect 3390 38770 3442 38782
rect 26126 38770 26178 38782
rect 26462 38834 26514 38846
rect 35198 38834 35250 38846
rect 29362 38782 29374 38834
rect 29426 38782 29438 38834
rect 33506 38782 33518 38834
rect 33570 38782 33582 38834
rect 43362 38782 43374 38834
rect 43426 38782 43438 38834
rect 26462 38770 26514 38782
rect 35198 38770 35250 38782
rect 25342 38722 25394 38734
rect 2146 38670 2158 38722
rect 2210 38670 2222 38722
rect 8418 38670 8430 38722
rect 8482 38670 8494 38722
rect 9538 38670 9550 38722
rect 9602 38670 9614 38722
rect 24210 38670 24222 38722
rect 24274 38670 24286 38722
rect 25342 38658 25394 38670
rect 30494 38722 30546 38734
rect 41022 38722 41074 38734
rect 33618 38670 33630 38722
rect 33682 38670 33694 38722
rect 43026 38670 43038 38722
rect 43090 38670 43102 38722
rect 30494 38658 30546 38670
rect 41022 38658 41074 38670
rect 43374 38610 43426 38622
rect 5058 38558 5070 38610
rect 5122 38607 5134 38610
rect 5506 38607 5518 38610
rect 5122 38561 5518 38607
rect 5122 38558 5134 38561
rect 5506 38558 5518 38561
rect 5570 38558 5582 38610
rect 33394 38558 33406 38610
rect 33458 38558 33470 38610
rect 43374 38546 43426 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 8206 38274 8258 38286
rect 8206 38210 8258 38222
rect 20750 38274 20802 38286
rect 20750 38210 20802 38222
rect 24894 38274 24946 38286
rect 24894 38210 24946 38222
rect 34190 38274 34242 38286
rect 34190 38210 34242 38222
rect 1822 38162 1874 38174
rect 1822 38098 1874 38110
rect 8430 38162 8482 38174
rect 34414 38162 34466 38174
rect 9650 38110 9662 38162
rect 9714 38110 9726 38162
rect 11778 38110 11790 38162
rect 11842 38110 11854 38162
rect 15362 38110 15374 38162
rect 15426 38110 15438 38162
rect 17490 38110 17502 38162
rect 17554 38110 17566 38162
rect 28466 38110 28478 38162
rect 28530 38110 28542 38162
rect 8430 38098 8482 38110
rect 34414 38098 34466 38110
rect 34974 38162 35026 38174
rect 38434 38110 38446 38162
rect 38498 38110 38510 38162
rect 34974 38098 35026 38110
rect 3838 38050 3890 38062
rect 25006 38050 25058 38062
rect 29598 38050 29650 38062
rect 8866 37998 8878 38050
rect 8930 37998 8942 38050
rect 14690 37998 14702 38050
rect 14754 37998 14766 38050
rect 18498 37998 18510 38050
rect 18562 37998 18574 38050
rect 19618 37998 19630 38050
rect 19682 37998 19694 38050
rect 27010 37998 27022 38050
rect 27074 37998 27086 38050
rect 27458 37998 27470 38050
rect 27522 37998 27534 38050
rect 3838 37986 3890 37998
rect 25006 37986 25058 37998
rect 29598 37986 29650 37998
rect 29822 38050 29874 38062
rect 29822 37986 29874 37998
rect 29934 38050 29986 38062
rect 29934 37986 29986 37998
rect 38782 38050 38834 38062
rect 39890 37998 39902 38050
rect 39954 37998 39966 38050
rect 38782 37986 38834 37998
rect 29486 37938 29538 37950
rect 18162 37886 18174 37938
rect 18226 37886 18238 37938
rect 29486 37874 29538 37886
rect 30718 37938 30770 37950
rect 30718 37874 30770 37886
rect 30830 37938 30882 37950
rect 30830 37874 30882 37886
rect 3726 37826 3778 37838
rect 24894 37826 24946 37838
rect 7858 37774 7870 37826
rect 7922 37774 7934 37826
rect 3726 37762 3778 37774
rect 24894 37762 24946 37774
rect 25566 37826 25618 37838
rect 25566 37762 25618 37774
rect 30494 37826 30546 37838
rect 38558 37826 38610 37838
rect 33842 37774 33854 37826
rect 33906 37774 33918 37826
rect 30494 37762 30546 37774
rect 38558 37762 38610 37774
rect 39230 37826 39282 37838
rect 39230 37762 39282 37774
rect 39678 37826 39730 37838
rect 39678 37762 39730 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 8990 37490 9042 37502
rect 8990 37426 9042 37438
rect 18062 37490 18114 37502
rect 18062 37426 18114 37438
rect 18286 37490 18338 37502
rect 18286 37426 18338 37438
rect 18510 37490 18562 37502
rect 18510 37426 18562 37438
rect 26574 37490 26626 37502
rect 26574 37426 26626 37438
rect 27246 37490 27298 37502
rect 27246 37426 27298 37438
rect 41918 37490 41970 37502
rect 41918 37426 41970 37438
rect 22654 37378 22706 37390
rect 5058 37326 5070 37378
rect 5122 37326 5134 37378
rect 12338 37326 12350 37378
rect 12402 37326 12414 37378
rect 19506 37326 19518 37378
rect 19570 37326 19582 37378
rect 22654 37314 22706 37326
rect 26686 37378 26738 37390
rect 39566 37378 39618 37390
rect 34962 37326 34974 37378
rect 35026 37326 35038 37378
rect 38098 37326 38110 37378
rect 38162 37326 38174 37378
rect 26686 37314 26738 37326
rect 39566 37314 39618 37326
rect 44270 37378 44322 37390
rect 45938 37326 45950 37378
rect 46002 37326 46014 37378
rect 44270 37314 44322 37326
rect 9550 37266 9602 37278
rect 4386 37214 4398 37266
rect 4450 37214 4462 37266
rect 9550 37202 9602 37214
rect 9774 37266 9826 37278
rect 15710 37266 15762 37278
rect 11554 37214 11566 37266
rect 11618 37214 11630 37266
rect 9774 37202 9826 37214
rect 15710 37202 15762 37214
rect 16270 37266 16322 37278
rect 16270 37202 16322 37214
rect 18622 37266 18674 37278
rect 28030 37266 28082 37278
rect 31502 37266 31554 37278
rect 40910 37266 40962 37278
rect 19842 37214 19854 37266
rect 19906 37214 19918 37266
rect 20850 37214 20862 37266
rect 20914 37214 20926 37266
rect 21970 37214 21982 37266
rect 22034 37214 22046 37266
rect 28130 37214 28142 37266
rect 28194 37214 28206 37266
rect 29586 37214 29598 37266
rect 29650 37214 29662 37266
rect 31266 37214 31278 37266
rect 31330 37214 31342 37266
rect 34738 37214 34750 37266
rect 34802 37214 34814 37266
rect 38434 37214 38446 37266
rect 38498 37214 38510 37266
rect 18622 37202 18674 37214
rect 28030 37202 28082 37214
rect 31502 37202 31554 37214
rect 40910 37202 40962 37214
rect 41134 37266 41186 37278
rect 41134 37202 41186 37214
rect 41806 37266 41858 37278
rect 41806 37202 41858 37214
rect 42142 37266 42194 37278
rect 43362 37214 43374 37266
rect 43426 37214 43438 37266
rect 46834 37214 46846 37266
rect 46898 37214 46910 37266
rect 42142 37202 42194 37214
rect 1822 37154 1874 37166
rect 7646 37154 7698 37166
rect 15374 37154 15426 37166
rect 26126 37154 26178 37166
rect 30158 37154 30210 37166
rect 7186 37102 7198 37154
rect 7250 37102 7262 37154
rect 14466 37102 14478 37154
rect 14530 37102 14542 37154
rect 19954 37102 19966 37154
rect 20018 37102 20030 37154
rect 20402 37102 20414 37154
rect 20466 37102 20478 37154
rect 28578 37102 28590 37154
rect 28642 37102 28654 37154
rect 29250 37102 29262 37154
rect 29314 37102 29326 37154
rect 1822 37090 1874 37102
rect 7646 37090 7698 37102
rect 15374 37090 15426 37102
rect 26126 37090 26178 37102
rect 30158 37090 30210 37102
rect 31838 37154 31890 37166
rect 40226 37102 40238 37154
rect 40290 37102 40302 37154
rect 43474 37102 43486 37154
rect 43538 37102 43550 37154
rect 45378 37102 45390 37154
rect 45442 37102 45454 37154
rect 47842 37102 47854 37154
rect 47906 37102 47918 37154
rect 31838 37090 31890 37102
rect 26574 37042 26626 37054
rect 32062 37042 32114 37054
rect 10098 36990 10110 37042
rect 10162 36990 10174 37042
rect 28466 36990 28478 37042
rect 28530 36990 28542 37042
rect 30818 36990 30830 37042
rect 30882 36990 30894 37042
rect 32386 36990 32398 37042
rect 32450 36990 32462 37042
rect 41458 36990 41470 37042
rect 41522 36990 41534 37042
rect 26574 36978 26626 36990
rect 32062 36978 32114 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 19742 36706 19794 36718
rect 45950 36706 46002 36718
rect 22194 36654 22206 36706
rect 22258 36703 22270 36706
rect 23090 36703 23102 36706
rect 22258 36657 23102 36703
rect 22258 36654 22270 36657
rect 23090 36654 23102 36657
rect 23154 36654 23166 36706
rect 28354 36654 28366 36706
rect 28418 36654 28430 36706
rect 19742 36642 19794 36654
rect 45950 36642 46002 36654
rect 2270 36594 2322 36606
rect 2270 36530 2322 36542
rect 4398 36594 4450 36606
rect 4398 36530 4450 36542
rect 8766 36594 8818 36606
rect 17950 36594 18002 36606
rect 10434 36542 10446 36594
rect 10498 36542 10510 36594
rect 12562 36542 12574 36594
rect 12626 36542 12638 36594
rect 14242 36542 14254 36594
rect 14306 36542 14318 36594
rect 8766 36530 8818 36542
rect 17950 36530 18002 36542
rect 18398 36594 18450 36606
rect 18398 36530 18450 36542
rect 19070 36594 19122 36606
rect 19070 36530 19122 36542
rect 20302 36594 20354 36606
rect 20302 36530 20354 36542
rect 22318 36594 22370 36606
rect 22318 36530 22370 36542
rect 22654 36594 22706 36606
rect 22654 36530 22706 36542
rect 23102 36594 23154 36606
rect 46398 36594 46450 36606
rect 27794 36542 27806 36594
rect 27858 36542 27870 36594
rect 29922 36542 29934 36594
rect 29986 36542 29998 36594
rect 30930 36542 30942 36594
rect 30994 36542 31006 36594
rect 23102 36530 23154 36542
rect 46398 36530 46450 36542
rect 4510 36482 4562 36494
rect 4510 36418 4562 36430
rect 5854 36482 5906 36494
rect 5854 36418 5906 36430
rect 7758 36482 7810 36494
rect 7758 36418 7810 36430
rect 7982 36482 8034 36494
rect 7982 36418 8034 36430
rect 8318 36482 8370 36494
rect 39454 36482 39506 36494
rect 9650 36430 9662 36482
rect 9714 36430 9726 36482
rect 14578 36430 14590 36482
rect 14642 36430 14654 36482
rect 23762 36430 23774 36482
rect 23826 36430 23838 36482
rect 25666 36430 25678 36482
rect 25730 36430 25742 36482
rect 26226 36430 26238 36482
rect 26290 36430 26302 36482
rect 27122 36430 27134 36482
rect 27186 36430 27198 36482
rect 28018 36430 28030 36482
rect 28082 36430 28094 36482
rect 30034 36430 30046 36482
rect 30098 36430 30110 36482
rect 32610 36430 32622 36482
rect 32674 36430 32686 36482
rect 8318 36418 8370 36430
rect 39454 36418 39506 36430
rect 39790 36482 39842 36494
rect 39790 36418 39842 36430
rect 41246 36482 41298 36494
rect 41246 36418 41298 36430
rect 41694 36482 41746 36494
rect 41694 36418 41746 36430
rect 45614 36482 45666 36494
rect 45614 36418 45666 36430
rect 46174 36482 46226 36494
rect 46174 36418 46226 36430
rect 46846 36482 46898 36494
rect 46846 36418 46898 36430
rect 3838 36370 3890 36382
rect 3838 36306 3890 36318
rect 5070 36370 5122 36382
rect 5070 36306 5122 36318
rect 17166 36370 17218 36382
rect 17166 36306 17218 36318
rect 19742 36370 19794 36382
rect 19742 36306 19794 36318
rect 19854 36370 19906 36382
rect 19854 36306 19906 36318
rect 23438 36370 23490 36382
rect 23438 36306 23490 36318
rect 30494 36370 30546 36382
rect 33070 36370 33122 36382
rect 31154 36318 31166 36370
rect 31218 36318 31230 36370
rect 30494 36306 30546 36318
rect 33070 36306 33122 36318
rect 39118 36370 39170 36382
rect 39118 36306 39170 36318
rect 39902 36370 39954 36382
rect 39902 36306 39954 36318
rect 40014 36370 40066 36382
rect 40014 36306 40066 36318
rect 40910 36370 40962 36382
rect 40910 36306 40962 36318
rect 1710 36258 1762 36270
rect 1710 36194 1762 36206
rect 4846 36258 4898 36270
rect 4846 36194 4898 36206
rect 5182 36258 5234 36270
rect 5182 36194 5234 36206
rect 5630 36258 5682 36270
rect 5630 36194 5682 36206
rect 5742 36258 5794 36270
rect 5742 36194 5794 36206
rect 6078 36258 6130 36270
rect 6078 36194 6130 36206
rect 7422 36258 7474 36270
rect 7422 36194 7474 36206
rect 8206 36258 8258 36270
rect 8206 36194 8258 36206
rect 17390 36258 17442 36270
rect 17390 36194 17442 36206
rect 24222 36258 24274 36270
rect 24222 36194 24274 36206
rect 25006 36258 25058 36270
rect 25006 36194 25058 36206
rect 38446 36258 38498 36270
rect 38446 36194 38498 36206
rect 38782 36258 38834 36270
rect 38782 36194 38834 36206
rect 40574 36258 40626 36270
rect 40574 36194 40626 36206
rect 46622 36258 46674 36270
rect 46622 36194 46674 36206
rect 46734 36258 46786 36270
rect 46734 36194 46786 36206
rect 48190 36258 48242 36270
rect 48190 36194 48242 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 17726 35922 17778 35934
rect 17726 35858 17778 35870
rect 20974 35922 21026 35934
rect 20974 35858 21026 35870
rect 26350 35922 26402 35934
rect 26350 35858 26402 35870
rect 40014 35922 40066 35934
rect 40014 35858 40066 35870
rect 40350 35922 40402 35934
rect 40350 35858 40402 35870
rect 11566 35810 11618 35822
rect 5282 35758 5294 35810
rect 5346 35758 5358 35810
rect 6850 35758 6862 35810
rect 6914 35758 6926 35810
rect 11566 35746 11618 35758
rect 17950 35810 18002 35822
rect 29374 35810 29426 35822
rect 19730 35758 19742 35810
rect 19794 35758 19806 35810
rect 17950 35746 18002 35758
rect 29374 35746 29426 35758
rect 29486 35810 29538 35822
rect 29486 35746 29538 35758
rect 29934 35810 29986 35822
rect 29934 35746 29986 35758
rect 39678 35810 39730 35822
rect 39678 35746 39730 35758
rect 39790 35810 39842 35822
rect 39790 35746 39842 35758
rect 41134 35810 41186 35822
rect 43038 35810 43090 35822
rect 42354 35758 42366 35810
rect 42418 35758 42430 35810
rect 41134 35746 41186 35758
rect 43038 35746 43090 35758
rect 45390 35810 45442 35822
rect 45390 35746 45442 35758
rect 46846 35810 46898 35822
rect 46846 35746 46898 35758
rect 27806 35698 27858 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 8082 35646 8094 35698
rect 8146 35646 8158 35698
rect 17490 35646 17502 35698
rect 17554 35646 17566 35698
rect 18162 35646 18174 35698
rect 18226 35646 18238 35698
rect 18834 35646 18846 35698
rect 18898 35646 18910 35698
rect 19170 35646 19182 35698
rect 19234 35646 19246 35698
rect 21746 35646 21758 35698
rect 21810 35646 21822 35698
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 27806 35634 27858 35646
rect 31054 35698 31106 35710
rect 31054 35634 31106 35646
rect 31838 35698 31890 35710
rect 41358 35698 41410 35710
rect 34402 35646 34414 35698
rect 34466 35646 34478 35698
rect 36418 35646 36430 35698
rect 36482 35646 36494 35698
rect 38098 35646 38110 35698
rect 38162 35646 38174 35698
rect 38994 35646 39006 35698
rect 39058 35646 39070 35698
rect 42466 35646 42478 35698
rect 42530 35646 42542 35698
rect 43362 35646 43374 35698
rect 43426 35646 43438 35698
rect 46162 35646 46174 35698
rect 46226 35646 46238 35698
rect 31838 35634 31890 35646
rect 41358 35634 41410 35646
rect 4958 35586 5010 35598
rect 2482 35534 2494 35586
rect 2546 35534 2558 35586
rect 4610 35534 4622 35586
rect 4674 35534 4686 35586
rect 4958 35522 5010 35534
rect 6974 35586 7026 35598
rect 17838 35586 17890 35598
rect 25902 35586 25954 35598
rect 8418 35534 8430 35586
rect 8482 35534 8494 35586
rect 11218 35534 11230 35586
rect 11282 35534 11294 35586
rect 19058 35534 19070 35586
rect 19122 35534 19134 35586
rect 21298 35534 21310 35586
rect 21362 35534 21374 35586
rect 23426 35534 23438 35586
rect 23490 35534 23502 35586
rect 6974 35522 7026 35534
rect 17838 35522 17890 35534
rect 25902 35522 25954 35534
rect 26798 35586 26850 35598
rect 26798 35522 26850 35534
rect 27358 35586 27410 35598
rect 27358 35522 27410 35534
rect 28254 35586 28306 35598
rect 28254 35522 28306 35534
rect 28702 35586 28754 35598
rect 28702 35522 28754 35534
rect 31390 35586 31442 35598
rect 34850 35534 34862 35586
rect 34914 35534 34926 35586
rect 38546 35534 38558 35586
rect 38610 35534 38622 35586
rect 42354 35534 42366 35586
rect 42418 35534 42430 35586
rect 43250 35534 43262 35586
rect 43314 35534 43326 35586
rect 46050 35534 46062 35586
rect 46114 35534 46126 35586
rect 31390 35522 31442 35534
rect 29486 35474 29538 35486
rect 39006 35474 39058 35486
rect 8642 35422 8654 35474
rect 8706 35422 8718 35474
rect 25778 35422 25790 35474
rect 25842 35471 25854 35474
rect 26338 35471 26350 35474
rect 25842 35425 26350 35471
rect 25842 35422 25854 35425
rect 26338 35422 26350 35425
rect 26402 35422 26414 35474
rect 30482 35422 30494 35474
rect 30546 35422 30558 35474
rect 37202 35422 37214 35474
rect 37266 35422 37278 35474
rect 29486 35410 29538 35422
rect 39006 35410 39058 35422
rect 39342 35474 39394 35486
rect 39342 35410 39394 35422
rect 41694 35474 41746 35486
rect 41694 35410 41746 35422
rect 45502 35474 45554 35486
rect 45502 35410 45554 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 4610 35086 4622 35138
rect 4674 35086 4686 35138
rect 18834 35086 18846 35138
rect 18898 35086 18910 35138
rect 20626 35086 20638 35138
rect 20690 35086 20702 35138
rect 32162 35086 32174 35138
rect 32226 35086 32238 35138
rect 39666 35086 39678 35138
rect 39730 35086 39742 35138
rect 4062 35026 4114 35038
rect 4062 34962 4114 34974
rect 5070 35026 5122 35038
rect 5070 34962 5122 34974
rect 8878 35026 8930 35038
rect 26350 35026 26402 35038
rect 20178 34974 20190 35026
rect 20242 34974 20254 35026
rect 28466 34974 28478 35026
rect 28530 34974 28542 35026
rect 32274 34974 32286 35026
rect 32338 34974 32350 35026
rect 33394 34974 33406 35026
rect 33458 34974 33470 35026
rect 45378 34974 45390 35026
rect 45442 34974 45454 35026
rect 8878 34962 8930 34974
rect 26350 34962 26402 34974
rect 4286 34914 4338 34926
rect 2258 34862 2270 34914
rect 2322 34862 2334 34914
rect 4286 34850 4338 34862
rect 5966 34914 6018 34926
rect 5966 34850 6018 34862
rect 6190 34914 6242 34926
rect 11566 34914 11618 34926
rect 8418 34862 8430 34914
rect 8482 34862 8494 34914
rect 6190 34850 6242 34862
rect 11566 34850 11618 34862
rect 16046 34914 16098 34926
rect 20414 34914 20466 34926
rect 17826 34862 17838 34914
rect 17890 34862 17902 34914
rect 18498 34862 18510 34914
rect 18562 34862 18574 34914
rect 18946 34862 18958 34914
rect 19010 34862 19022 34914
rect 16046 34850 16098 34862
rect 20414 34850 20466 34862
rect 21646 34914 21698 34926
rect 21646 34850 21698 34862
rect 21982 34914 22034 34926
rect 31166 34914 31218 34926
rect 38446 34914 38498 34926
rect 41246 34914 41298 34926
rect 22306 34862 22318 34914
rect 22370 34862 22382 34914
rect 22754 34862 22766 34914
rect 22818 34862 22830 34914
rect 23426 34862 23438 34914
rect 23490 34862 23502 34914
rect 24210 34862 24222 34914
rect 24274 34862 24286 34914
rect 24882 34862 24894 34914
rect 24946 34862 24958 34914
rect 25778 34862 25790 34914
rect 25842 34862 25854 34914
rect 27010 34862 27022 34914
rect 27074 34862 27086 34914
rect 31826 34862 31838 34914
rect 31890 34862 31902 34914
rect 32050 34862 32062 34914
rect 32114 34862 32126 34914
rect 33282 34862 33294 34914
rect 33346 34862 33358 34914
rect 34962 34862 34974 34914
rect 35026 34862 35038 34914
rect 37762 34862 37774 34914
rect 37826 34862 37838 34914
rect 39218 34862 39230 34914
rect 39282 34862 39294 34914
rect 21982 34850 22034 34862
rect 31166 34850 31218 34862
rect 38446 34850 38498 34862
rect 41246 34850 41298 34862
rect 41470 34914 41522 34926
rect 41470 34850 41522 34862
rect 42030 34914 42082 34926
rect 42030 34850 42082 34862
rect 42478 34914 42530 34926
rect 42914 34862 42926 34914
rect 42978 34862 42990 34914
rect 45154 34862 45166 34914
rect 45218 34862 45230 34914
rect 42478 34850 42530 34862
rect 2494 34802 2546 34814
rect 2494 34738 2546 34750
rect 3838 34802 3890 34814
rect 7534 34802 7586 34814
rect 6626 34750 6638 34802
rect 6690 34750 6702 34802
rect 6850 34750 6862 34802
rect 6914 34750 6926 34802
rect 3838 34738 3890 34750
rect 7534 34738 7586 34750
rect 7758 34802 7810 34814
rect 17950 34802 18002 34814
rect 16706 34750 16718 34802
rect 16770 34750 16782 34802
rect 7758 34738 7810 34750
rect 17950 34738 18002 34750
rect 21310 34802 21362 34814
rect 21310 34738 21362 34750
rect 21422 34802 21474 34814
rect 29822 34802 29874 34814
rect 35646 34802 35698 34814
rect 27906 34750 27918 34802
rect 27970 34750 27982 34802
rect 30818 34750 30830 34802
rect 30882 34750 30894 34802
rect 21422 34738 21474 34750
rect 29822 34738 29874 34750
rect 35646 34738 35698 34750
rect 36094 34802 36146 34814
rect 36094 34738 36146 34750
rect 36206 34802 36258 34814
rect 36206 34738 36258 34750
rect 40910 34802 40962 34814
rect 40910 34738 40962 34750
rect 41022 34802 41074 34814
rect 41022 34738 41074 34750
rect 43374 34802 43426 34814
rect 43374 34738 43426 34750
rect 45838 34802 45890 34814
rect 45838 34738 45890 34750
rect 5742 34690 5794 34702
rect 5742 34626 5794 34638
rect 7982 34690 8034 34702
rect 7982 34626 8034 34638
rect 8094 34690 8146 34702
rect 8094 34626 8146 34638
rect 9326 34690 9378 34702
rect 9326 34626 9378 34638
rect 9774 34690 9826 34702
rect 15486 34690 15538 34702
rect 11890 34638 11902 34690
rect 11954 34638 11966 34690
rect 9774 34626 9826 34638
rect 15486 34626 15538 34638
rect 16382 34690 16434 34702
rect 16382 34626 16434 34638
rect 17390 34690 17442 34702
rect 17390 34626 17442 34638
rect 29262 34690 29314 34702
rect 35310 34690 35362 34702
rect 34738 34638 34750 34690
rect 34802 34638 34814 34690
rect 29262 34626 29314 34638
rect 35310 34626 35362 34638
rect 35534 34690 35586 34702
rect 35534 34626 35586 34638
rect 35870 34690 35922 34702
rect 35870 34626 35922 34638
rect 37102 34690 37154 34702
rect 37102 34626 37154 34638
rect 40350 34690 40402 34702
rect 40350 34626 40402 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 2718 34354 2770 34366
rect 2718 34290 2770 34302
rect 4286 34354 4338 34366
rect 4286 34290 4338 34302
rect 4622 34354 4674 34366
rect 4622 34290 4674 34302
rect 9102 34354 9154 34366
rect 21422 34354 21474 34366
rect 17714 34302 17726 34354
rect 17778 34302 17790 34354
rect 9102 34290 9154 34302
rect 21422 34290 21474 34302
rect 24558 34354 24610 34366
rect 24558 34290 24610 34302
rect 27022 34354 27074 34366
rect 27022 34290 27074 34302
rect 29038 34354 29090 34366
rect 29038 34290 29090 34302
rect 29486 34354 29538 34366
rect 29486 34290 29538 34302
rect 40238 34354 40290 34366
rect 40238 34290 40290 34302
rect 43598 34354 43650 34366
rect 43598 34290 43650 34302
rect 44830 34354 44882 34366
rect 44830 34290 44882 34302
rect 45502 34354 45554 34366
rect 45502 34290 45554 34302
rect 47742 34354 47794 34366
rect 47742 34290 47794 34302
rect 8542 34242 8594 34254
rect 16494 34242 16546 34254
rect 23662 34242 23714 34254
rect 5170 34190 5182 34242
rect 5234 34190 5246 34242
rect 5730 34190 5742 34242
rect 5794 34190 5806 34242
rect 13906 34190 13918 34242
rect 13970 34190 13982 34242
rect 15922 34190 15934 34242
rect 15986 34190 15998 34242
rect 22082 34190 22094 34242
rect 22146 34190 22158 34242
rect 8542 34178 8594 34190
rect 16494 34178 16546 34190
rect 23662 34178 23714 34190
rect 34190 34242 34242 34254
rect 34190 34178 34242 34190
rect 34638 34242 34690 34254
rect 34638 34178 34690 34190
rect 35198 34242 35250 34254
rect 45054 34242 45106 34254
rect 35858 34190 35870 34242
rect 35922 34190 35934 34242
rect 38098 34190 38110 34242
rect 38162 34190 38174 34242
rect 35198 34178 35250 34190
rect 45054 34178 45106 34190
rect 45726 34242 45778 34254
rect 45726 34178 45778 34190
rect 46622 34242 46674 34254
rect 46622 34178 46674 34190
rect 47182 34242 47234 34254
rect 47182 34178 47234 34190
rect 48190 34242 48242 34254
rect 48190 34178 48242 34190
rect 1710 34130 1762 34142
rect 1710 34066 1762 34078
rect 2270 34130 2322 34142
rect 12462 34130 12514 34142
rect 16270 34130 16322 34142
rect 17390 34130 17442 34142
rect 42926 34130 42978 34142
rect 5058 34078 5070 34130
rect 5122 34078 5134 34130
rect 6514 34078 6526 34130
rect 6578 34078 6590 34130
rect 6850 34078 6862 34130
rect 6914 34078 6926 34130
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 14690 34078 14702 34130
rect 14754 34078 14766 34130
rect 16818 34078 16830 34130
rect 16882 34078 16894 34130
rect 18834 34078 18846 34130
rect 18898 34078 18910 34130
rect 25442 34078 25454 34130
rect 25506 34078 25518 34130
rect 27906 34078 27918 34130
rect 27970 34078 27982 34130
rect 33282 34078 33294 34130
rect 33346 34078 33358 34130
rect 36866 34078 36878 34130
rect 36930 34078 36942 34130
rect 37762 34078 37774 34130
rect 37826 34078 37838 34130
rect 41010 34078 41022 34130
rect 41074 34078 41086 34130
rect 2270 34066 2322 34078
rect 12462 34066 12514 34078
rect 16270 34066 16322 34078
rect 17390 34066 17442 34078
rect 42926 34066 42978 34078
rect 43262 34130 43314 34142
rect 43262 34066 43314 34078
rect 43486 34130 43538 34142
rect 44718 34130 44770 34142
rect 44258 34078 44270 34130
rect 44322 34127 44334 34130
rect 44482 34127 44494 34130
rect 44322 34081 44494 34127
rect 44322 34078 44334 34081
rect 44482 34078 44494 34081
rect 44546 34078 44558 34130
rect 43486 34066 43538 34078
rect 44718 34066 44770 34078
rect 45278 34130 45330 34142
rect 45278 34066 45330 34078
rect 3390 34018 3442 34030
rect 2706 33966 2718 34018
rect 2770 33966 2782 34018
rect 3390 33954 3442 33966
rect 6190 34018 6242 34030
rect 16382 34018 16434 34030
rect 7970 33966 7982 34018
rect 8034 33966 8046 34018
rect 13570 33966 13582 34018
rect 13634 33966 13646 34018
rect 6190 33954 6242 33966
rect 16382 33954 16434 33966
rect 19294 34018 19346 34030
rect 26574 34018 26626 34030
rect 28590 34018 28642 34030
rect 34750 34018 34802 34030
rect 22306 33966 22318 34018
rect 22370 33966 22382 34018
rect 25554 33966 25566 34018
rect 25618 33966 25630 34018
rect 28242 33966 28254 34018
rect 28306 33966 28318 34018
rect 33394 33966 33406 34018
rect 33458 33966 33470 34018
rect 19294 33954 19346 33966
rect 26574 33954 26626 33966
rect 28590 33954 28642 33966
rect 34750 33954 34802 33966
rect 39678 34018 39730 34030
rect 45390 34018 45442 34030
rect 41682 33966 41694 34018
rect 41746 33966 41758 34018
rect 39678 33954 39730 33966
rect 45390 33954 45442 33966
rect 2942 33906 2994 33918
rect 2942 33842 2994 33854
rect 8430 33906 8482 33918
rect 34862 33906 34914 33918
rect 8866 33854 8878 33906
rect 8930 33903 8942 33906
rect 9090 33903 9102 33906
rect 8930 33857 9102 33903
rect 8930 33854 8942 33857
rect 9090 33854 9102 33857
rect 9154 33854 9166 33906
rect 25890 33854 25902 33906
rect 25954 33854 25966 33906
rect 8430 33842 8482 33854
rect 34862 33842 34914 33854
rect 35310 33906 35362 33918
rect 35310 33842 35362 33854
rect 42702 33906 42754 33918
rect 42702 33842 42754 33854
rect 46510 33906 46562 33918
rect 46510 33842 46562 33854
rect 46846 33906 46898 33918
rect 46846 33842 46898 33854
rect 47294 33906 47346 33918
rect 47294 33842 47346 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 2158 33570 2210 33582
rect 2158 33506 2210 33518
rect 12686 33570 12738 33582
rect 12686 33506 12738 33518
rect 13806 33570 13858 33582
rect 13806 33506 13858 33518
rect 14142 33570 14194 33582
rect 14142 33506 14194 33518
rect 19630 33570 19682 33582
rect 19630 33506 19682 33518
rect 19966 33570 20018 33582
rect 19966 33506 20018 33518
rect 2942 33458 2994 33470
rect 2482 33406 2494 33458
rect 2546 33406 2558 33458
rect 2942 33394 2994 33406
rect 3390 33458 3442 33470
rect 3390 33394 3442 33406
rect 3838 33458 3890 33470
rect 18174 33458 18226 33470
rect 37998 33458 38050 33470
rect 14690 33406 14702 33458
rect 14754 33406 14766 33458
rect 25330 33406 25342 33458
rect 25394 33406 25406 33458
rect 27458 33406 27470 33458
rect 27522 33406 27534 33458
rect 37090 33406 37102 33458
rect 37154 33406 37166 33458
rect 3838 33394 3890 33406
rect 18174 33394 18226 33406
rect 37998 33394 38050 33406
rect 44270 33458 44322 33470
rect 44270 33394 44322 33406
rect 1934 33346 1986 33358
rect 6750 33346 6802 33358
rect 9550 33346 9602 33358
rect 5954 33294 5966 33346
rect 6018 33294 6030 33346
rect 7074 33294 7086 33346
rect 7138 33294 7150 33346
rect 1934 33282 1986 33294
rect 6750 33282 6802 33294
rect 9550 33282 9602 33294
rect 12238 33346 12290 33358
rect 12238 33282 12290 33294
rect 12574 33346 12626 33358
rect 30382 33346 30434 33358
rect 38446 33346 38498 33358
rect 42702 33346 42754 33358
rect 14914 33294 14926 33346
rect 14978 33294 14990 33346
rect 21298 33294 21310 33346
rect 21362 33294 21374 33346
rect 24546 33294 24558 33346
rect 24610 33294 24622 33346
rect 29922 33294 29934 33346
rect 29986 33294 29998 33346
rect 33842 33294 33854 33346
rect 33906 33294 33918 33346
rect 34402 33294 34414 33346
rect 34466 33294 34478 33346
rect 34738 33294 34750 33346
rect 34802 33294 34814 33346
rect 37426 33294 37438 33346
rect 37490 33294 37502 33346
rect 38770 33294 38782 33346
rect 38834 33294 38846 33346
rect 41234 33294 41246 33346
rect 41298 33294 41310 33346
rect 12574 33282 12626 33294
rect 30382 33282 30434 33294
rect 38446 33282 38498 33294
rect 42702 33282 42754 33294
rect 43374 33346 43426 33358
rect 43586 33294 43598 33346
rect 43650 33294 43662 33346
rect 46162 33294 46174 33346
rect 46226 33294 46238 33346
rect 46722 33294 46734 33346
rect 46786 33294 46798 33346
rect 47058 33294 47070 33346
rect 47122 33294 47134 33346
rect 43374 33282 43426 33294
rect 2382 33234 2434 33246
rect 2382 33170 2434 33182
rect 5742 33234 5794 33246
rect 5742 33170 5794 33182
rect 6638 33234 6690 33246
rect 6638 33170 6690 33182
rect 9326 33234 9378 33246
rect 9326 33170 9378 33182
rect 9886 33234 9938 33246
rect 9886 33170 9938 33182
rect 10334 33234 10386 33246
rect 10334 33170 10386 33182
rect 12686 33234 12738 33246
rect 12686 33170 12738 33182
rect 13582 33234 13634 33246
rect 38334 33234 38386 33246
rect 14802 33182 14814 33234
rect 14866 33182 14878 33234
rect 16258 33182 16270 33234
rect 16322 33182 16334 33234
rect 18722 33182 18734 33234
rect 18786 33182 18798 33234
rect 21522 33182 21534 33234
rect 21586 33182 21598 33234
rect 21970 33182 21982 33234
rect 22034 33182 22046 33234
rect 39778 33182 39790 33234
rect 39842 33182 39854 33234
rect 41010 33182 41022 33234
rect 41074 33182 41086 33234
rect 41346 33182 41358 33234
rect 41410 33182 41422 33234
rect 13582 33170 13634 33182
rect 38334 33170 38386 33182
rect 9550 33122 9602 33134
rect 9550 33058 9602 33070
rect 10222 33122 10274 33134
rect 10222 33058 10274 33070
rect 10446 33122 10498 33134
rect 10446 33058 10498 33070
rect 10670 33122 10722 33134
rect 18398 33122 18450 33134
rect 17154 33070 17166 33122
rect 17218 33070 17230 33122
rect 10670 33058 10722 33070
rect 18398 33058 18450 33070
rect 19406 33122 19458 33134
rect 19406 33058 19458 33070
rect 19854 33122 19906 33134
rect 40126 33122 40178 33134
rect 34738 33070 34750 33122
rect 34802 33070 34814 33122
rect 19854 33058 19906 33070
rect 40126 33058 40178 33070
rect 42478 33122 42530 33134
rect 42478 33058 42530 33070
rect 42814 33122 42866 33134
rect 42814 33058 42866 33070
rect 42926 33122 42978 33134
rect 42926 33058 42978 33070
rect 45726 33122 45778 33134
rect 45726 33058 45778 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 1822 32786 1874 32798
rect 1822 32722 1874 32734
rect 4286 32786 4338 32798
rect 4286 32722 4338 32734
rect 4734 32786 4786 32798
rect 4734 32722 4786 32734
rect 8654 32786 8706 32798
rect 8654 32722 8706 32734
rect 9886 32786 9938 32798
rect 19630 32786 19682 32798
rect 12114 32734 12126 32786
rect 12178 32734 12190 32786
rect 14354 32734 14366 32786
rect 14418 32734 14430 32786
rect 9886 32722 9938 32734
rect 19630 32722 19682 32734
rect 21086 32786 21138 32798
rect 21086 32722 21138 32734
rect 22094 32786 22146 32798
rect 38558 32786 38610 32798
rect 28242 32734 28254 32786
rect 28306 32734 28318 32786
rect 34962 32734 34974 32786
rect 35026 32734 35038 32786
rect 22094 32722 22146 32734
rect 38558 32722 38610 32734
rect 39566 32786 39618 32798
rect 39566 32722 39618 32734
rect 41694 32786 41746 32798
rect 41694 32722 41746 32734
rect 3166 32674 3218 32686
rect 9550 32674 9602 32686
rect 8194 32622 8206 32674
rect 8258 32622 8270 32674
rect 3166 32610 3218 32622
rect 9550 32610 9602 32622
rect 11006 32674 11058 32686
rect 11006 32610 11058 32622
rect 15822 32674 15874 32686
rect 15822 32610 15874 32622
rect 17390 32674 17442 32686
rect 20414 32674 20466 32686
rect 19954 32622 19966 32674
rect 20018 32622 20030 32674
rect 17390 32610 17442 32622
rect 20414 32610 20466 32622
rect 20526 32674 20578 32686
rect 37214 32674 37266 32686
rect 30706 32622 30718 32674
rect 30770 32622 30782 32674
rect 33506 32622 33518 32674
rect 33570 32622 33582 32674
rect 20526 32610 20578 32622
rect 37214 32610 37266 32622
rect 38222 32674 38274 32686
rect 38222 32610 38274 32622
rect 38446 32674 38498 32686
rect 38446 32610 38498 32622
rect 39790 32674 39842 32686
rect 39790 32610 39842 32622
rect 40350 32674 40402 32686
rect 40350 32610 40402 32622
rect 40910 32674 40962 32686
rect 40910 32610 40962 32622
rect 41246 32674 41298 32686
rect 48190 32674 48242 32686
rect 46050 32622 46062 32674
rect 46114 32622 46126 32674
rect 41246 32610 41298 32622
rect 48190 32610 48242 32622
rect 2718 32562 2770 32574
rect 5630 32562 5682 32574
rect 2482 32510 2494 32562
rect 2546 32510 2558 32562
rect 2930 32510 2942 32562
rect 2994 32510 3006 32562
rect 2718 32498 2770 32510
rect 5630 32498 5682 32510
rect 6302 32562 6354 32574
rect 13806 32562 13858 32574
rect 7186 32510 7198 32562
rect 7250 32510 7262 32562
rect 7746 32510 7758 32562
rect 7810 32510 7822 32562
rect 12338 32510 12350 32562
rect 12402 32510 12414 32562
rect 6302 32498 6354 32510
rect 13806 32498 13858 32510
rect 14030 32562 14082 32574
rect 18846 32562 18898 32574
rect 17602 32510 17614 32562
rect 17666 32510 17678 32562
rect 14030 32498 14082 32510
rect 18846 32498 18898 32510
rect 21870 32562 21922 32574
rect 21870 32498 21922 32510
rect 22542 32562 22594 32574
rect 22542 32498 22594 32510
rect 22766 32562 22818 32574
rect 38894 32562 38946 32574
rect 23090 32510 23102 32562
rect 23154 32510 23166 32562
rect 25218 32510 25230 32562
rect 25282 32510 25294 32562
rect 31042 32510 31054 32562
rect 31106 32510 31118 32562
rect 32050 32510 32062 32562
rect 32114 32510 32126 32562
rect 33842 32510 33854 32562
rect 33906 32510 33918 32562
rect 34850 32510 34862 32562
rect 34914 32510 34926 32562
rect 37426 32510 37438 32562
rect 37490 32510 37502 32562
rect 47282 32510 47294 32562
rect 47346 32510 47358 32562
rect 22766 32498 22818 32510
rect 38894 32498 38946 32510
rect 3054 32450 3106 32462
rect 3054 32386 3106 32398
rect 3838 32450 3890 32462
rect 3838 32386 3890 32398
rect 5070 32450 5122 32462
rect 5070 32386 5122 32398
rect 6526 32450 6578 32462
rect 18510 32450 18562 32462
rect 7410 32398 7422 32450
rect 7474 32398 7486 32450
rect 6526 32386 6578 32398
rect 18510 32386 18562 32398
rect 21982 32450 22034 32462
rect 21982 32386 22034 32398
rect 22878 32450 22930 32462
rect 22878 32386 22930 32398
rect 24670 32450 24722 32462
rect 26002 32398 26014 32450
rect 26066 32398 26078 32450
rect 30034 32398 30046 32450
rect 30098 32398 30110 32450
rect 31938 32398 31950 32450
rect 32002 32398 32014 32450
rect 47058 32398 47070 32450
rect 47122 32398 47134 32450
rect 24670 32386 24722 32398
rect 11230 32338 11282 32350
rect 5954 32286 5966 32338
rect 6018 32286 6030 32338
rect 11230 32274 11282 32286
rect 11566 32338 11618 32350
rect 11566 32274 11618 32286
rect 16046 32338 16098 32350
rect 16046 32274 16098 32286
rect 16382 32338 16434 32350
rect 16382 32274 16434 32286
rect 18958 32338 19010 32350
rect 18958 32274 19010 32286
rect 20414 32338 20466 32350
rect 20414 32274 20466 32286
rect 31726 32338 31778 32350
rect 31726 32274 31778 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 42702 32002 42754 32014
rect 2706 31950 2718 32002
rect 2770 31950 2782 32002
rect 11442 31950 11454 32002
rect 11506 31950 11518 32002
rect 42702 31938 42754 31950
rect 41134 31890 41186 31902
rect 6402 31838 6414 31890
rect 6466 31838 6478 31890
rect 7298 31838 7310 31890
rect 7362 31838 7374 31890
rect 15698 31838 15710 31890
rect 15762 31838 15774 31890
rect 23314 31838 23326 31890
rect 23378 31838 23390 31890
rect 29250 31838 29262 31890
rect 29314 31838 29326 31890
rect 31714 31838 31726 31890
rect 31778 31838 31790 31890
rect 35634 31838 35646 31890
rect 35698 31838 35710 31890
rect 41134 31826 41186 31838
rect 41358 31890 41410 31902
rect 41358 31826 41410 31838
rect 42254 31890 42306 31902
rect 42254 31826 42306 31838
rect 2158 31778 2210 31790
rect 2158 31714 2210 31726
rect 2494 31778 2546 31790
rect 3838 31778 3890 31790
rect 10670 31778 10722 31790
rect 2818 31726 2830 31778
rect 2882 31726 2894 31778
rect 6626 31726 6638 31778
rect 6690 31726 6702 31778
rect 7410 31726 7422 31778
rect 7474 31726 7486 31778
rect 9314 31726 9326 31778
rect 9378 31726 9390 31778
rect 2494 31714 2546 31726
rect 3838 31714 3890 31726
rect 10670 31714 10722 31726
rect 10894 31778 10946 31790
rect 10894 31714 10946 31726
rect 14590 31778 14642 31790
rect 23550 31778 23602 31790
rect 34414 31778 34466 31790
rect 14914 31726 14926 31778
rect 14978 31726 14990 31778
rect 17378 31726 17390 31778
rect 17442 31726 17454 31778
rect 22082 31726 22094 31778
rect 22146 31726 22158 31778
rect 22642 31726 22654 31778
rect 22706 31726 22718 31778
rect 30706 31726 30718 31778
rect 30770 31726 30782 31778
rect 35522 31726 35534 31778
rect 35586 31726 35598 31778
rect 14590 31714 14642 31726
rect 23550 31714 23602 31726
rect 34414 31714 34466 31726
rect 1934 31666 1986 31678
rect 1934 31602 1986 31614
rect 4846 31666 4898 31678
rect 9550 31666 9602 31678
rect 7746 31614 7758 31666
rect 7810 31614 7822 31666
rect 4846 31602 4898 31614
rect 9550 31602 9602 31614
rect 11118 31666 11170 31678
rect 23886 31666 23938 31678
rect 16034 31614 16046 31666
rect 16098 31614 16110 31666
rect 18386 31614 18398 31666
rect 18450 31614 18462 31666
rect 11118 31602 11170 31614
rect 23886 31602 23938 31614
rect 28590 31666 28642 31678
rect 33294 31666 33346 31678
rect 29474 31614 29486 31666
rect 29538 31614 29550 31666
rect 28590 31602 28642 31614
rect 33294 31602 33346 31614
rect 34526 31666 34578 31678
rect 34526 31602 34578 31614
rect 35982 31666 36034 31678
rect 42590 31666 42642 31678
rect 39778 31614 39790 31666
rect 39842 31614 39854 31666
rect 35982 31602 36034 31614
rect 42590 31602 42642 31614
rect 3278 31554 3330 31566
rect 2594 31502 2606 31554
rect 2658 31502 2670 31554
rect 3278 31490 3330 31502
rect 4622 31554 4674 31566
rect 4622 31490 4674 31502
rect 4958 31554 5010 31566
rect 4958 31490 5010 31502
rect 5182 31554 5234 31566
rect 5182 31490 5234 31502
rect 5966 31554 6018 31566
rect 5966 31490 6018 31502
rect 9998 31554 10050 31566
rect 9998 31490 10050 31502
rect 11902 31554 11954 31566
rect 23774 31554 23826 31566
rect 12226 31502 12238 31554
rect 12290 31502 12302 31554
rect 11902 31490 11954 31502
rect 23774 31490 23826 31502
rect 32958 31554 33010 31566
rect 32958 31490 33010 31502
rect 34750 31554 34802 31566
rect 48190 31554 48242 31566
rect 40674 31502 40686 31554
rect 40738 31502 40750 31554
rect 41682 31502 41694 31554
rect 41746 31502 41758 31554
rect 34750 31490 34802 31502
rect 48190 31490 48242 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 23326 31218 23378 31230
rect 23326 31154 23378 31166
rect 25790 31218 25842 31230
rect 25790 31154 25842 31166
rect 27246 31218 27298 31230
rect 27246 31154 27298 31166
rect 7870 31106 7922 31118
rect 6850 31054 6862 31106
rect 6914 31054 6926 31106
rect 7870 31042 7922 31054
rect 8094 31106 8146 31118
rect 8094 31042 8146 31054
rect 10894 31106 10946 31118
rect 10894 31042 10946 31054
rect 11230 31106 11282 31118
rect 20750 31106 20802 31118
rect 17490 31054 17502 31106
rect 17554 31054 17566 31106
rect 11230 31042 11282 31054
rect 20750 31042 20802 31054
rect 21422 31106 21474 31118
rect 21422 31042 21474 31054
rect 27470 31106 27522 31118
rect 34414 31106 34466 31118
rect 29922 31054 29934 31106
rect 29986 31054 29998 31106
rect 32050 31054 32062 31106
rect 32114 31054 32126 31106
rect 27470 31042 27522 31054
rect 34414 31042 34466 31054
rect 42478 31106 42530 31118
rect 42478 31042 42530 31054
rect 8318 30994 8370 31006
rect 1698 30942 1710 30994
rect 1762 30942 1774 30994
rect 5506 30942 5518 30994
rect 5570 30942 5582 30994
rect 6402 30942 6414 30994
rect 6466 30942 6478 30994
rect 8318 30930 8370 30942
rect 8430 30994 8482 31006
rect 8430 30930 8482 30942
rect 9662 30994 9714 31006
rect 14030 30994 14082 31006
rect 9874 30942 9886 30994
rect 9938 30942 9950 30994
rect 12226 30942 12238 30994
rect 12290 30942 12302 30994
rect 13234 30942 13246 30994
rect 13298 30942 13310 30994
rect 9662 30930 9714 30942
rect 14030 30930 14082 30942
rect 14366 30994 14418 31006
rect 14366 30930 14418 30942
rect 14926 30994 14978 31006
rect 14926 30930 14978 30942
rect 16158 30994 16210 31006
rect 28814 30994 28866 31006
rect 17378 30942 17390 30994
rect 17442 30942 17454 30994
rect 18274 30942 18286 30994
rect 18338 30942 18350 30994
rect 20066 30942 20078 30994
rect 20130 30942 20142 30994
rect 21186 30942 21198 30994
rect 21250 30942 21262 30994
rect 23538 30942 23550 30994
rect 23602 30942 23614 30994
rect 25554 30942 25566 30994
rect 25618 30942 25630 30994
rect 28466 30942 28478 30994
rect 28530 30942 28542 30994
rect 16158 30930 16210 30942
rect 28814 30930 28866 30942
rect 29038 30994 29090 31006
rect 41806 30994 41858 31006
rect 30818 30942 30830 30994
rect 30882 30942 30894 30994
rect 31826 30942 31838 30994
rect 31890 30942 31902 30994
rect 36194 30942 36206 30994
rect 36258 30942 36270 30994
rect 36530 30942 36542 30994
rect 36594 30942 36606 30994
rect 37538 30942 37550 30994
rect 37602 30942 37614 30994
rect 37874 30942 37886 30994
rect 37938 30942 37950 30994
rect 38546 30942 38558 30994
rect 38610 30942 38622 30994
rect 41570 30942 41582 30994
rect 41634 30942 41646 30994
rect 29038 30930 29090 30942
rect 41806 30930 41858 30942
rect 4958 30882 5010 30894
rect 2482 30830 2494 30882
rect 2546 30830 2558 30882
rect 4610 30830 4622 30882
rect 4674 30830 4686 30882
rect 4958 30818 5010 30830
rect 10558 30882 10610 30894
rect 15374 30882 15426 30894
rect 40910 30882 40962 30894
rect 11778 30830 11790 30882
rect 11842 30830 11854 30882
rect 16706 30830 16718 30882
rect 16770 30830 16782 30882
rect 18050 30830 18062 30882
rect 18114 30830 18126 30882
rect 20514 30830 20526 30882
rect 20578 30830 20590 30882
rect 42578 30830 42590 30882
rect 42642 30830 42654 30882
rect 10558 30818 10610 30830
rect 15374 30818 15426 30830
rect 40910 30818 40962 30830
rect 16382 30770 16434 30782
rect 8866 30718 8878 30770
rect 8930 30718 8942 30770
rect 16382 30706 16434 30718
rect 29150 30770 29202 30782
rect 29150 30706 29202 30718
rect 34526 30770 34578 30782
rect 42254 30770 42306 30782
rect 35298 30718 35310 30770
rect 35362 30718 35374 30770
rect 34526 30706 34578 30718
rect 42254 30706 42306 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 14142 30322 14194 30334
rect 16046 30322 16098 30334
rect 4498 30270 4510 30322
rect 4562 30270 4574 30322
rect 6626 30270 6638 30322
rect 6690 30270 6702 30322
rect 15138 30270 15150 30322
rect 15202 30270 15214 30322
rect 14142 30258 14194 30270
rect 16046 30258 16098 30270
rect 16382 30322 16434 30334
rect 29934 30322 29986 30334
rect 16594 30270 16606 30322
rect 16658 30270 16670 30322
rect 18050 30270 18062 30322
rect 18114 30270 18126 30322
rect 20738 30270 20750 30322
rect 20802 30270 20814 30322
rect 16382 30258 16434 30270
rect 29934 30258 29986 30270
rect 1934 30210 1986 30222
rect 1934 30146 1986 30158
rect 2942 30210 2994 30222
rect 12910 30210 12962 30222
rect 4386 30158 4398 30210
rect 4450 30158 4462 30210
rect 5170 30158 5182 30210
rect 5234 30158 5246 30210
rect 6514 30158 6526 30210
rect 6578 30158 6590 30210
rect 8530 30158 8542 30210
rect 8594 30158 8606 30210
rect 10098 30158 10110 30210
rect 10162 30158 10174 30210
rect 12114 30158 12126 30210
rect 12178 30158 12190 30210
rect 14814 30210 14866 30222
rect 27246 30210 27298 30222
rect 2942 30146 2994 30158
rect 12910 30146 12962 30158
rect 14478 30154 14530 30166
rect 2606 30098 2658 30110
rect 12574 30098 12626 30110
rect 4274 30046 4286 30098
rect 4338 30046 4350 30098
rect 7746 30046 7758 30098
rect 7810 30046 7822 30098
rect 8082 30046 8094 30098
rect 8146 30046 8158 30098
rect 11330 30046 11342 30098
rect 11394 30046 11406 30098
rect 2606 30034 2658 30046
rect 12574 30034 12626 30046
rect 12686 30098 12738 30110
rect 15586 30158 15598 30210
rect 15650 30158 15662 30210
rect 16706 30158 16718 30210
rect 16770 30158 16782 30210
rect 19394 30158 19406 30210
rect 19458 30158 19470 30210
rect 21410 30158 21422 30210
rect 21474 30158 21486 30210
rect 23538 30158 23550 30210
rect 23602 30158 23614 30210
rect 14814 30146 14866 30158
rect 27246 30146 27298 30158
rect 27582 30210 27634 30222
rect 28478 30210 28530 30222
rect 35422 30210 35474 30222
rect 28242 30158 28254 30210
rect 28306 30158 28318 30210
rect 31938 30158 31950 30210
rect 32002 30158 32014 30210
rect 32610 30158 32622 30210
rect 32674 30158 32686 30210
rect 33058 30158 33070 30210
rect 33122 30158 33134 30210
rect 27582 30146 27634 30158
rect 28478 30146 28530 30158
rect 35422 30146 35474 30158
rect 36990 30210 37042 30222
rect 36990 30146 37042 30158
rect 37102 30210 37154 30222
rect 37426 30158 37438 30210
rect 37490 30158 37502 30210
rect 40338 30158 40350 30210
rect 40402 30158 40414 30210
rect 41122 30158 41134 30210
rect 41186 30158 41198 30210
rect 41794 30158 41806 30210
rect 41858 30158 41870 30210
rect 42354 30158 42366 30210
rect 42418 30158 42430 30210
rect 37102 30146 37154 30158
rect 14478 30090 14530 30102
rect 17278 30098 17330 30110
rect 12686 30034 12738 30046
rect 17278 30034 17330 30046
rect 17390 30098 17442 30110
rect 29262 30098 29314 30110
rect 18162 30046 18174 30098
rect 18226 30046 18238 30098
rect 21746 30046 21758 30098
rect 21810 30046 21822 30098
rect 22642 30046 22654 30098
rect 22706 30046 22718 30098
rect 23202 30046 23214 30098
rect 23266 30046 23278 30098
rect 17390 30034 17442 30046
rect 29262 30034 29314 30046
rect 29374 30098 29426 30110
rect 35870 30098 35922 30110
rect 32050 30046 32062 30098
rect 32114 30046 32126 30098
rect 29374 30034 29426 30046
rect 35870 30034 35922 30046
rect 36094 30098 36146 30110
rect 36094 30034 36146 30046
rect 40574 30098 40626 30110
rect 40574 30034 40626 30046
rect 40686 30098 40738 30110
rect 43934 30098 43986 30110
rect 41570 30046 41582 30098
rect 41634 30046 41646 30098
rect 40686 30034 40738 30046
rect 43934 30034 43986 30046
rect 2270 29986 2322 29998
rect 2270 29922 2322 29934
rect 3502 29986 3554 29998
rect 3502 29922 3554 29934
rect 5742 29986 5794 29998
rect 5742 29922 5794 29934
rect 9662 29986 9714 29998
rect 9662 29922 9714 29934
rect 14590 29986 14642 29998
rect 14590 29922 14642 29934
rect 17614 29986 17666 29998
rect 29038 29986 29090 29998
rect 21858 29934 21870 29986
rect 21922 29934 21934 29986
rect 22754 29934 22766 29986
rect 22818 29934 22830 29986
rect 17614 29922 17666 29934
rect 29038 29922 29090 29934
rect 35982 29986 36034 29998
rect 35982 29922 36034 29934
rect 38446 29986 38498 29998
rect 38446 29922 38498 29934
rect 40014 29986 40066 29998
rect 44046 29986 44098 29998
rect 42466 29934 42478 29986
rect 42530 29934 42542 29986
rect 40014 29922 40066 29934
rect 44046 29922 44098 29934
rect 44270 29986 44322 29998
rect 44270 29922 44322 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 5406 29650 5458 29662
rect 5406 29586 5458 29598
rect 5966 29650 6018 29662
rect 5966 29586 6018 29598
rect 7534 29650 7586 29662
rect 7534 29586 7586 29598
rect 7982 29650 8034 29662
rect 7982 29586 8034 29598
rect 8990 29650 9042 29662
rect 8990 29586 9042 29598
rect 12014 29650 12066 29662
rect 12014 29586 12066 29598
rect 12574 29650 12626 29662
rect 12574 29586 12626 29598
rect 20638 29650 20690 29662
rect 20638 29586 20690 29598
rect 24670 29650 24722 29662
rect 39566 29650 39618 29662
rect 30034 29598 30046 29650
rect 30098 29598 30110 29650
rect 24670 29586 24722 29598
rect 39566 29586 39618 29598
rect 40350 29650 40402 29662
rect 40350 29586 40402 29598
rect 41246 29650 41298 29662
rect 47506 29598 47518 29650
rect 47570 29598 47582 29650
rect 41246 29586 41298 29598
rect 5630 29538 5682 29550
rect 5630 29474 5682 29486
rect 5742 29538 5794 29550
rect 14702 29538 14754 29550
rect 11218 29486 11230 29538
rect 11282 29486 11294 29538
rect 5742 29474 5794 29486
rect 14702 29474 14754 29486
rect 14814 29538 14866 29550
rect 14814 29474 14866 29486
rect 18622 29538 18674 29550
rect 18622 29474 18674 29486
rect 18846 29538 18898 29550
rect 18846 29474 18898 29486
rect 21758 29538 21810 29550
rect 32510 29538 32562 29550
rect 39118 29538 39170 29550
rect 27346 29486 27358 29538
rect 27410 29486 27422 29538
rect 28242 29486 28254 29538
rect 28306 29486 28318 29538
rect 36418 29486 36430 29538
rect 36482 29486 36494 29538
rect 38322 29486 38334 29538
rect 38386 29486 38398 29538
rect 21758 29474 21810 29486
rect 32510 29474 32562 29486
rect 39118 29474 39170 29486
rect 41358 29538 41410 29550
rect 41358 29474 41410 29486
rect 42590 29538 42642 29550
rect 45278 29538 45330 29550
rect 43362 29486 43374 29538
rect 43426 29486 43438 29538
rect 45938 29486 45950 29538
rect 46002 29486 46014 29538
rect 42590 29474 42642 29486
rect 45278 29474 45330 29486
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 2270 29426 2322 29438
rect 2270 29362 2322 29374
rect 9550 29426 9602 29438
rect 9550 29362 9602 29374
rect 9774 29426 9826 29438
rect 9774 29362 9826 29374
rect 10446 29426 10498 29438
rect 10446 29362 10498 29374
rect 10670 29426 10722 29438
rect 10670 29362 10722 29374
rect 10894 29426 10946 29438
rect 10894 29362 10946 29374
rect 11902 29426 11954 29438
rect 11902 29362 11954 29374
rect 12238 29426 12290 29438
rect 12238 29362 12290 29374
rect 22094 29426 22146 29438
rect 31614 29426 31666 29438
rect 40910 29426 40962 29438
rect 25442 29374 25454 29426
rect 25506 29374 25518 29426
rect 26786 29374 26798 29426
rect 26850 29374 26862 29426
rect 29698 29374 29710 29426
rect 29762 29374 29774 29426
rect 31938 29374 31950 29426
rect 32002 29374 32014 29426
rect 37314 29374 37326 29426
rect 37378 29374 37390 29426
rect 22094 29362 22146 29374
rect 31614 29362 31666 29374
rect 40910 29362 40962 29374
rect 41470 29426 41522 29438
rect 41470 29362 41522 29374
rect 42702 29426 42754 29438
rect 43922 29374 43934 29426
rect 43986 29374 43998 29426
rect 44594 29374 44606 29426
rect 44658 29374 44670 29426
rect 47170 29374 47182 29426
rect 47234 29374 47246 29426
rect 42702 29362 42754 29374
rect 4846 29314 4898 29326
rect 4846 29250 4898 29262
rect 15374 29314 15426 29326
rect 18834 29262 18846 29314
rect 18898 29262 18910 29314
rect 25890 29262 25902 29314
rect 25954 29262 25966 29314
rect 28018 29262 28030 29314
rect 28082 29262 28094 29314
rect 35858 29262 35870 29314
rect 35922 29262 35934 29314
rect 45714 29262 45726 29314
rect 45778 29262 45790 29314
rect 15374 29250 15426 29262
rect 9998 29202 10050 29214
rect 9998 29138 10050 29150
rect 14814 29202 14866 29214
rect 14814 29138 14866 29150
rect 39006 29202 39058 29214
rect 39006 29138 39058 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 10782 28866 10834 28878
rect 33742 28866 33794 28878
rect 27570 28814 27582 28866
rect 27634 28814 27646 28866
rect 10782 28802 10834 28814
rect 33742 28802 33794 28814
rect 35534 28866 35586 28878
rect 35534 28802 35586 28814
rect 39454 28866 39506 28878
rect 39454 28802 39506 28814
rect 40462 28866 40514 28878
rect 47058 28814 47070 28866
rect 47122 28814 47134 28866
rect 40462 28802 40514 28814
rect 12014 28754 12066 28766
rect 2482 28702 2494 28754
rect 2546 28702 2558 28754
rect 4610 28702 4622 28754
rect 4674 28702 4686 28754
rect 12014 28690 12066 28702
rect 17054 28754 17106 28766
rect 17054 28690 17106 28702
rect 18510 28754 18562 28766
rect 18510 28690 18562 28702
rect 20190 28754 20242 28766
rect 27022 28754 27074 28766
rect 24210 28702 24222 28754
rect 24274 28702 24286 28754
rect 20190 28690 20242 28702
rect 27022 28690 27074 28702
rect 27470 28754 27522 28766
rect 40238 28754 40290 28766
rect 38658 28702 38670 28754
rect 38722 28702 38734 28754
rect 27470 28690 27522 28702
rect 40238 28690 40290 28702
rect 41246 28754 41298 28766
rect 41246 28690 41298 28702
rect 43486 28754 43538 28766
rect 45278 28754 45330 28766
rect 43698 28702 43710 28754
rect 43762 28702 43774 28754
rect 46610 28702 46622 28754
rect 46674 28702 46686 28754
rect 43486 28690 43538 28702
rect 45278 28690 45330 28702
rect 5070 28642 5122 28654
rect 11230 28642 11282 28654
rect 1698 28590 1710 28642
rect 1762 28590 1774 28642
rect 5730 28590 5742 28642
rect 5794 28590 5806 28642
rect 9538 28590 9550 28642
rect 9602 28590 9614 28642
rect 5070 28578 5122 28590
rect 11230 28578 11282 28590
rect 14590 28642 14642 28654
rect 14590 28578 14642 28590
rect 18846 28642 18898 28654
rect 18846 28578 18898 28590
rect 18958 28642 19010 28654
rect 18958 28578 19010 28590
rect 19182 28642 19234 28654
rect 19182 28578 19234 28590
rect 19294 28642 19346 28654
rect 20414 28642 20466 28654
rect 19842 28590 19854 28642
rect 19906 28590 19918 28642
rect 19294 28578 19346 28590
rect 20414 28578 20466 28590
rect 21534 28642 21586 28654
rect 44718 28642 44770 28654
rect 22642 28590 22654 28642
rect 22706 28590 22718 28642
rect 25442 28590 25454 28642
rect 25506 28590 25518 28642
rect 25778 28590 25790 28642
rect 25842 28590 25854 28642
rect 27570 28590 27582 28642
rect 27634 28590 27646 28642
rect 28690 28590 28702 28642
rect 28754 28590 28766 28642
rect 38546 28590 38558 28642
rect 38610 28590 38622 28642
rect 46722 28590 46734 28642
rect 46786 28590 46798 28642
rect 21534 28578 21586 28590
rect 44718 28578 44770 28590
rect 10670 28530 10722 28542
rect 10098 28478 10110 28530
rect 10162 28478 10174 28530
rect 10670 28466 10722 28478
rect 10782 28530 10834 28542
rect 14702 28530 14754 28542
rect 11554 28478 11566 28530
rect 11618 28478 11630 28530
rect 10782 28466 10834 28478
rect 14702 28466 14754 28478
rect 16494 28530 16546 28542
rect 16494 28466 16546 28478
rect 16606 28530 16658 28542
rect 16606 28466 16658 28478
rect 22094 28530 22146 28542
rect 22094 28466 22146 28478
rect 22430 28530 22482 28542
rect 22430 28466 22482 28478
rect 32622 28530 32674 28542
rect 32622 28466 32674 28478
rect 33630 28530 33682 28542
rect 33630 28466 33682 28478
rect 33742 28530 33794 28542
rect 33742 28466 33794 28478
rect 35198 28530 35250 28542
rect 35198 28466 35250 28478
rect 35422 28530 35474 28542
rect 35422 28466 35474 28478
rect 35870 28530 35922 28542
rect 35870 28466 35922 28478
rect 35982 28530 36034 28542
rect 35982 28466 36034 28478
rect 37326 28530 37378 28542
rect 37326 28466 37378 28478
rect 37662 28530 37714 28542
rect 37662 28466 37714 28478
rect 39006 28530 39058 28542
rect 39006 28466 39058 28478
rect 39342 28530 39394 28542
rect 39342 28466 39394 28478
rect 45166 28530 45218 28542
rect 45166 28466 45218 28478
rect 45390 28530 45442 28542
rect 45390 28466 45442 28478
rect 48190 28530 48242 28542
rect 48190 28466 48242 28478
rect 5742 28418 5794 28430
rect 14926 28418 14978 28430
rect 9762 28366 9774 28418
rect 9826 28366 9838 28418
rect 5742 28354 5794 28366
rect 14926 28354 14978 28366
rect 16270 28418 16322 28430
rect 16270 28354 16322 28366
rect 32734 28418 32786 28430
rect 32734 28354 32786 28366
rect 32958 28418 33010 28430
rect 32958 28354 33010 28366
rect 36206 28418 36258 28430
rect 36206 28354 36258 28366
rect 39454 28418 39506 28430
rect 43710 28418 43762 28430
rect 40786 28366 40798 28418
rect 40850 28366 40862 28418
rect 39454 28354 39506 28366
rect 43710 28354 43762 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 3390 28082 3442 28094
rect 2482 28030 2494 28082
rect 2546 28030 2558 28082
rect 3390 28018 3442 28030
rect 8542 28082 8594 28094
rect 8542 28018 8594 28030
rect 11566 28082 11618 28094
rect 11566 28018 11618 28030
rect 12350 28082 12402 28094
rect 12350 28018 12402 28030
rect 12574 28082 12626 28094
rect 12574 28018 12626 28030
rect 25902 28082 25954 28094
rect 25902 28018 25954 28030
rect 33182 28082 33234 28094
rect 33182 28018 33234 28030
rect 40238 28082 40290 28094
rect 40238 28018 40290 28030
rect 46510 28082 46562 28094
rect 46510 28018 46562 28030
rect 8878 27970 8930 27982
rect 8878 27906 8930 27918
rect 8990 27970 9042 27982
rect 11342 27970 11394 27982
rect 10098 27918 10110 27970
rect 10162 27918 10174 27970
rect 8990 27906 9042 27918
rect 11342 27906 11394 27918
rect 11678 27970 11730 27982
rect 11678 27906 11730 27918
rect 14478 27970 14530 27982
rect 14478 27906 14530 27918
rect 20414 27970 20466 27982
rect 20414 27906 20466 27918
rect 20638 27970 20690 27982
rect 25678 27970 25730 27982
rect 21522 27918 21534 27970
rect 21586 27918 21598 27970
rect 23090 27918 23102 27970
rect 23154 27918 23166 27970
rect 20638 27906 20690 27918
rect 25678 27906 25730 27918
rect 26014 27970 26066 27982
rect 26014 27906 26066 27918
rect 27582 27970 27634 27982
rect 27582 27906 27634 27918
rect 29710 27970 29762 27982
rect 29710 27906 29762 27918
rect 33070 27970 33122 27982
rect 33954 27918 33966 27970
rect 34018 27918 34030 27970
rect 36082 27918 36094 27970
rect 36146 27918 36158 27970
rect 37538 27918 37550 27970
rect 37602 27918 37614 27970
rect 39778 27918 39790 27970
rect 39842 27918 39854 27970
rect 33070 27906 33122 27918
rect 2942 27858 2994 27870
rect 2258 27806 2270 27858
rect 2322 27806 2334 27858
rect 2942 27794 2994 27806
rect 8654 27858 8706 27870
rect 10446 27858 10498 27870
rect 9874 27806 9886 27858
rect 9938 27806 9950 27858
rect 8654 27794 8706 27806
rect 10446 27794 10498 27806
rect 11006 27858 11058 27870
rect 11006 27794 11058 27806
rect 11790 27858 11842 27870
rect 14814 27858 14866 27870
rect 19406 27858 19458 27870
rect 26126 27858 26178 27870
rect 28478 27858 28530 27870
rect 40350 27858 40402 27870
rect 12002 27806 12014 27858
rect 12066 27806 12078 27858
rect 12898 27806 12910 27858
rect 12962 27806 12974 27858
rect 15810 27806 15822 27858
rect 15874 27806 15886 27858
rect 16482 27806 16494 27858
rect 16546 27806 16558 27858
rect 19058 27806 19070 27858
rect 19122 27806 19134 27858
rect 21858 27806 21870 27858
rect 21922 27806 21934 27858
rect 28018 27806 28030 27858
rect 28082 27806 28094 27858
rect 30146 27806 30158 27858
rect 30210 27806 30222 27858
rect 34962 27806 34974 27858
rect 35026 27806 35038 27858
rect 35746 27806 35758 27858
rect 35810 27806 35822 27858
rect 38546 27806 38558 27858
rect 38610 27806 38622 27858
rect 11790 27794 11842 27806
rect 14814 27794 14866 27806
rect 19406 27794 19458 27806
rect 26126 27794 26178 27806
rect 28478 27794 28530 27806
rect 40350 27794 40402 27806
rect 46622 27858 46674 27870
rect 46622 27794 46674 27806
rect 1822 27746 1874 27758
rect 1822 27682 1874 27694
rect 12462 27746 12514 27758
rect 12462 27682 12514 27694
rect 15710 27746 15762 27758
rect 20526 27746 20578 27758
rect 19842 27694 19854 27746
rect 19906 27694 19918 27746
rect 15710 27682 15762 27694
rect 20526 27682 20578 27694
rect 23438 27746 23490 27758
rect 23438 27682 23490 27694
rect 23774 27746 23826 27758
rect 30594 27694 30606 27746
rect 30658 27694 30670 27746
rect 36978 27694 36990 27746
rect 37042 27694 37054 27746
rect 23774 27682 23826 27694
rect 16382 27634 16434 27646
rect 16382 27570 16434 27582
rect 18062 27634 18114 27646
rect 18062 27570 18114 27582
rect 23998 27634 24050 27646
rect 23998 27570 24050 27582
rect 24334 27634 24386 27646
rect 24334 27570 24386 27582
rect 33182 27634 33234 27646
rect 33182 27570 33234 27582
rect 40238 27634 40290 27646
rect 40238 27570 40290 27582
rect 46510 27634 46562 27646
rect 46510 27570 46562 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 21870 27298 21922 27310
rect 37662 27298 37714 27310
rect 41246 27298 41298 27310
rect 18386 27246 18398 27298
rect 18450 27246 18462 27298
rect 19170 27246 19182 27298
rect 19234 27295 19246 27298
rect 19842 27295 19854 27298
rect 19234 27249 19854 27295
rect 19234 27246 19246 27249
rect 19842 27246 19854 27249
rect 19906 27246 19918 27298
rect 35298 27246 35310 27298
rect 35362 27246 35374 27298
rect 37986 27246 37998 27298
rect 38050 27246 38062 27298
rect 21870 27234 21922 27246
rect 37662 27234 37714 27246
rect 41246 27234 41298 27246
rect 6750 27186 6802 27198
rect 2146 27134 2158 27186
rect 2210 27134 2222 27186
rect 6750 27122 6802 27134
rect 8878 27186 8930 27198
rect 8878 27122 8930 27134
rect 12910 27186 12962 27198
rect 19406 27186 19458 27198
rect 17714 27134 17726 27186
rect 17778 27134 17790 27186
rect 12910 27122 12962 27134
rect 19406 27122 19458 27134
rect 19966 27186 20018 27198
rect 31950 27186 32002 27198
rect 20626 27134 20638 27186
rect 20690 27134 20702 27186
rect 22754 27134 22766 27186
rect 22818 27134 22830 27186
rect 25554 27134 25566 27186
rect 25618 27134 25630 27186
rect 31042 27134 31054 27186
rect 31106 27134 31118 27186
rect 35522 27134 35534 27186
rect 35586 27134 35598 27186
rect 19966 27122 20018 27134
rect 31950 27122 32002 27134
rect 3278 27074 3330 27086
rect 12350 27074 12402 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 8418 27022 8430 27074
rect 8482 27022 8494 27074
rect 3278 27010 3330 27022
rect 12350 27010 12402 27022
rect 12798 27074 12850 27086
rect 12798 27010 12850 27022
rect 13582 27074 13634 27086
rect 21646 27074 21698 27086
rect 28254 27074 28306 27086
rect 37438 27074 37490 27086
rect 13794 27022 13806 27074
rect 13858 27022 13870 27074
rect 15922 27022 15934 27074
rect 15986 27022 15998 27074
rect 17042 27022 17054 27074
rect 17106 27022 17118 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 20738 27022 20750 27074
rect 20802 27022 20814 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 30818 27022 30830 27074
rect 30882 27022 30894 27074
rect 31602 27022 31614 27074
rect 31666 27022 31678 27074
rect 32610 27022 32622 27074
rect 32674 27022 32686 27074
rect 33394 27022 33406 27074
rect 33458 27022 33470 27074
rect 35410 27022 35422 27074
rect 35474 27022 35486 27074
rect 36194 27022 36206 27074
rect 36258 27022 36270 27074
rect 38994 27022 39006 27074
rect 39058 27022 39070 27074
rect 39890 27022 39902 27074
rect 39954 27022 39966 27074
rect 13582 27010 13634 27022
rect 21646 27010 21698 27022
rect 28254 27010 28306 27022
rect 37438 27010 37490 27022
rect 2606 26962 2658 26974
rect 2606 26898 2658 26910
rect 2942 26962 2994 26974
rect 4062 26962 4114 26974
rect 3602 26910 3614 26962
rect 3666 26910 3678 26962
rect 2942 26898 2994 26910
rect 4062 26898 4114 26910
rect 5854 26962 5906 26974
rect 10334 26962 10386 26974
rect 7746 26910 7758 26962
rect 7810 26910 7822 26962
rect 8194 26910 8206 26962
rect 8258 26910 8270 26962
rect 5854 26898 5906 26910
rect 10334 26898 10386 26910
rect 10670 26962 10722 26974
rect 10670 26898 10722 26910
rect 11006 26962 11058 26974
rect 11006 26898 11058 26910
rect 12126 26962 12178 26974
rect 12126 26898 12178 26910
rect 14478 26962 14530 26974
rect 28142 26962 28194 26974
rect 45614 26962 45666 26974
rect 16930 26910 16942 26962
rect 16994 26910 17006 26962
rect 22978 26910 22990 26962
rect 23042 26910 23054 26962
rect 30258 26910 30270 26962
rect 30322 26910 30334 26962
rect 33842 26910 33854 26962
rect 33906 26910 33918 26962
rect 38770 26910 38782 26962
rect 38834 26910 38846 26962
rect 14478 26898 14530 26910
rect 28142 26898 28194 26910
rect 45614 26898 45666 26910
rect 45726 26962 45778 26974
rect 45726 26898 45778 26910
rect 6190 26850 6242 26862
rect 6190 26786 6242 26798
rect 9998 26850 10050 26862
rect 9998 26786 10050 26798
rect 12574 26850 12626 26862
rect 27694 26850 27746 26862
rect 16146 26798 16158 26850
rect 16210 26798 16222 26850
rect 22194 26798 22206 26850
rect 22258 26798 22270 26850
rect 12574 26786 12626 26798
rect 27694 26786 27746 26798
rect 27918 26850 27970 26862
rect 27918 26786 27970 26798
rect 45950 26850 46002 26862
rect 45950 26786 46002 26798
rect 48190 26850 48242 26862
rect 48190 26786 48242 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 14478 26514 14530 26526
rect 13794 26462 13806 26514
rect 13858 26462 13870 26514
rect 14478 26450 14530 26462
rect 22094 26514 22146 26526
rect 22094 26450 22146 26462
rect 30942 26514 30994 26526
rect 30942 26450 30994 26462
rect 31054 26514 31106 26526
rect 31054 26450 31106 26462
rect 31614 26514 31666 26526
rect 31614 26450 31666 26462
rect 31838 26514 31890 26526
rect 31838 26450 31890 26462
rect 38334 26514 38386 26526
rect 38334 26450 38386 26462
rect 12686 26402 12738 26414
rect 16270 26402 16322 26414
rect 28926 26402 28978 26414
rect 2706 26350 2718 26402
rect 2770 26350 2782 26402
rect 6402 26350 6414 26402
rect 6466 26350 6478 26402
rect 10098 26350 10110 26402
rect 10162 26350 10174 26402
rect 10882 26350 10894 26402
rect 10946 26350 10958 26402
rect 12450 26350 12462 26402
rect 12514 26350 12526 26402
rect 14130 26350 14142 26402
rect 14194 26350 14206 26402
rect 18946 26350 18958 26402
rect 19010 26350 19022 26402
rect 20850 26350 20862 26402
rect 20914 26350 20926 26402
rect 12686 26338 12738 26350
rect 16270 26338 16322 26350
rect 28926 26338 28978 26350
rect 31502 26402 31554 26414
rect 31502 26338 31554 26350
rect 33070 26402 33122 26414
rect 45154 26350 45166 26402
rect 45218 26350 45230 26402
rect 47394 26350 47406 26402
rect 47458 26350 47470 26402
rect 33070 26338 33122 26350
rect 8990 26290 9042 26302
rect 13246 26290 13298 26302
rect 2034 26238 2046 26290
rect 2098 26238 2110 26290
rect 5618 26238 5630 26290
rect 5682 26238 5694 26290
rect 9874 26238 9886 26290
rect 9938 26238 9950 26290
rect 8990 26226 9042 26238
rect 13246 26226 13298 26238
rect 13470 26290 13522 26302
rect 22430 26290 22482 26302
rect 23774 26290 23826 26302
rect 27694 26290 27746 26302
rect 15250 26238 15262 26290
rect 15314 26238 15326 26290
rect 20178 26238 20190 26290
rect 20242 26238 20254 26290
rect 23090 26238 23102 26290
rect 23154 26238 23166 26290
rect 23426 26238 23438 26290
rect 23490 26238 23502 26290
rect 23986 26238 23998 26290
rect 24050 26238 24062 26290
rect 13470 26226 13522 26238
rect 22430 26226 22482 26238
rect 23774 26226 23826 26238
rect 27694 26226 27746 26238
rect 28142 26290 28194 26302
rect 29038 26290 29090 26302
rect 28466 26238 28478 26290
rect 28530 26238 28542 26290
rect 28142 26226 28194 26238
rect 29038 26226 29090 26238
rect 29150 26290 29202 26302
rect 33506 26238 33518 26290
rect 33570 26238 33582 26290
rect 43698 26238 43710 26290
rect 43762 26238 43774 26290
rect 46274 26238 46286 26290
rect 46338 26238 46350 26290
rect 29150 26226 29202 26238
rect 5294 26178 5346 26190
rect 27134 26178 27186 26190
rect 44158 26178 44210 26190
rect 4834 26126 4846 26178
rect 4898 26126 4910 26178
rect 8530 26126 8542 26178
rect 8594 26126 8606 26178
rect 10546 26126 10558 26178
rect 10610 26126 10622 26178
rect 15138 26126 15150 26178
rect 15202 26126 15214 26178
rect 18498 26126 18510 26178
rect 18562 26126 18574 26178
rect 33842 26126 33854 26178
rect 33906 26126 33918 26178
rect 43362 26126 43374 26178
rect 43426 26126 43438 26178
rect 44818 26126 44830 26178
rect 44882 26126 44894 26178
rect 5294 26114 5346 26126
rect 27134 26114 27186 26126
rect 44158 26114 44210 26126
rect 16494 26066 16546 26078
rect 15810 26014 15822 26066
rect 15874 26014 15886 26066
rect 16494 26002 16546 26014
rect 16830 26066 16882 26078
rect 31166 26066 31218 26078
rect 24098 26014 24110 26066
rect 24162 26014 24174 26066
rect 27458 26014 27470 26066
rect 27522 26014 27534 26066
rect 16830 26002 16882 26014
rect 31166 26002 31218 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 14254 25730 14306 25742
rect 25778 25678 25790 25730
rect 25842 25678 25854 25730
rect 14254 25666 14306 25678
rect 5070 25618 5122 25630
rect 11790 25618 11842 25630
rect 16606 25618 16658 25630
rect 34078 25618 34130 25630
rect 4274 25566 4286 25618
rect 4338 25566 4350 25618
rect 7746 25566 7758 25618
rect 7810 25566 7822 25618
rect 9986 25566 9998 25618
rect 10050 25566 10062 25618
rect 15810 25566 15822 25618
rect 15874 25566 15886 25618
rect 18386 25566 18398 25618
rect 18450 25566 18462 25618
rect 27570 25566 27582 25618
rect 27634 25566 27646 25618
rect 32274 25566 32286 25618
rect 32338 25566 32350 25618
rect 5070 25554 5122 25566
rect 11790 25554 11842 25566
rect 16606 25554 16658 25566
rect 34078 25554 34130 25566
rect 37214 25618 37266 25630
rect 37214 25554 37266 25566
rect 43710 25618 43762 25630
rect 45838 25618 45890 25630
rect 45378 25566 45390 25618
rect 45442 25566 45454 25618
rect 43710 25554 43762 25566
rect 45838 25554 45890 25566
rect 5630 25506 5682 25518
rect 8094 25506 8146 25518
rect 12126 25506 12178 25518
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 5842 25454 5854 25506
rect 5906 25454 5918 25506
rect 6290 25454 6302 25506
rect 6354 25454 6366 25506
rect 7410 25454 7422 25506
rect 7474 25454 7486 25506
rect 8530 25454 8542 25506
rect 8594 25454 8606 25506
rect 9090 25454 9102 25506
rect 9154 25454 9166 25506
rect 5630 25442 5682 25454
rect 8094 25442 8146 25454
rect 12126 25442 12178 25454
rect 14142 25506 14194 25518
rect 14142 25442 14194 25454
rect 14702 25506 14754 25518
rect 16942 25506 16994 25518
rect 20750 25506 20802 25518
rect 16146 25454 16158 25506
rect 16210 25454 16222 25506
rect 18274 25454 18286 25506
rect 18338 25454 18350 25506
rect 14702 25442 14754 25454
rect 16942 25442 16994 25454
rect 20750 25442 20802 25454
rect 21534 25506 21586 25518
rect 25230 25506 25282 25518
rect 23314 25454 23326 25506
rect 23378 25454 23390 25506
rect 21534 25442 21586 25454
rect 25230 25442 25282 25454
rect 25454 25506 25506 25518
rect 42814 25506 42866 25518
rect 46398 25506 46450 25518
rect 28018 25454 28030 25506
rect 28082 25454 28094 25506
rect 28578 25454 28590 25506
rect 28642 25454 28654 25506
rect 32162 25454 32174 25506
rect 32226 25454 32238 25506
rect 41010 25454 41022 25506
rect 41074 25454 41086 25506
rect 41682 25454 41694 25506
rect 41746 25454 41758 25506
rect 43138 25454 43150 25506
rect 43202 25454 43214 25506
rect 45154 25454 45166 25506
rect 45218 25454 45230 25506
rect 25454 25442 25506 25454
rect 42814 25442 42866 25454
rect 46398 25442 46450 25454
rect 14814 25394 14866 25406
rect 14814 25330 14866 25342
rect 15038 25394 15090 25406
rect 15038 25330 15090 25342
rect 19070 25394 19122 25406
rect 19070 25330 19122 25342
rect 20414 25394 20466 25406
rect 20414 25330 20466 25342
rect 21422 25394 21474 25406
rect 21422 25330 21474 25342
rect 23102 25394 23154 25406
rect 32622 25394 32674 25406
rect 46286 25394 46338 25406
rect 27906 25342 27918 25394
rect 27970 25342 27982 25394
rect 40562 25342 40574 25394
rect 40626 25342 40638 25394
rect 23102 25330 23154 25342
rect 32622 25330 32674 25342
rect 46286 25330 46338 25342
rect 12238 25282 12290 25294
rect 12238 25218 12290 25230
rect 12462 25282 12514 25294
rect 12462 25218 12514 25230
rect 14254 25282 14306 25294
rect 21198 25282 21250 25294
rect 17266 25230 17278 25282
rect 17330 25230 17342 25282
rect 14254 25218 14306 25230
rect 21198 25218 21250 25230
rect 26462 25282 26514 25294
rect 26462 25218 26514 25230
rect 29262 25282 29314 25294
rect 29262 25218 29314 25230
rect 33966 25282 34018 25294
rect 46062 25282 46114 25294
rect 42130 25230 42142 25282
rect 42194 25230 42206 25282
rect 33966 25218 34018 25230
rect 46062 25218 46114 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 5294 24946 5346 24958
rect 5294 24882 5346 24894
rect 6862 24946 6914 24958
rect 18174 24946 18226 24958
rect 11106 24894 11118 24946
rect 11170 24894 11182 24946
rect 6862 24882 6914 24894
rect 18174 24882 18226 24894
rect 18398 24946 18450 24958
rect 18398 24882 18450 24894
rect 18958 24946 19010 24958
rect 18958 24882 19010 24894
rect 21310 24946 21362 24958
rect 21310 24882 21362 24894
rect 23550 24946 23602 24958
rect 32398 24946 32450 24958
rect 28690 24894 28702 24946
rect 28754 24894 28766 24946
rect 23550 24882 23602 24894
rect 32398 24882 32450 24894
rect 36878 24946 36930 24958
rect 36878 24882 36930 24894
rect 37886 24946 37938 24958
rect 37886 24882 37938 24894
rect 38446 24946 38498 24958
rect 38446 24882 38498 24894
rect 39118 24946 39170 24958
rect 39118 24882 39170 24894
rect 39566 24946 39618 24958
rect 39566 24882 39618 24894
rect 4734 24834 4786 24846
rect 4734 24770 4786 24782
rect 5182 24834 5234 24846
rect 6750 24834 6802 24846
rect 5842 24782 5854 24834
rect 5906 24782 5918 24834
rect 5182 24770 5234 24782
rect 6750 24770 6802 24782
rect 12798 24834 12850 24846
rect 19630 24834 19682 24846
rect 14690 24782 14702 24834
rect 14754 24782 14766 24834
rect 12798 24770 12850 24782
rect 19630 24770 19682 24782
rect 20862 24834 20914 24846
rect 20862 24770 20914 24782
rect 25230 24834 25282 24846
rect 31950 24834 32002 24846
rect 27122 24782 27134 24834
rect 27186 24782 27198 24834
rect 28802 24782 28814 24834
rect 28866 24782 28878 24834
rect 25230 24770 25282 24782
rect 31950 24770 32002 24782
rect 32286 24834 32338 24846
rect 37998 24834 38050 24846
rect 37426 24782 37438 24834
rect 37490 24782 37502 24834
rect 32286 24770 32338 24782
rect 37998 24770 38050 24782
rect 39454 24834 39506 24846
rect 39454 24770 39506 24782
rect 40014 24834 40066 24846
rect 40014 24770 40066 24782
rect 42254 24834 42306 24846
rect 43026 24782 43038 24834
rect 43090 24782 43102 24834
rect 42254 24770 42306 24782
rect 4846 24722 4898 24734
rect 7086 24722 7138 24734
rect 10782 24722 10834 24734
rect 18062 24722 18114 24734
rect 6066 24670 6078 24722
rect 6130 24670 6142 24722
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 8306 24670 8318 24722
rect 8370 24670 8382 24722
rect 14354 24670 14366 24722
rect 14418 24670 14430 24722
rect 4846 24658 4898 24670
rect 7086 24658 7138 24670
rect 10782 24658 10834 24670
rect 18062 24658 18114 24670
rect 19406 24722 19458 24734
rect 19406 24658 19458 24670
rect 20078 24722 20130 24734
rect 20078 24658 20130 24670
rect 20302 24722 20354 24734
rect 23214 24722 23266 24734
rect 31838 24722 31890 24734
rect 22978 24670 22990 24722
rect 23042 24670 23054 24722
rect 25442 24670 25454 24722
rect 25506 24670 25518 24722
rect 25890 24670 25902 24722
rect 25954 24670 25966 24722
rect 27570 24670 27582 24722
rect 27634 24670 27646 24722
rect 31490 24670 31502 24722
rect 31554 24670 31566 24722
rect 20302 24658 20354 24670
rect 23214 24658 23266 24670
rect 31838 24658 31890 24670
rect 32622 24722 32674 24734
rect 39790 24722 39842 24734
rect 43822 24722 43874 24734
rect 32946 24670 32958 24722
rect 33010 24670 33022 24722
rect 33954 24670 33966 24722
rect 34018 24670 34030 24722
rect 35410 24670 35422 24722
rect 35474 24670 35486 24722
rect 37202 24670 37214 24722
rect 37266 24670 37278 24722
rect 40338 24670 40350 24722
rect 40402 24670 40414 24722
rect 42466 24670 42478 24722
rect 42530 24670 42542 24722
rect 42914 24670 42926 24722
rect 42978 24670 42990 24722
rect 32622 24658 32674 24670
rect 39790 24658 39842 24670
rect 43822 24658 43874 24670
rect 44046 24722 44098 24734
rect 44718 24722 44770 24734
rect 44370 24670 44382 24722
rect 44434 24670 44446 24722
rect 44046 24658 44098 24670
rect 44718 24658 44770 24670
rect 45054 24722 45106 24734
rect 45054 24658 45106 24670
rect 45390 24722 45442 24734
rect 45390 24658 45442 24670
rect 19854 24610 19906 24622
rect 8194 24558 8206 24610
rect 8258 24558 8270 24610
rect 14578 24558 14590 24610
rect 14642 24558 14654 24610
rect 19058 24558 19070 24610
rect 19122 24558 19134 24610
rect 19854 24546 19906 24558
rect 29486 24610 29538 24622
rect 29486 24546 29538 24558
rect 29934 24610 29986 24622
rect 35870 24610 35922 24622
rect 45166 24610 45218 24622
rect 33618 24558 33630 24610
rect 33682 24558 33694 24610
rect 34962 24558 34974 24610
rect 35026 24558 35038 24610
rect 43138 24558 43150 24610
rect 43202 24558 43214 24610
rect 29934 24546 29986 24558
rect 35870 24546 35922 24558
rect 45166 24546 45218 24558
rect 4734 24498 4786 24510
rect 4734 24434 4786 24446
rect 5294 24498 5346 24510
rect 18734 24498 18786 24510
rect 37886 24498 37938 24510
rect 8306 24446 8318 24498
rect 8370 24446 8382 24498
rect 13794 24446 13806 24498
rect 13858 24446 13870 24498
rect 33730 24446 33742 24498
rect 33794 24446 33806 24498
rect 5294 24434 5346 24446
rect 18734 24434 18786 24446
rect 37886 24434 37938 24446
rect 40350 24498 40402 24510
rect 40350 24434 40402 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 43698 24110 43710 24162
rect 43762 24159 43774 24162
rect 44146 24159 44158 24162
rect 43762 24113 44158 24159
rect 43762 24110 43774 24113
rect 44146 24110 44158 24113
rect 44210 24110 44222 24162
rect 2270 24050 2322 24062
rect 2270 23986 2322 23998
rect 29150 24050 29202 24062
rect 39230 24050 39282 24062
rect 43710 24050 43762 24062
rect 29586 23998 29598 24050
rect 29650 23998 29662 24050
rect 31826 23998 31838 24050
rect 31890 23998 31902 24050
rect 36082 23998 36094 24050
rect 36146 23998 36158 24050
rect 41234 23998 41246 24050
rect 41298 23998 41310 24050
rect 43026 23998 43038 24050
rect 43090 23998 43102 24050
rect 29150 23986 29202 23998
rect 39230 23986 39282 23998
rect 43710 23986 43762 23998
rect 44158 24050 44210 24062
rect 44158 23986 44210 23998
rect 46734 24050 46786 24062
rect 46734 23986 46786 23998
rect 6414 23938 6466 23950
rect 6414 23874 6466 23886
rect 6750 23938 6802 23950
rect 6750 23874 6802 23886
rect 11454 23938 11506 23950
rect 11454 23874 11506 23886
rect 11678 23938 11730 23950
rect 11678 23874 11730 23886
rect 11902 23938 11954 23950
rect 11902 23874 11954 23886
rect 12126 23938 12178 23950
rect 20638 23938 20690 23950
rect 13570 23886 13582 23938
rect 13634 23886 13646 23938
rect 12126 23874 12178 23886
rect 20638 23874 20690 23886
rect 21534 23938 21586 23950
rect 21534 23874 21586 23886
rect 23214 23938 23266 23950
rect 32958 23938 33010 23950
rect 37326 23938 37378 23950
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 23874 23886 23886 23938
rect 23938 23886 23950 23938
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 26338 23886 26350 23938
rect 26402 23886 26414 23938
rect 29810 23886 29822 23938
rect 29874 23886 29886 23938
rect 31154 23886 31166 23938
rect 31218 23886 31230 23938
rect 31938 23886 31950 23938
rect 32002 23886 32014 23938
rect 34178 23886 34190 23938
rect 34242 23886 34254 23938
rect 35186 23886 35198 23938
rect 35250 23886 35262 23938
rect 23214 23874 23266 23886
rect 32958 23874 33010 23886
rect 37326 23874 37378 23886
rect 37662 23938 37714 23950
rect 37662 23874 37714 23886
rect 38334 23938 38386 23950
rect 38334 23874 38386 23886
rect 38894 23938 38946 23950
rect 39666 23886 39678 23938
rect 39730 23886 39742 23938
rect 40338 23886 40350 23938
rect 40402 23886 40414 23938
rect 40786 23886 40798 23938
rect 40850 23886 40862 23938
rect 41682 23886 41694 23938
rect 41746 23886 41758 23938
rect 42914 23886 42926 23938
rect 42978 23886 42990 23938
rect 46946 23886 46958 23938
rect 47010 23886 47022 23938
rect 38894 23874 38946 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 6638 23826 6690 23838
rect 6638 23762 6690 23774
rect 10222 23826 10274 23838
rect 10222 23762 10274 23774
rect 10670 23826 10722 23838
rect 10670 23762 10722 23774
rect 13806 23826 13858 23838
rect 20862 23826 20914 23838
rect 19954 23774 19966 23826
rect 20018 23774 20030 23826
rect 20178 23774 20190 23826
rect 20242 23774 20254 23826
rect 13806 23762 13858 23774
rect 20862 23762 20914 23774
rect 21310 23826 21362 23838
rect 21310 23762 21362 23774
rect 22878 23826 22930 23838
rect 37998 23826 38050 23838
rect 41918 23826 41970 23838
rect 25106 23774 25118 23826
rect 25170 23774 25182 23826
rect 25666 23774 25678 23826
rect 25730 23774 25742 23826
rect 32610 23774 32622 23826
rect 32674 23774 32686 23826
rect 33842 23774 33854 23826
rect 33906 23774 33918 23826
rect 40898 23774 40910 23826
rect 40962 23774 40974 23826
rect 42690 23774 42702 23826
rect 42754 23774 42766 23826
rect 48066 23774 48078 23826
rect 48130 23774 48142 23826
rect 22878 23762 22930 23774
rect 37998 23762 38050 23774
rect 41918 23762 41970 23774
rect 9662 23714 9714 23726
rect 9662 23650 9714 23662
rect 10894 23714 10946 23726
rect 10894 23650 10946 23662
rect 11006 23714 11058 23726
rect 11006 23650 11058 23662
rect 11118 23714 11170 23726
rect 11118 23650 11170 23662
rect 11342 23714 11394 23726
rect 22990 23714 23042 23726
rect 30942 23714 30994 23726
rect 21858 23662 21870 23714
rect 21922 23662 21934 23714
rect 26450 23662 26462 23714
rect 26514 23662 26526 23714
rect 11342 23650 11394 23662
rect 22990 23650 23042 23662
rect 30942 23650 30994 23662
rect 33070 23714 33122 23726
rect 33070 23650 33122 23662
rect 37662 23714 37714 23726
rect 37662 23650 37714 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 1822 23378 1874 23390
rect 1822 23314 1874 23326
rect 6862 23378 6914 23390
rect 6862 23314 6914 23326
rect 14702 23378 14754 23390
rect 14702 23314 14754 23326
rect 23998 23378 24050 23390
rect 23998 23314 24050 23326
rect 29822 23378 29874 23390
rect 29822 23314 29874 23326
rect 38782 23378 38834 23390
rect 38782 23314 38834 23326
rect 40798 23378 40850 23390
rect 40798 23314 40850 23326
rect 41022 23378 41074 23390
rect 41022 23314 41074 23326
rect 41582 23378 41634 23390
rect 41582 23314 41634 23326
rect 45838 23378 45890 23390
rect 45838 23314 45890 23326
rect 9550 23266 9602 23278
rect 14590 23266 14642 23278
rect 5842 23214 5854 23266
rect 5906 23214 5918 23266
rect 13346 23214 13358 23266
rect 13410 23214 13422 23266
rect 13906 23214 13918 23266
rect 13970 23214 13982 23266
rect 9550 23202 9602 23214
rect 14590 23202 14642 23214
rect 15486 23266 15538 23278
rect 15486 23202 15538 23214
rect 15598 23266 15650 23278
rect 15598 23202 15650 23214
rect 16158 23266 16210 23278
rect 22878 23266 22930 23278
rect 19282 23214 19294 23266
rect 19346 23214 19358 23266
rect 21298 23214 21310 23266
rect 21362 23214 21374 23266
rect 16158 23202 16210 23214
rect 22878 23202 22930 23214
rect 23886 23266 23938 23278
rect 29710 23266 29762 23278
rect 41134 23266 41186 23278
rect 26114 23214 26126 23266
rect 26178 23214 26190 23266
rect 35522 23214 35534 23266
rect 35586 23214 35598 23266
rect 38098 23214 38110 23266
rect 38162 23214 38174 23266
rect 23886 23202 23938 23214
rect 29710 23202 29762 23214
rect 41134 23202 41186 23214
rect 15822 23154 15874 23166
rect 27582 23154 27634 23166
rect 29150 23154 29202 23166
rect 4722 23102 4734 23154
rect 4786 23102 4798 23154
rect 11778 23102 11790 23154
rect 11842 23102 11854 23154
rect 12786 23102 12798 23154
rect 12850 23102 12862 23154
rect 14242 23102 14254 23154
rect 14306 23102 14318 23154
rect 21410 23102 21422 23154
rect 21474 23102 21486 23154
rect 22306 23102 22318 23154
rect 22370 23102 22382 23154
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 25330 23102 25342 23154
rect 25394 23102 25406 23154
rect 26674 23102 26686 23154
rect 26738 23102 26750 23154
rect 27234 23102 27246 23154
rect 27298 23102 27310 23154
rect 28466 23102 28478 23154
rect 28530 23102 28542 23154
rect 15822 23090 15874 23102
rect 27582 23090 27634 23102
rect 29150 23090 29202 23102
rect 30046 23154 30098 23166
rect 45726 23154 45778 23166
rect 33954 23102 33966 23154
rect 34018 23102 34030 23154
rect 37090 23102 37102 23154
rect 37154 23102 37166 23154
rect 39330 23102 39342 23154
rect 39394 23102 39406 23154
rect 39666 23102 39678 23154
rect 39730 23102 39742 23154
rect 40226 23102 40238 23154
rect 40290 23102 40302 23154
rect 30046 23090 30098 23102
rect 45726 23090 45778 23102
rect 4062 23042 4114 23054
rect 13022 23042 13074 23054
rect 25790 23042 25842 23054
rect 6178 22990 6190 23042
rect 6242 22990 6254 23042
rect 12226 22990 12238 23042
rect 12290 22990 12302 23042
rect 20290 22990 20302 23042
rect 20354 22990 20366 23042
rect 26226 22990 26238 23042
rect 26290 22990 26302 23042
rect 28130 22990 28142 23042
rect 28194 22990 28206 23042
rect 34066 22990 34078 23042
rect 34130 22990 34142 23042
rect 35298 22990 35310 23042
rect 35362 22990 35374 23042
rect 4062 22978 4114 22990
rect 13022 22978 13074 22990
rect 25790 22978 25842 22990
rect 14702 22930 14754 22942
rect 45838 22930 45890 22942
rect 10546 22878 10558 22930
rect 10610 22878 10622 22930
rect 12114 22878 12126 22930
rect 12178 22878 12190 22930
rect 34738 22878 34750 22930
rect 34802 22878 34814 22930
rect 39554 22878 39566 22930
rect 39618 22878 39630 22930
rect 14702 22866 14754 22878
rect 45838 22866 45890 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 15710 22594 15762 22606
rect 42578 22542 42590 22594
rect 42642 22542 42654 22594
rect 15710 22530 15762 22542
rect 11790 22482 11842 22494
rect 8530 22430 8542 22482
rect 8594 22430 8606 22482
rect 11790 22418 11842 22430
rect 12910 22482 12962 22494
rect 15038 22482 15090 22494
rect 14690 22430 14702 22482
rect 14754 22430 14766 22482
rect 12910 22418 12962 22430
rect 15038 22418 15090 22430
rect 15486 22482 15538 22494
rect 15486 22418 15538 22430
rect 19406 22482 19458 22494
rect 20302 22482 20354 22494
rect 25902 22482 25954 22494
rect 19730 22430 19742 22482
rect 19794 22430 19806 22482
rect 22082 22430 22094 22482
rect 22146 22430 22158 22482
rect 19406 22418 19458 22430
rect 20302 22418 20354 22430
rect 25902 22418 25954 22430
rect 29262 22482 29314 22494
rect 29262 22418 29314 22430
rect 36990 22482 37042 22494
rect 38446 22482 38498 22494
rect 40574 22482 40626 22494
rect 37426 22430 37438 22482
rect 37490 22430 37502 22482
rect 40002 22430 40014 22482
rect 40066 22430 40078 22482
rect 36990 22418 37042 22430
rect 38446 22418 38498 22430
rect 40574 22418 40626 22430
rect 41022 22482 41074 22494
rect 41022 22418 41074 22430
rect 42254 22482 42306 22494
rect 42254 22418 42306 22430
rect 45502 22482 45554 22494
rect 45938 22430 45950 22482
rect 46002 22430 46014 22482
rect 45502 22418 45554 22430
rect 7086 22370 7138 22382
rect 7086 22306 7138 22318
rect 7422 22370 7474 22382
rect 7422 22306 7474 22318
rect 7758 22370 7810 22382
rect 9326 22370 9378 22382
rect 8418 22318 8430 22370
rect 8482 22318 8494 22370
rect 7758 22306 7810 22318
rect 9326 22306 9378 22318
rect 9774 22370 9826 22382
rect 11566 22370 11618 22382
rect 9986 22318 9998 22370
rect 10050 22318 10062 22370
rect 9774 22306 9826 22318
rect 11566 22306 11618 22318
rect 11678 22370 11730 22382
rect 11678 22306 11730 22318
rect 11902 22370 11954 22382
rect 11902 22306 11954 22318
rect 12014 22370 12066 22382
rect 16718 22370 16770 22382
rect 14578 22318 14590 22370
rect 14642 22318 14654 22370
rect 12014 22306 12066 22318
rect 16718 22306 16770 22318
rect 18174 22370 18226 22382
rect 18174 22306 18226 22318
rect 20078 22370 20130 22382
rect 27246 22370 27298 22382
rect 42030 22370 42082 22382
rect 21746 22318 21758 22370
rect 21810 22318 21822 22370
rect 22194 22318 22206 22370
rect 22258 22318 22270 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 39442 22318 39454 22370
rect 39506 22318 39518 22370
rect 46162 22318 46174 22370
rect 46226 22318 46238 22370
rect 20078 22306 20130 22318
rect 27246 22306 27298 22318
rect 42030 22306 42082 22318
rect 10670 22258 10722 22270
rect 38334 22258 38386 22270
rect 17602 22206 17614 22258
rect 17666 22206 17678 22258
rect 22866 22206 22878 22258
rect 22930 22206 22942 22258
rect 10670 22194 10722 22206
rect 38334 22194 38386 22206
rect 38558 22258 38610 22270
rect 46846 22258 46898 22270
rect 39778 22206 39790 22258
rect 39842 22206 39854 22258
rect 38558 22194 38610 22206
rect 46846 22194 46898 22206
rect 47070 22258 47122 22270
rect 47070 22194 47122 22206
rect 7534 22146 7586 22158
rect 16830 22146 16882 22158
rect 16034 22094 16046 22146
rect 16098 22094 16110 22146
rect 7534 22082 7586 22094
rect 16830 22082 16882 22094
rect 17054 22146 17106 22158
rect 17054 22082 17106 22094
rect 17278 22146 17330 22158
rect 18846 22146 18898 22158
rect 18498 22094 18510 22146
rect 18562 22094 18574 22146
rect 17278 22082 17330 22094
rect 18846 22082 18898 22094
rect 27582 22146 27634 22158
rect 27582 22082 27634 22094
rect 40462 22146 40514 22158
rect 40462 22082 40514 22094
rect 46958 22146 47010 22158
rect 46958 22082 47010 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 10222 21810 10274 21822
rect 10222 21746 10274 21758
rect 10782 21810 10834 21822
rect 10782 21746 10834 21758
rect 10894 21810 10946 21822
rect 10894 21746 10946 21758
rect 11454 21810 11506 21822
rect 11454 21746 11506 21758
rect 13582 21810 13634 21822
rect 14926 21810 14978 21822
rect 13906 21758 13918 21810
rect 13970 21758 13982 21810
rect 13582 21746 13634 21758
rect 14926 21746 14978 21758
rect 18398 21810 18450 21822
rect 18398 21746 18450 21758
rect 20190 21810 20242 21822
rect 20190 21746 20242 21758
rect 20526 21810 20578 21822
rect 20526 21746 20578 21758
rect 45278 21810 45330 21822
rect 45278 21746 45330 21758
rect 45502 21810 45554 21822
rect 45502 21746 45554 21758
rect 46398 21810 46450 21822
rect 46398 21746 46450 21758
rect 17726 21698 17778 21710
rect 17726 21634 17778 21646
rect 18286 21698 18338 21710
rect 29038 21698 29090 21710
rect 26114 21646 26126 21698
rect 26178 21646 26190 21698
rect 18286 21634 18338 21646
rect 29038 21634 29090 21646
rect 30494 21698 30546 21710
rect 30494 21634 30546 21646
rect 30606 21698 30658 21710
rect 30606 21634 30658 21646
rect 31726 21698 31778 21710
rect 42242 21646 42254 21698
rect 42306 21646 42318 21698
rect 44818 21646 44830 21698
rect 44882 21646 44894 21698
rect 31726 21634 31778 21646
rect 1710 21586 1762 21598
rect 1710 21522 1762 21534
rect 2270 21586 2322 21598
rect 8318 21586 8370 21598
rect 5058 21534 5070 21586
rect 5122 21534 5134 21586
rect 2270 21522 2322 21534
rect 8318 21522 8370 21534
rect 14814 21586 14866 21598
rect 14814 21522 14866 21534
rect 15150 21586 15202 21598
rect 16494 21586 16546 21598
rect 15698 21534 15710 21586
rect 15762 21534 15774 21586
rect 15150 21522 15202 21534
rect 16494 21522 16546 21534
rect 17614 21586 17666 21598
rect 17614 21522 17666 21534
rect 18622 21586 18674 21598
rect 18622 21522 18674 21534
rect 20638 21586 20690 21598
rect 30270 21586 30322 21598
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 27346 21534 27358 21586
rect 27410 21534 27422 21586
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 42690 21534 42702 21586
rect 42754 21534 42766 21586
rect 43474 21534 43486 21586
rect 43538 21534 43550 21586
rect 45826 21534 45838 21586
rect 45890 21534 45902 21586
rect 46946 21534 46958 21586
rect 47010 21534 47022 21586
rect 20638 21522 20690 21534
rect 30270 21522 30322 21534
rect 9662 21474 9714 21486
rect 25790 21474 25842 21486
rect 28366 21474 28418 21486
rect 45390 21474 45442 21486
rect 5730 21422 5742 21474
rect 5794 21422 5806 21474
rect 7858 21422 7870 21474
rect 7922 21422 7934 21474
rect 15810 21422 15822 21474
rect 15874 21422 15886 21474
rect 27010 21422 27022 21474
rect 27074 21422 27086 21474
rect 29922 21422 29934 21474
rect 29986 21422 29998 21474
rect 48066 21422 48078 21474
rect 48130 21422 48142 21474
rect 9662 21410 9714 21422
rect 25790 21410 25842 21422
rect 28366 21410 28418 21422
rect 45390 21410 45442 21422
rect 10670 21362 10722 21374
rect 10670 21298 10722 21310
rect 17726 21362 17778 21374
rect 17726 21298 17778 21310
rect 20526 21362 20578 21374
rect 20526 21298 20578 21310
rect 31614 21362 31666 21374
rect 31614 21298 31666 21310
rect 31950 21362 32002 21374
rect 31950 21298 32002 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 37774 21026 37826 21038
rect 41470 21026 41522 21038
rect 17378 20974 17390 21026
rect 17442 20974 17454 21026
rect 27010 20974 27022 21026
rect 27074 20974 27086 21026
rect 29586 20974 29598 21026
rect 29650 20974 29662 21026
rect 31266 20974 31278 21026
rect 31330 20974 31342 21026
rect 37986 20974 37998 21026
rect 38050 21023 38062 21026
rect 38546 21023 38558 21026
rect 38050 20977 38558 21023
rect 38050 20974 38062 20977
rect 38546 20974 38558 20977
rect 38610 20974 38622 21026
rect 37774 20962 37826 20974
rect 41470 20962 41522 20974
rect 1822 20914 1874 20926
rect 19630 20914 19682 20926
rect 17154 20862 17166 20914
rect 17218 20862 17230 20914
rect 18946 20862 18958 20914
rect 19010 20862 19022 20914
rect 1822 20850 1874 20862
rect 19630 20850 19682 20862
rect 25230 20914 25282 20926
rect 28590 20914 28642 20926
rect 39118 20914 39170 20926
rect 27346 20862 27358 20914
rect 27410 20862 27422 20914
rect 30034 20862 30046 20914
rect 30098 20862 30110 20914
rect 32610 20862 32622 20914
rect 32674 20862 32686 20914
rect 45602 20862 45614 20914
rect 45666 20862 45678 20914
rect 25230 20850 25282 20862
rect 28590 20850 28642 20862
rect 39118 20850 39170 20862
rect 15486 20802 15538 20814
rect 5954 20750 5966 20802
rect 6018 20750 6030 20802
rect 10098 20750 10110 20802
rect 10162 20750 10174 20802
rect 15486 20738 15538 20750
rect 15710 20802 15762 20814
rect 20302 20802 20354 20814
rect 16034 20750 16046 20802
rect 16098 20750 16110 20802
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 19282 20750 19294 20802
rect 19346 20750 19358 20802
rect 15710 20738 15762 20750
rect 20302 20738 20354 20750
rect 25902 20802 25954 20814
rect 25902 20738 25954 20750
rect 26126 20802 26178 20814
rect 46734 20802 46786 20814
rect 27234 20750 27246 20802
rect 27298 20750 27310 20802
rect 30146 20750 30158 20802
rect 30210 20750 30222 20802
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 32946 20750 32958 20802
rect 33010 20750 33022 20802
rect 45378 20750 45390 20802
rect 45442 20750 45454 20802
rect 26126 20738 26178 20750
rect 46734 20738 46786 20750
rect 5742 20690 5794 20702
rect 5742 20626 5794 20638
rect 10558 20690 10610 20702
rect 10558 20626 10610 20638
rect 15598 20690 15650 20702
rect 15598 20626 15650 20638
rect 19966 20690 20018 20702
rect 19966 20626 20018 20638
rect 28030 20690 28082 20702
rect 28030 20626 28082 20638
rect 28142 20690 28194 20702
rect 28142 20626 28194 20638
rect 37662 20690 37714 20702
rect 44830 20690 44882 20702
rect 41682 20638 41694 20690
rect 41746 20638 41758 20690
rect 42130 20638 42142 20690
rect 42194 20638 42206 20690
rect 37662 20626 37714 20638
rect 44830 20626 44882 20638
rect 20190 20578 20242 20590
rect 20190 20514 20242 20526
rect 22542 20578 22594 20590
rect 22542 20514 22594 20526
rect 25678 20578 25730 20590
rect 25678 20514 25730 20526
rect 26014 20578 26066 20590
rect 26014 20514 26066 20526
rect 27806 20578 27858 20590
rect 27806 20514 27858 20526
rect 36094 20578 36146 20590
rect 36094 20514 36146 20526
rect 38222 20578 38274 20590
rect 38222 20514 38274 20526
rect 38670 20578 38722 20590
rect 38670 20514 38722 20526
rect 41134 20578 41186 20590
rect 41134 20514 41186 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 17726 20242 17778 20254
rect 17726 20178 17778 20190
rect 21198 20242 21250 20254
rect 21198 20178 21250 20190
rect 22094 20242 22146 20254
rect 22094 20178 22146 20190
rect 30158 20242 30210 20254
rect 30158 20178 30210 20190
rect 31278 20242 31330 20254
rect 31278 20178 31330 20190
rect 32286 20242 32338 20254
rect 32286 20178 32338 20190
rect 33406 20242 33458 20254
rect 33406 20178 33458 20190
rect 37886 20242 37938 20254
rect 41022 20242 41074 20254
rect 37886 20178 37938 20190
rect 38670 20186 38722 20198
rect 9886 20130 9938 20142
rect 9886 20066 9938 20078
rect 12798 20130 12850 20142
rect 12798 20066 12850 20078
rect 14590 20130 14642 20142
rect 14590 20066 14642 20078
rect 17950 20130 18002 20142
rect 22318 20130 22370 20142
rect 21522 20078 21534 20130
rect 21586 20078 21598 20130
rect 17950 20066 18002 20078
rect 22318 20066 22370 20078
rect 24222 20130 24274 20142
rect 24222 20066 24274 20078
rect 26014 20130 26066 20142
rect 28590 20130 28642 20142
rect 27234 20078 27246 20130
rect 27298 20078 27310 20130
rect 26014 20066 26066 20078
rect 28590 20066 28642 20078
rect 29934 20130 29986 20142
rect 29934 20066 29986 20078
rect 31502 20130 31554 20142
rect 31502 20066 31554 20078
rect 32062 20130 32114 20142
rect 32062 20066 32114 20078
rect 32398 20130 32450 20142
rect 36430 20130 36482 20142
rect 35074 20078 35086 20130
rect 35138 20078 35150 20130
rect 32398 20066 32450 20078
rect 36430 20066 36482 20078
rect 38110 20130 38162 20142
rect 41022 20178 41074 20190
rect 43262 20242 43314 20254
rect 43262 20178 43314 20190
rect 45390 20242 45442 20254
rect 45390 20178 45442 20190
rect 38670 20122 38722 20134
rect 45166 20130 45218 20142
rect 39778 20078 39790 20130
rect 39842 20078 39854 20130
rect 38110 20066 38162 20078
rect 45166 20066 45218 20078
rect 45502 20130 45554 20142
rect 45502 20066 45554 20078
rect 47406 20130 47458 20142
rect 47406 20066 47458 20078
rect 11902 20018 11954 20030
rect 10546 19966 10558 20018
rect 10610 19966 10622 20018
rect 11902 19954 11954 19966
rect 17278 20018 17330 20030
rect 20414 20018 20466 20030
rect 23214 20018 23266 20030
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 21858 19966 21870 20018
rect 21922 19966 21934 20018
rect 22754 19966 22766 20018
rect 22818 19966 22830 20018
rect 17278 19954 17330 19966
rect 20414 19954 20466 19966
rect 23214 19954 23266 19966
rect 30270 20018 30322 20030
rect 30270 19954 30322 19966
rect 30606 20018 30658 20030
rect 30606 19954 30658 19966
rect 31390 20018 31442 20030
rect 31390 19954 31442 19966
rect 31950 20018 32002 20030
rect 36206 20018 36258 20030
rect 34290 19966 34302 20018
rect 34354 19966 34366 20018
rect 35186 19966 35198 20018
rect 35250 19966 35262 20018
rect 31950 19954 32002 19966
rect 36206 19954 36258 19966
rect 36878 20018 36930 20030
rect 36878 19954 36930 19966
rect 37102 20018 37154 20030
rect 37102 19954 37154 19966
rect 38222 20018 38274 20030
rect 38222 19954 38274 19966
rect 38782 20018 38834 20030
rect 44382 20018 44434 20030
rect 39330 19966 39342 20018
rect 39394 19966 39406 20018
rect 40226 19966 40238 20018
rect 40290 19966 40302 20018
rect 42242 19966 42254 20018
rect 42306 19966 42318 20018
rect 38782 19954 38834 19966
rect 44382 19954 44434 19966
rect 44606 20018 44658 20030
rect 44606 19954 44658 19966
rect 45054 20018 45106 20030
rect 47618 19966 47630 20018
rect 47682 19966 47694 20018
rect 45054 19954 45106 19966
rect 15150 19906 15202 19918
rect 11106 19854 11118 19906
rect 11170 19854 11182 19906
rect 12338 19854 12350 19906
rect 12402 19854 12414 19906
rect 15150 19842 15202 19854
rect 17838 19906 17890 19918
rect 29038 19906 29090 19918
rect 25218 19854 25230 19906
rect 25282 19854 25294 19906
rect 27906 19854 27918 19906
rect 27970 19854 27982 19906
rect 17838 19842 17890 19854
rect 29038 19842 29090 19854
rect 30718 19906 30770 19918
rect 30718 19842 30770 19854
rect 36318 19906 36370 19918
rect 42702 19906 42754 19918
rect 37538 19854 37550 19906
rect 37602 19854 37614 19906
rect 39890 19854 39902 19906
rect 39954 19854 39966 19906
rect 41794 19854 41806 19906
rect 41858 19854 41870 19906
rect 36318 19842 36370 19854
rect 42702 19842 42754 19854
rect 43038 19906 43090 19918
rect 43038 19842 43090 19854
rect 44494 19906 44546 19918
rect 44494 19842 44546 19854
rect 47182 19906 47234 19918
rect 47182 19842 47234 19854
rect 9998 19794 10050 19806
rect 22430 19794 22482 19806
rect 13794 19742 13806 19794
rect 13858 19742 13870 19794
rect 20290 19742 20302 19794
rect 20354 19742 20366 19794
rect 9998 19730 10050 19742
rect 22430 19730 22482 19742
rect 38670 19794 38722 19806
rect 38670 19730 38722 19742
rect 43374 19794 43426 19806
rect 43374 19730 43426 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 14030 19458 14082 19470
rect 14030 19394 14082 19406
rect 22766 19458 22818 19470
rect 22766 19394 22818 19406
rect 37550 19458 37602 19470
rect 41570 19406 41582 19458
rect 41634 19406 41646 19458
rect 37550 19394 37602 19406
rect 15038 19346 15090 19358
rect 15038 19282 15090 19294
rect 21534 19346 21586 19358
rect 21534 19282 21586 19294
rect 23998 19346 24050 19358
rect 23998 19282 24050 19294
rect 25566 19346 25618 19358
rect 25566 19282 25618 19294
rect 32622 19346 32674 19358
rect 32622 19282 32674 19294
rect 33742 19346 33794 19358
rect 33742 19282 33794 19294
rect 34190 19346 34242 19358
rect 34190 19282 34242 19294
rect 34750 19346 34802 19358
rect 34750 19282 34802 19294
rect 35310 19346 35362 19358
rect 37214 19346 37266 19358
rect 45838 19346 45890 19358
rect 36194 19294 36206 19346
rect 36258 19294 36270 19346
rect 41010 19294 41022 19346
rect 41074 19294 41086 19346
rect 35310 19282 35362 19294
rect 37214 19282 37266 19294
rect 45838 19282 45890 19294
rect 11230 19234 11282 19246
rect 9762 19182 9774 19234
rect 9826 19182 9838 19234
rect 10322 19182 10334 19234
rect 10386 19182 10398 19234
rect 11230 19170 11282 19182
rect 11790 19234 11842 19246
rect 11790 19170 11842 19182
rect 12014 19234 12066 19246
rect 12014 19170 12066 19182
rect 12462 19234 12514 19246
rect 22318 19234 22370 19246
rect 21970 19182 21982 19234
rect 22034 19182 22046 19234
rect 12462 19170 12514 19182
rect 22318 19170 22370 19182
rect 22542 19234 22594 19246
rect 25454 19234 25506 19246
rect 23538 19182 23550 19234
rect 23602 19182 23614 19234
rect 24882 19182 24894 19234
rect 24946 19182 24958 19234
rect 22542 19170 22594 19182
rect 25454 19170 25506 19182
rect 26126 19234 26178 19246
rect 26126 19170 26178 19182
rect 33406 19234 33458 19246
rect 33406 19170 33458 19182
rect 33630 19234 33682 19246
rect 33630 19170 33682 19182
rect 33966 19234 34018 19246
rect 33966 19170 34018 19182
rect 34526 19234 34578 19246
rect 36990 19234 37042 19246
rect 35970 19182 35982 19234
rect 36034 19182 36046 19234
rect 34526 19170 34578 19182
rect 36990 19170 37042 19182
rect 38334 19234 38386 19246
rect 44942 19234 44994 19246
rect 38658 19182 38670 19234
rect 38722 19182 38734 19234
rect 38994 19182 39006 19234
rect 39058 19182 39070 19234
rect 39666 19182 39678 19234
rect 39730 19182 39742 19234
rect 40226 19182 40238 19234
rect 40290 19182 40302 19234
rect 40898 19182 40910 19234
rect 40962 19182 40974 19234
rect 45378 19182 45390 19234
rect 45442 19182 45454 19234
rect 47170 19182 47182 19234
rect 47234 19182 47246 19234
rect 38334 19170 38386 19182
rect 44942 19170 44994 19182
rect 11342 19122 11394 19134
rect 9874 19070 9886 19122
rect 9938 19070 9950 19122
rect 11342 19058 11394 19070
rect 13470 19122 13522 19134
rect 13470 19058 13522 19070
rect 13918 19122 13970 19134
rect 13918 19058 13970 19070
rect 21758 19122 21810 19134
rect 39778 19070 39790 19122
rect 39842 19070 39854 19122
rect 48066 19070 48078 19122
rect 48130 19070 48142 19122
rect 21758 19058 21810 19070
rect 9214 19010 9266 19022
rect 11006 19010 11058 19022
rect 10434 18958 10446 19010
rect 10498 18958 10510 19010
rect 9214 18946 9266 18958
rect 11006 18946 11058 18958
rect 11454 19010 11506 19022
rect 11454 18946 11506 18958
rect 12238 19010 12290 19022
rect 12238 18946 12290 18958
rect 12574 19010 12626 19022
rect 12574 18946 12626 18958
rect 12910 19010 12962 19022
rect 12910 18946 12962 18958
rect 13694 19010 13746 19022
rect 13694 18946 13746 18958
rect 22206 19010 22258 19022
rect 38110 19010 38162 19022
rect 23090 18958 23102 19010
rect 23154 18958 23166 19010
rect 22206 18946 22258 18958
rect 38110 18946 38162 18958
rect 38222 19010 38274 19022
rect 38222 18946 38274 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 9774 18674 9826 18686
rect 9774 18610 9826 18622
rect 11230 18674 11282 18686
rect 31950 18674 32002 18686
rect 34862 18674 34914 18686
rect 36318 18674 36370 18686
rect 15250 18622 15262 18674
rect 15314 18622 15326 18674
rect 33394 18622 33406 18674
rect 33458 18622 33470 18674
rect 36082 18622 36094 18674
rect 36146 18622 36158 18674
rect 11230 18610 11282 18622
rect 31950 18610 32002 18622
rect 34862 18610 34914 18622
rect 36318 18610 36370 18622
rect 38222 18674 38274 18686
rect 38222 18610 38274 18622
rect 38334 18618 38386 18630
rect 10670 18562 10722 18574
rect 10670 18498 10722 18510
rect 11006 18562 11058 18574
rect 20974 18562 21026 18574
rect 31726 18562 31778 18574
rect 12226 18510 12238 18562
rect 12290 18510 12302 18562
rect 14578 18510 14590 18562
rect 14642 18510 14654 18562
rect 29026 18510 29038 18562
rect 29090 18510 29102 18562
rect 11006 18498 11058 18510
rect 20974 18498 21026 18510
rect 31726 18498 31778 18510
rect 36542 18562 36594 18574
rect 36542 18498 36594 18510
rect 36654 18562 36706 18574
rect 38334 18554 38386 18566
rect 38782 18562 38834 18574
rect 36654 18498 36706 18510
rect 38782 18498 38834 18510
rect 40350 18562 40402 18574
rect 40350 18498 40402 18510
rect 10334 18450 10386 18462
rect 10098 18398 10110 18450
rect 10162 18398 10174 18450
rect 10334 18386 10386 18398
rect 10558 18450 10610 18462
rect 14926 18450 14978 18462
rect 32286 18450 32338 18462
rect 12450 18398 12462 18450
rect 12514 18398 12526 18450
rect 13234 18398 13246 18450
rect 13298 18398 13310 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 20290 18398 20302 18450
rect 20354 18398 20366 18450
rect 21746 18398 21758 18450
rect 21810 18398 21822 18450
rect 22530 18398 22542 18450
rect 22594 18398 22606 18450
rect 28802 18398 28814 18450
rect 28866 18398 28878 18450
rect 10558 18386 10610 18398
rect 14926 18386 14978 18398
rect 32286 18386 32338 18398
rect 35534 18450 35586 18462
rect 35534 18386 35586 18398
rect 35758 18450 35810 18462
rect 38670 18450 38722 18462
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 35758 18386 35810 18398
rect 38670 18386 38722 18398
rect 39006 18450 39058 18462
rect 39006 18386 39058 18398
rect 39454 18450 39506 18462
rect 39890 18398 39902 18450
rect 39954 18398 39966 18450
rect 39454 18386 39506 18398
rect 15710 18338 15762 18350
rect 19182 18338 19234 18350
rect 21422 18338 21474 18350
rect 25342 18338 25394 18350
rect 18722 18286 18734 18338
rect 18786 18286 18798 18338
rect 20066 18286 20078 18338
rect 20130 18286 20142 18338
rect 24658 18286 24670 18338
rect 24722 18286 24734 18338
rect 15710 18274 15762 18286
rect 19182 18274 19234 18286
rect 21422 18274 21474 18286
rect 25342 18274 25394 18286
rect 29934 18338 29986 18350
rect 29934 18274 29986 18286
rect 31166 18338 31218 18350
rect 33966 18338 34018 18350
rect 31826 18286 31838 18338
rect 31890 18286 31902 18338
rect 31166 18274 31218 18286
rect 33966 18274 34018 18286
rect 34414 18338 34466 18350
rect 34414 18274 34466 18286
rect 37214 18338 37266 18350
rect 37214 18274 37266 18286
rect 11342 18226 11394 18238
rect 11342 18162 11394 18174
rect 15934 18226 15986 18238
rect 15934 18162 15986 18174
rect 16270 18226 16322 18238
rect 16270 18162 16322 18174
rect 33742 18226 33794 18238
rect 38222 18226 38274 18238
rect 34402 18174 34414 18226
rect 34466 18223 34478 18226
rect 34850 18223 34862 18226
rect 34466 18177 34862 18223
rect 34466 18174 34478 18177
rect 34850 18174 34862 18177
rect 34914 18174 34926 18226
rect 33742 18162 33794 18174
rect 38222 18162 38274 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 18734 17890 18786 17902
rect 18734 17826 18786 17838
rect 36094 17890 36146 17902
rect 36094 17826 36146 17838
rect 11118 17778 11170 17790
rect 11118 17714 11170 17726
rect 14590 17778 14642 17790
rect 29374 17778 29426 17790
rect 26226 17726 26238 17778
rect 26290 17726 26302 17778
rect 28354 17726 28366 17778
rect 28418 17726 28430 17778
rect 14590 17714 14642 17726
rect 29374 17714 29426 17726
rect 31278 17778 31330 17790
rect 31278 17714 31330 17726
rect 31726 17778 31778 17790
rect 31726 17714 31778 17726
rect 32398 17778 32450 17790
rect 32398 17714 32450 17726
rect 34526 17778 34578 17790
rect 34526 17714 34578 17726
rect 35422 17778 35474 17790
rect 35422 17714 35474 17726
rect 37214 17778 37266 17790
rect 37214 17714 37266 17726
rect 39678 17778 39730 17790
rect 39678 17714 39730 17726
rect 40126 17778 40178 17790
rect 42130 17726 42142 17778
rect 42194 17726 42206 17778
rect 40126 17714 40178 17726
rect 18510 17666 18562 17678
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 14354 17614 14366 17666
rect 14418 17614 14430 17666
rect 15810 17614 15822 17666
rect 15874 17614 15886 17666
rect 16706 17614 16718 17666
rect 16770 17614 16782 17666
rect 18510 17602 18562 17614
rect 20302 17666 20354 17678
rect 20302 17602 20354 17614
rect 20526 17666 20578 17678
rect 20526 17602 20578 17614
rect 25118 17666 25170 17678
rect 30270 17666 30322 17678
rect 25554 17614 25566 17666
rect 25618 17614 25630 17666
rect 25118 17602 25170 17614
rect 30270 17602 30322 17614
rect 34862 17666 34914 17678
rect 34862 17602 34914 17614
rect 39006 17666 39058 17678
rect 39006 17602 39058 17614
rect 39342 17666 39394 17678
rect 42018 17614 42030 17666
rect 42082 17614 42094 17666
rect 39342 17602 39394 17614
rect 17390 17554 17442 17566
rect 19966 17554 20018 17566
rect 14578 17502 14590 17554
rect 14642 17502 14654 17554
rect 15586 17502 15598 17554
rect 15650 17502 15662 17554
rect 19058 17502 19070 17554
rect 19122 17502 19134 17554
rect 17390 17490 17442 17502
rect 19966 17490 20018 17502
rect 36206 17554 36258 17566
rect 36206 17490 36258 17502
rect 37886 17554 37938 17566
rect 37886 17490 37938 17502
rect 39118 17554 39170 17566
rect 39118 17490 39170 17502
rect 42702 17554 42754 17566
rect 42702 17490 42754 17502
rect 43038 17554 43090 17566
rect 43038 17490 43090 17502
rect 43262 17554 43314 17566
rect 43262 17490 43314 17502
rect 20414 17442 20466 17454
rect 20414 17378 20466 17390
rect 29934 17442 29986 17454
rect 29934 17378 29986 17390
rect 30382 17442 30434 17454
rect 30382 17378 30434 17390
rect 30494 17442 30546 17454
rect 30494 17378 30546 17390
rect 30718 17442 30770 17454
rect 30718 17378 30770 17390
rect 31166 17442 31218 17454
rect 31166 17378 31218 17390
rect 36094 17442 36146 17454
rect 36094 17378 36146 17390
rect 38334 17442 38386 17454
rect 38334 17378 38386 17390
rect 43150 17442 43202 17454
rect 43150 17378 43202 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 13918 17106 13970 17118
rect 13918 17042 13970 17054
rect 14814 17106 14866 17118
rect 14814 17042 14866 17054
rect 16382 17106 16434 17118
rect 16382 17042 16434 17054
rect 16606 17106 16658 17118
rect 16606 17042 16658 17054
rect 21646 17106 21698 17118
rect 21646 17042 21698 17054
rect 28590 17106 28642 17118
rect 28590 17042 28642 17054
rect 32286 17106 32338 17118
rect 32286 17042 32338 17054
rect 33630 17106 33682 17118
rect 33630 17042 33682 17054
rect 34190 17106 34242 17118
rect 34190 17042 34242 17054
rect 36542 17106 36594 17118
rect 36542 17042 36594 17054
rect 38782 17106 38834 17118
rect 38782 17042 38834 17054
rect 11118 16994 11170 17006
rect 11118 16930 11170 16942
rect 11230 16994 11282 17006
rect 11230 16930 11282 16942
rect 14254 16994 14306 17006
rect 14254 16930 14306 16942
rect 14702 16994 14754 17006
rect 14702 16930 14754 16942
rect 15038 16994 15090 17006
rect 15038 16930 15090 16942
rect 21422 16994 21474 17006
rect 21422 16930 21474 16942
rect 22206 16994 22258 17006
rect 45726 16994 45778 17006
rect 33282 16942 33294 16994
rect 33346 16942 33358 16994
rect 22206 16930 22258 16942
rect 45726 16930 45778 16942
rect 11454 16882 11506 16894
rect 11454 16818 11506 16830
rect 14142 16882 14194 16894
rect 14142 16818 14194 16830
rect 14478 16882 14530 16894
rect 14478 16818 14530 16830
rect 15262 16882 15314 16894
rect 15262 16818 15314 16830
rect 15486 16882 15538 16894
rect 16158 16882 16210 16894
rect 21086 16882 21138 16894
rect 31838 16882 31890 16894
rect 15810 16830 15822 16882
rect 15874 16830 15886 16882
rect 18722 16830 18734 16882
rect 18786 16830 18798 16882
rect 29922 16830 29934 16882
rect 29986 16830 29998 16882
rect 30594 16830 30606 16882
rect 30658 16830 30670 16882
rect 15486 16818 15538 16830
rect 16158 16818 16210 16830
rect 21086 16818 21138 16830
rect 31838 16818 31890 16830
rect 32062 16882 32114 16894
rect 32062 16818 32114 16830
rect 32398 16882 32450 16894
rect 47742 16882 47794 16894
rect 41570 16830 41582 16882
rect 41634 16830 41646 16882
rect 43250 16830 43262 16882
rect 43314 16830 43326 16882
rect 45042 16830 45054 16882
rect 45106 16830 45118 16882
rect 47058 16830 47070 16882
rect 47122 16830 47134 16882
rect 32398 16818 32450 16830
rect 47742 16818 47794 16830
rect 16270 16770 16322 16782
rect 19182 16770 19234 16782
rect 18834 16718 18846 16770
rect 18898 16718 18910 16770
rect 16270 16706 16322 16718
rect 19182 16706 19234 16718
rect 29822 16770 29874 16782
rect 29822 16706 29874 16718
rect 31278 16770 31330 16782
rect 42142 16770 42194 16782
rect 41682 16718 41694 16770
rect 41746 16718 41758 16770
rect 43026 16718 43038 16770
rect 43090 16718 43102 16770
rect 44930 16718 44942 16770
rect 44994 16718 45006 16770
rect 31278 16706 31330 16718
rect 42142 16706 42194 16718
rect 21310 16658 21362 16670
rect 30258 16606 30270 16658
rect 30322 16606 30334 16658
rect 43586 16606 43598 16658
rect 43650 16606 43662 16658
rect 21310 16594 21362 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 12350 16322 12402 16334
rect 43262 16322 43314 16334
rect 24546 16270 24558 16322
rect 24610 16319 24622 16322
rect 24882 16319 24894 16322
rect 24610 16273 24894 16319
rect 24610 16270 24622 16273
rect 24882 16270 24894 16273
rect 24946 16270 24958 16322
rect 32386 16270 32398 16322
rect 32450 16319 32462 16322
rect 32946 16319 32958 16322
rect 32450 16273 32958 16319
rect 32450 16270 32462 16273
rect 32946 16270 32958 16273
rect 33010 16270 33022 16322
rect 12350 16258 12402 16270
rect 43262 16258 43314 16270
rect 15262 16210 15314 16222
rect 20862 16210 20914 16222
rect 23102 16210 23154 16222
rect 14690 16158 14702 16210
rect 14754 16158 14766 16210
rect 20178 16158 20190 16210
rect 20242 16158 20254 16210
rect 22082 16158 22094 16210
rect 22146 16158 22158 16210
rect 15262 16146 15314 16158
rect 20862 16146 20914 16158
rect 23102 16146 23154 16158
rect 24446 16210 24498 16222
rect 24446 16146 24498 16158
rect 24894 16210 24946 16222
rect 29374 16210 29426 16222
rect 32510 16210 32562 16222
rect 25890 16158 25902 16210
rect 25954 16158 25966 16210
rect 28018 16158 28030 16210
rect 28082 16158 28094 16210
rect 31266 16158 31278 16210
rect 31330 16158 31342 16210
rect 24894 16146 24946 16158
rect 29374 16146 29426 16158
rect 32510 16146 32562 16158
rect 36206 16210 36258 16222
rect 36206 16146 36258 16158
rect 37102 16210 37154 16222
rect 45614 16210 45666 16222
rect 42242 16158 42254 16210
rect 42306 16158 42318 16210
rect 43026 16158 43038 16210
rect 43090 16158 43102 16210
rect 37102 16146 37154 16158
rect 45614 16146 45666 16158
rect 47070 16210 47122 16222
rect 47070 16146 47122 16158
rect 10446 16098 10498 16110
rect 10446 16034 10498 16046
rect 10670 16098 10722 16110
rect 10670 16034 10722 16046
rect 11454 16098 11506 16110
rect 11454 16034 11506 16046
rect 11566 16098 11618 16110
rect 11566 16034 11618 16046
rect 11902 16098 11954 16110
rect 11902 16034 11954 16046
rect 12238 16098 12290 16110
rect 29710 16098 29762 16110
rect 14354 16046 14366 16098
rect 14418 16046 14430 16098
rect 19954 16046 19966 16098
rect 20018 16046 20030 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 21970 16046 21982 16098
rect 22034 16046 22046 16098
rect 25106 16046 25118 16098
rect 25170 16046 25182 16098
rect 12238 16034 12290 16046
rect 29710 16034 29762 16046
rect 29822 16098 29874 16110
rect 29822 16034 29874 16046
rect 29934 16098 29986 16110
rect 29934 16034 29986 16046
rect 30382 16098 30434 16110
rect 32846 16098 32898 16110
rect 31154 16046 31166 16098
rect 31218 16046 31230 16098
rect 32050 16046 32062 16098
rect 32114 16046 32126 16098
rect 42914 16046 42926 16098
rect 42978 16046 42990 16098
rect 44818 16046 44830 16098
rect 44882 16046 44894 16098
rect 47618 16046 47630 16098
rect 47682 16046 47694 16098
rect 30382 16034 30434 16046
rect 32846 16034 32898 16046
rect 19294 15986 19346 15998
rect 41918 15986 41970 15998
rect 22642 15934 22654 15986
rect 22706 15934 22718 15986
rect 30706 15934 30718 15986
rect 30770 15934 30782 15986
rect 19294 15922 19346 15934
rect 41918 15922 41970 15934
rect 42142 15986 42194 15998
rect 45166 15986 45218 15998
rect 42354 15934 42366 15986
rect 42418 15983 42430 15986
rect 42802 15983 42814 15986
rect 42418 15937 42814 15983
rect 42418 15934 42430 15937
rect 42802 15934 42814 15937
rect 42866 15934 42878 15986
rect 42142 15922 42194 15934
rect 45166 15922 45218 15934
rect 45502 15986 45554 15998
rect 45502 15922 45554 15934
rect 47406 15986 47458 15998
rect 47406 15922 47458 15934
rect 11790 15874 11842 15886
rect 10994 15822 11006 15874
rect 11058 15822 11070 15874
rect 11790 15810 11842 15822
rect 12350 15874 12402 15886
rect 12350 15810 12402 15822
rect 23438 15874 23490 15886
rect 45054 15874 45106 15886
rect 23762 15822 23774 15874
rect 23826 15822 23838 15874
rect 23438 15810 23490 15822
rect 45054 15810 45106 15822
rect 45726 15874 45778 15886
rect 45726 15810 45778 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 12126 15538 12178 15550
rect 12126 15474 12178 15486
rect 12350 15538 12402 15550
rect 12350 15474 12402 15486
rect 12574 15538 12626 15550
rect 12574 15474 12626 15486
rect 13134 15538 13186 15550
rect 24334 15538 24386 15550
rect 21522 15486 21534 15538
rect 21586 15486 21598 15538
rect 13134 15474 13186 15486
rect 24334 15474 24386 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 25790 15538 25842 15550
rect 25790 15474 25842 15486
rect 30606 15538 30658 15550
rect 30606 15474 30658 15486
rect 37550 15538 37602 15550
rect 37550 15474 37602 15486
rect 11454 15426 11506 15438
rect 11454 15362 11506 15374
rect 11566 15426 11618 15438
rect 11566 15362 11618 15374
rect 11678 15426 11730 15438
rect 11678 15362 11730 15374
rect 13022 15426 13074 15438
rect 13022 15362 13074 15374
rect 16270 15426 16322 15438
rect 16270 15362 16322 15374
rect 18398 15426 18450 15438
rect 18398 15362 18450 15374
rect 22878 15426 22930 15438
rect 22878 15362 22930 15374
rect 24446 15426 24498 15438
rect 24446 15362 24498 15374
rect 35310 15426 35362 15438
rect 35310 15362 35362 15374
rect 35758 15426 35810 15438
rect 35758 15362 35810 15374
rect 35982 15426 36034 15438
rect 35982 15362 36034 15374
rect 36542 15426 36594 15438
rect 36542 15362 36594 15374
rect 36878 15426 36930 15438
rect 40350 15426 40402 15438
rect 38434 15374 38446 15426
rect 38498 15374 38510 15426
rect 40114 15374 40126 15426
rect 40178 15374 40190 15426
rect 36878 15362 36930 15374
rect 40350 15362 40402 15374
rect 13358 15314 13410 15326
rect 21198 15314 21250 15326
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 13358 15250 13410 15262
rect 21198 15250 21250 15262
rect 22766 15314 22818 15326
rect 22766 15250 22818 15262
rect 24110 15314 24162 15326
rect 31838 15314 31890 15326
rect 31154 15262 31166 15314
rect 31218 15262 31230 15314
rect 24110 15250 24162 15262
rect 31838 15250 31890 15262
rect 36094 15314 36146 15326
rect 36094 15250 36146 15262
rect 37438 15314 37490 15326
rect 37438 15250 37490 15262
rect 37774 15314 37826 15326
rect 37774 15250 37826 15262
rect 12238 15202 12290 15214
rect 26350 15202 26402 15214
rect 17938 15150 17950 15202
rect 18002 15150 18014 15202
rect 12238 15138 12290 15150
rect 26350 15138 26402 15150
rect 35422 15202 35474 15214
rect 35422 15138 35474 15150
rect 38334 15202 38386 15214
rect 38334 15138 38386 15150
rect 22878 15090 22930 15102
rect 35534 15090 35586 15102
rect 10994 15038 11006 15090
rect 11058 15038 11070 15090
rect 31938 15038 31950 15090
rect 32002 15038 32014 15090
rect 22878 15026 22930 15038
rect 35534 15026 35586 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 22430 14754 22482 14766
rect 22430 14690 22482 14702
rect 43710 14754 43762 14766
rect 43710 14690 43762 14702
rect 12350 14642 12402 14654
rect 11554 14590 11566 14642
rect 11618 14590 11630 14642
rect 12350 14578 12402 14590
rect 13470 14642 13522 14654
rect 13470 14578 13522 14590
rect 14702 14642 14754 14654
rect 29710 14642 29762 14654
rect 27458 14590 27470 14642
rect 27522 14590 27534 14642
rect 14702 14578 14754 14590
rect 29710 14578 29762 14590
rect 30158 14642 30210 14654
rect 30158 14578 30210 14590
rect 31166 14642 31218 14654
rect 31166 14578 31218 14590
rect 31614 14642 31666 14654
rect 31614 14578 31666 14590
rect 32062 14642 32114 14654
rect 36542 14642 36594 14654
rect 40462 14642 40514 14654
rect 41806 14642 41858 14654
rect 35858 14590 35870 14642
rect 35922 14590 35934 14642
rect 38322 14590 38334 14642
rect 38386 14590 38398 14642
rect 40002 14590 40014 14642
rect 40066 14590 40078 14642
rect 40898 14590 40910 14642
rect 40962 14590 40974 14642
rect 32062 14578 32114 14590
rect 36542 14578 36594 14590
rect 40462 14578 40514 14590
rect 41806 14578 41858 14590
rect 44830 14642 44882 14654
rect 44830 14578 44882 14590
rect 46734 14642 46786 14654
rect 46734 14578 46786 14590
rect 11118 14530 11170 14542
rect 11118 14466 11170 14478
rect 12574 14530 12626 14542
rect 12574 14466 12626 14478
rect 13022 14530 13074 14542
rect 13022 14466 13074 14478
rect 15710 14530 15762 14542
rect 15710 14466 15762 14478
rect 17614 14530 17666 14542
rect 17614 14466 17666 14478
rect 17838 14530 17890 14542
rect 17838 14466 17890 14478
rect 21534 14530 21586 14542
rect 21534 14466 21586 14478
rect 21758 14530 21810 14542
rect 27918 14530 27970 14542
rect 22866 14478 22878 14530
rect 22930 14478 22942 14530
rect 23314 14478 23326 14530
rect 23378 14478 23390 14530
rect 21758 14466 21810 14478
rect 27918 14466 27970 14478
rect 29150 14530 29202 14542
rect 29150 14466 29202 14478
rect 30494 14530 30546 14542
rect 37214 14530 37266 14542
rect 39118 14530 39170 14542
rect 43822 14530 43874 14542
rect 33282 14478 33294 14530
rect 33346 14478 33358 14530
rect 35410 14478 35422 14530
rect 35474 14478 35486 14530
rect 38210 14478 38222 14530
rect 38274 14478 38286 14530
rect 39778 14478 39790 14530
rect 39842 14478 39854 14530
rect 41122 14478 41134 14530
rect 41186 14478 41198 14530
rect 30494 14466 30546 14478
rect 37214 14466 37266 14478
rect 39118 14466 39170 14478
rect 43822 14466 43874 14478
rect 44046 14530 44098 14542
rect 45054 14530 45106 14542
rect 44258 14478 44270 14530
rect 44322 14478 44334 14530
rect 45378 14478 45390 14530
rect 45442 14478 45454 14530
rect 46946 14478 46958 14530
rect 47010 14478 47022 14530
rect 44046 14466 44098 14478
rect 45054 14466 45106 14478
rect 13582 14418 13634 14430
rect 13582 14354 13634 14366
rect 15374 14418 15426 14430
rect 16494 14418 16546 14430
rect 16034 14366 16046 14418
rect 16098 14366 16110 14418
rect 15374 14354 15426 14366
rect 16494 14354 16546 14366
rect 16606 14418 16658 14430
rect 16606 14354 16658 14366
rect 21422 14418 21474 14430
rect 21422 14354 21474 14366
rect 22318 14418 22370 14430
rect 22318 14354 22370 14366
rect 22654 14418 22706 14430
rect 22654 14354 22706 14366
rect 26574 14418 26626 14430
rect 30606 14418 30658 14430
rect 34974 14418 35026 14430
rect 26898 14366 26910 14418
rect 26962 14366 26974 14418
rect 32722 14366 32734 14418
rect 32786 14366 32798 14418
rect 34402 14366 34414 14418
rect 34466 14366 34478 14418
rect 26574 14354 26626 14366
rect 30606 14354 30658 14366
rect 34974 14354 35026 14366
rect 37102 14418 37154 14430
rect 48066 14366 48078 14418
rect 48130 14366 48142 14418
rect 37102 14354 37154 14366
rect 16270 14306 16322 14318
rect 16270 14242 16322 14254
rect 17390 14306 17442 14318
rect 17390 14242 17442 14254
rect 17726 14306 17778 14318
rect 17726 14242 17778 14254
rect 21198 14306 21250 14318
rect 21198 14242 21250 14254
rect 22094 14306 22146 14318
rect 22094 14242 22146 14254
rect 30830 14306 30882 14318
rect 36878 14306 36930 14318
rect 34290 14254 34302 14306
rect 34354 14254 34366 14306
rect 30830 14242 30882 14254
rect 36878 14242 36930 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 14926 13970 14978 13982
rect 14926 13906 14978 13918
rect 16494 13970 16546 13982
rect 16494 13906 16546 13918
rect 18734 13970 18786 13982
rect 18734 13906 18786 13918
rect 22878 13970 22930 13982
rect 22878 13906 22930 13918
rect 23438 13970 23490 13982
rect 23438 13906 23490 13918
rect 23998 13970 24050 13982
rect 23998 13906 24050 13918
rect 32286 13970 32338 13982
rect 32286 13906 32338 13918
rect 37102 13970 37154 13982
rect 37102 13906 37154 13918
rect 37662 13970 37714 13982
rect 37662 13906 37714 13918
rect 38222 13970 38274 13982
rect 45378 13918 45390 13970
rect 45442 13918 45454 13970
rect 38222 13906 38274 13918
rect 12686 13858 12738 13870
rect 12002 13806 12014 13858
rect 12066 13806 12078 13858
rect 12686 13794 12738 13806
rect 14814 13858 14866 13870
rect 14814 13794 14866 13806
rect 15150 13858 15202 13870
rect 15150 13794 15202 13806
rect 16606 13858 16658 13870
rect 16606 13794 16658 13806
rect 18846 13858 18898 13870
rect 18846 13794 18898 13806
rect 22766 13858 22818 13870
rect 34750 13858 34802 13870
rect 37214 13858 37266 13870
rect 30482 13806 30494 13858
rect 30546 13806 30558 13858
rect 36306 13806 36318 13858
rect 36370 13806 36382 13858
rect 22766 13794 22818 13806
rect 34750 13794 34802 13806
rect 37214 13794 37266 13806
rect 37550 13858 37602 13870
rect 37550 13794 37602 13806
rect 38110 13858 38162 13870
rect 43810 13806 43822 13858
rect 43874 13806 43886 13858
rect 38110 13794 38162 13806
rect 13246 13746 13298 13758
rect 11778 13694 11790 13746
rect 11842 13694 11854 13746
rect 13246 13682 13298 13694
rect 14254 13746 14306 13758
rect 15822 13746 15874 13758
rect 15474 13694 15486 13746
rect 15538 13694 15550 13746
rect 14254 13682 14306 13694
rect 15822 13682 15874 13694
rect 16046 13746 16098 13758
rect 16046 13682 16098 13694
rect 16270 13746 16322 13758
rect 20638 13746 20690 13758
rect 22206 13746 22258 13758
rect 23550 13746 23602 13758
rect 25230 13746 25282 13758
rect 29710 13746 29762 13758
rect 31838 13746 31890 13758
rect 36654 13746 36706 13758
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 21074 13694 21086 13746
rect 21138 13694 21150 13746
rect 22530 13694 22542 13746
rect 22594 13694 22606 13746
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 25666 13694 25678 13746
rect 25730 13694 25742 13746
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 30146 13694 30158 13746
rect 30210 13694 30222 13746
rect 35186 13694 35198 13746
rect 35250 13694 35262 13746
rect 16270 13682 16322 13694
rect 20638 13682 20690 13694
rect 22206 13682 22258 13694
rect 23550 13682 23602 13694
rect 25230 13682 25282 13694
rect 29710 13682 29762 13694
rect 31838 13682 31890 13694
rect 36654 13682 36706 13694
rect 36878 13746 36930 13758
rect 36878 13682 36930 13694
rect 38446 13746 38498 13758
rect 38446 13682 38498 13694
rect 38782 13746 38834 13758
rect 38782 13682 38834 13694
rect 39678 13746 39730 13758
rect 44034 13694 44046 13746
rect 44098 13694 44110 13746
rect 45042 13694 45054 13746
rect 45106 13694 45118 13746
rect 39678 13682 39730 13694
rect 14478 13634 14530 13646
rect 11890 13582 11902 13634
rect 11954 13582 11966 13634
rect 14478 13570 14530 13582
rect 15934 13634 15986 13646
rect 24446 13634 24498 13646
rect 19506 13582 19518 13634
rect 19570 13582 19582 13634
rect 21186 13582 21198 13634
rect 21250 13582 21262 13634
rect 35522 13582 35534 13634
rect 35586 13582 35598 13634
rect 15934 13570 15986 13582
rect 24446 13570 24498 13582
rect 18734 13522 18786 13534
rect 23438 13522 23490 13534
rect 29374 13522 29426 13534
rect 31614 13522 31666 13534
rect 13906 13470 13918 13522
rect 13970 13470 13982 13522
rect 19282 13470 19294 13522
rect 19346 13470 19358 13522
rect 25890 13470 25902 13522
rect 25954 13470 25966 13522
rect 31266 13470 31278 13522
rect 31330 13470 31342 13522
rect 18734 13458 18786 13470
rect 23438 13458 23490 13470
rect 29374 13458 29426 13470
rect 31614 13458 31666 13470
rect 37662 13522 37714 13534
rect 37662 13458 37714 13470
rect 39006 13522 39058 13534
rect 39902 13522 39954 13534
rect 39330 13470 39342 13522
rect 39394 13470 39406 13522
rect 39006 13458 39058 13470
rect 39902 13458 39954 13470
rect 40238 13522 40290 13534
rect 40238 13458 40290 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 18958 13186 19010 13198
rect 18958 13122 19010 13134
rect 15934 13074 15986 13086
rect 20078 13074 20130 13086
rect 26014 13074 26066 13086
rect 37102 13074 37154 13086
rect 14690 13022 14702 13074
rect 14754 13022 14766 13074
rect 17042 13022 17054 13074
rect 17106 13022 17118 13074
rect 24434 13022 24446 13074
rect 24498 13022 24510 13074
rect 25554 13022 25566 13074
rect 25618 13022 25630 13074
rect 29362 13022 29374 13074
rect 29426 13022 29438 13074
rect 30594 13022 30606 13074
rect 30658 13022 30670 13074
rect 32386 13022 32398 13074
rect 32450 13022 32462 13074
rect 15934 13010 15986 13022
rect 20078 13010 20130 13022
rect 26014 13010 26066 13022
rect 37102 13010 37154 13022
rect 41246 13074 41298 13086
rect 41246 13010 41298 13022
rect 43262 13074 43314 13086
rect 43262 13010 43314 13022
rect 12238 12962 12290 12974
rect 12238 12898 12290 12910
rect 13694 12962 13746 12974
rect 19406 12962 19458 12974
rect 34750 12962 34802 12974
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 14802 12910 14814 12962
rect 14866 12910 14878 12962
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 24546 12910 24558 12962
rect 24610 12910 24622 12962
rect 29698 12910 29710 12962
rect 29762 12910 29774 12962
rect 30818 12910 30830 12962
rect 30882 12910 30894 12962
rect 32162 12910 32174 12962
rect 32226 12910 32238 12962
rect 13694 12898 13746 12910
rect 19406 12898 19458 12910
rect 34750 12898 34802 12910
rect 34974 12962 35026 12974
rect 34974 12898 35026 12910
rect 35310 12962 35362 12974
rect 35310 12898 35362 12910
rect 36206 12962 36258 12974
rect 36206 12898 36258 12910
rect 39790 12962 39842 12974
rect 39790 12898 39842 12910
rect 40014 12962 40066 12974
rect 40338 12910 40350 12962
rect 40402 12910 40414 12962
rect 42578 12910 42590 12962
rect 42642 12910 42654 12962
rect 40014 12898 40066 12910
rect 13582 12850 13634 12862
rect 16158 12850 16210 12862
rect 15362 12798 15374 12850
rect 15426 12798 15438 12850
rect 13582 12786 13634 12798
rect 16158 12786 16210 12798
rect 19070 12850 19122 12862
rect 19070 12786 19122 12798
rect 30158 12850 30210 12862
rect 30158 12786 30210 12798
rect 31502 12850 31554 12862
rect 31502 12786 31554 12798
rect 32846 12850 32898 12862
rect 32846 12786 32898 12798
rect 36094 12850 36146 12862
rect 36094 12786 36146 12798
rect 39902 12850 39954 12862
rect 41682 12798 41694 12850
rect 41746 12798 41758 12850
rect 39902 12786 39954 12798
rect 13358 12738 13410 12750
rect 12562 12686 12574 12738
rect 12626 12686 12638 12738
rect 13358 12674 13410 12686
rect 18958 12738 19010 12750
rect 18958 12674 19010 12686
rect 19518 12738 19570 12750
rect 19518 12674 19570 12686
rect 19742 12738 19794 12750
rect 19742 12674 19794 12686
rect 34974 12738 35026 12750
rect 34974 12674 35026 12686
rect 35870 12738 35922 12750
rect 35870 12674 35922 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 14030 12402 14082 12414
rect 14030 12338 14082 12350
rect 15934 12402 15986 12414
rect 15934 12338 15986 12350
rect 16046 12402 16098 12414
rect 16046 12338 16098 12350
rect 16606 12402 16658 12414
rect 16606 12338 16658 12350
rect 20414 12402 20466 12414
rect 20414 12338 20466 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 26350 12402 26402 12414
rect 26350 12338 26402 12350
rect 26910 12402 26962 12414
rect 26910 12338 26962 12350
rect 27582 12402 27634 12414
rect 27582 12338 27634 12350
rect 28142 12402 28194 12414
rect 36542 12402 36594 12414
rect 31266 12350 31278 12402
rect 31330 12350 31342 12402
rect 28142 12338 28194 12350
rect 36542 12338 36594 12350
rect 12350 12290 12402 12302
rect 12350 12226 12402 12238
rect 19070 12290 19122 12302
rect 19070 12226 19122 12238
rect 19406 12290 19458 12302
rect 19406 12226 19458 12238
rect 25342 12290 25394 12302
rect 25342 12226 25394 12238
rect 27806 12290 27858 12302
rect 27806 12226 27858 12238
rect 31838 12290 31890 12302
rect 31838 12226 31890 12238
rect 33182 12290 33234 12302
rect 33182 12226 33234 12238
rect 41022 12290 41074 12302
rect 41022 12226 41074 12238
rect 15150 12178 15202 12190
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 14690 12126 14702 12178
rect 14754 12126 14766 12178
rect 15150 12114 15202 12126
rect 15486 12178 15538 12190
rect 15486 12114 15538 12126
rect 16158 12178 16210 12190
rect 19630 12178 19682 12190
rect 18162 12126 18174 12178
rect 18226 12126 18238 12178
rect 16158 12114 16210 12126
rect 19630 12114 19682 12126
rect 25678 12178 25730 12190
rect 25678 12114 25730 12126
rect 26238 12178 26290 12190
rect 26238 12114 26290 12126
rect 26574 12178 26626 12190
rect 26574 12114 26626 12126
rect 27470 12178 27522 12190
rect 27470 12114 27522 12126
rect 31614 12178 31666 12190
rect 31614 12114 31666 12126
rect 33294 12178 33346 12190
rect 46734 12178 46786 12190
rect 43362 12126 43374 12178
rect 43426 12126 43438 12178
rect 43810 12126 43822 12178
rect 43874 12126 43886 12178
rect 33294 12114 33346 12126
rect 46734 12114 46786 12126
rect 46958 12178 47010 12190
rect 46958 12114 47010 12126
rect 14254 12066 14306 12078
rect 41134 12066 41186 12078
rect 18722 12014 18734 12066
rect 18786 12014 18798 12066
rect 14254 12002 14306 12014
rect 41134 12002 41186 12014
rect 41470 12066 41522 12078
rect 41470 12002 41522 12014
rect 42366 12066 42418 12078
rect 42366 12002 42418 12014
rect 12686 11954 12738 11966
rect 12686 11890 12738 11902
rect 19966 11954 20018 11966
rect 19966 11890 20018 11902
rect 33182 11954 33234 11966
rect 33182 11890 33234 11902
rect 41694 11954 41746 11966
rect 41694 11890 41746 11902
rect 42030 11954 42082 11966
rect 42030 11890 42082 11902
rect 42590 11954 42642 11966
rect 47742 11954 47794 11966
rect 42914 11902 42926 11954
rect 42978 11902 42990 11954
rect 43362 11902 43374 11954
rect 43426 11902 43438 11954
rect 42590 11890 42642 11902
rect 47742 11890 47794 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 15138 11566 15150 11618
rect 15202 11566 15214 11618
rect 25678 11506 25730 11518
rect 29822 11506 29874 11518
rect 15026 11454 15038 11506
rect 15090 11454 15102 11506
rect 24322 11454 24334 11506
rect 24386 11454 24398 11506
rect 27122 11454 27134 11506
rect 27186 11454 27198 11506
rect 25678 11442 25730 11454
rect 29822 11442 29874 11454
rect 11230 11394 11282 11406
rect 11230 11330 11282 11342
rect 11566 11394 11618 11406
rect 18734 11394 18786 11406
rect 11778 11342 11790 11394
rect 11842 11342 11854 11394
rect 12674 11342 12686 11394
rect 12738 11342 12750 11394
rect 14690 11342 14702 11394
rect 14754 11342 14766 11394
rect 11566 11330 11618 11342
rect 18734 11330 18786 11342
rect 19406 11394 19458 11406
rect 24670 11394 24722 11406
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 23202 11342 23214 11394
rect 23266 11342 23278 11394
rect 19406 11330 19458 11342
rect 24670 11330 24722 11342
rect 25902 11394 25954 11406
rect 27582 11394 27634 11406
rect 26898 11342 26910 11394
rect 26962 11342 26974 11394
rect 25902 11330 25954 11342
rect 27582 11330 27634 11342
rect 28142 11394 28194 11406
rect 28142 11330 28194 11342
rect 29150 11394 29202 11406
rect 32846 11394 32898 11406
rect 32274 11342 32286 11394
rect 32338 11342 32350 11394
rect 29150 11330 29202 11342
rect 32846 11330 32898 11342
rect 32958 11394 33010 11406
rect 34190 11394 34242 11406
rect 37774 11394 37826 11406
rect 33730 11342 33742 11394
rect 33794 11342 33806 11394
rect 37314 11342 37326 11394
rect 37378 11342 37390 11394
rect 32958 11330 33010 11342
rect 34190 11330 34242 11342
rect 37774 11330 37826 11342
rect 41918 11394 41970 11406
rect 41918 11330 41970 11342
rect 42254 11394 42306 11406
rect 42254 11330 42306 11342
rect 42478 11394 42530 11406
rect 42478 11330 42530 11342
rect 11342 11282 11394 11294
rect 28030 11282 28082 11294
rect 12226 11230 12238 11282
rect 12290 11230 12302 11282
rect 24994 11230 25006 11282
rect 25058 11230 25070 11282
rect 11342 11218 11394 11230
rect 28030 11218 28082 11230
rect 28590 11282 28642 11294
rect 28590 11218 28642 11230
rect 29262 11282 29314 11294
rect 29262 11218 29314 11230
rect 30270 11282 30322 11294
rect 30270 11218 30322 11230
rect 33294 11282 33346 11294
rect 33294 11218 33346 11230
rect 36206 11282 36258 11294
rect 36206 11218 36258 11230
rect 36318 11282 36370 11294
rect 36318 11218 36370 11230
rect 18846 11170 18898 11182
rect 12786 11118 12798 11170
rect 12850 11118 12862 11170
rect 18846 11106 18898 11118
rect 18958 11170 19010 11182
rect 27806 11170 27858 11182
rect 26226 11118 26238 11170
rect 26290 11118 26302 11170
rect 18958 11106 19010 11118
rect 27806 11106 27858 11118
rect 29486 11170 29538 11182
rect 29486 11106 29538 11118
rect 36542 11170 36594 11182
rect 36542 11106 36594 11118
rect 42142 11170 42194 11182
rect 42142 11106 42194 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 23662 10834 23714 10846
rect 23662 10770 23714 10782
rect 24558 10834 24610 10846
rect 24558 10770 24610 10782
rect 24782 10834 24834 10846
rect 24782 10770 24834 10782
rect 26798 10834 26850 10846
rect 26798 10770 26850 10782
rect 26910 10834 26962 10846
rect 30034 10782 30046 10834
rect 30098 10782 30110 10834
rect 34178 10782 34190 10834
rect 34242 10782 34254 10834
rect 26910 10770 26962 10782
rect 21534 10722 21586 10734
rect 23774 10722 23826 10734
rect 12114 10670 12126 10722
rect 12178 10670 12190 10722
rect 23202 10670 23214 10722
rect 23266 10670 23278 10722
rect 21534 10658 21586 10670
rect 23774 10658 23826 10670
rect 24446 10722 24498 10734
rect 32286 10722 32338 10734
rect 28466 10670 28478 10722
rect 28530 10670 28542 10722
rect 24446 10658 24498 10670
rect 32286 10658 32338 10670
rect 32398 10722 32450 10734
rect 32398 10658 32450 10670
rect 32622 10722 32674 10734
rect 32622 10658 32674 10670
rect 33182 10722 33234 10734
rect 33182 10658 33234 10670
rect 33294 10722 33346 10734
rect 44382 10722 44434 10734
rect 35634 10670 35646 10722
rect 35698 10670 35710 10722
rect 33294 10658 33346 10670
rect 44382 10658 44434 10670
rect 18622 10610 18674 10622
rect 20078 10610 20130 10622
rect 27022 10610 27074 10622
rect 43262 10610 43314 10622
rect 12338 10558 12350 10610
rect 12402 10558 12414 10610
rect 13010 10558 13022 10610
rect 13074 10558 13086 10610
rect 17938 10558 17950 10610
rect 18002 10558 18014 10610
rect 19618 10558 19630 10610
rect 19682 10558 19694 10610
rect 20850 10558 20862 10610
rect 20914 10558 20926 10610
rect 22194 10558 22206 10610
rect 22258 10558 22270 10610
rect 22866 10558 22878 10610
rect 22930 10558 22942 10610
rect 25778 10558 25790 10610
rect 25842 10558 25854 10610
rect 27346 10558 27358 10610
rect 27410 10558 27422 10610
rect 29586 10558 29598 10610
rect 29650 10558 29662 10610
rect 34738 10558 34750 10610
rect 34802 10558 34814 10610
rect 35410 10558 35422 10610
rect 35474 10558 35486 10610
rect 37538 10558 37550 10610
rect 37602 10558 37614 10610
rect 38994 10558 39006 10610
rect 39058 10558 39070 10610
rect 18622 10546 18674 10558
rect 20078 10546 20130 10558
rect 27022 10546 27074 10558
rect 43262 10546 43314 10558
rect 43486 10610 43538 10622
rect 44034 10558 44046 10610
rect 44098 10558 44110 10610
rect 43486 10546 43538 10558
rect 13694 10498 13746 10510
rect 26462 10498 26514 10510
rect 36766 10498 36818 10510
rect 17714 10446 17726 10498
rect 17778 10446 17790 10498
rect 19170 10446 19182 10498
rect 19234 10446 19246 10498
rect 20738 10446 20750 10498
rect 20802 10446 20814 10498
rect 22754 10446 22766 10498
rect 22818 10446 22830 10498
rect 26002 10446 26014 10498
rect 26066 10446 26078 10498
rect 28130 10446 28142 10498
rect 28194 10446 28206 10498
rect 37986 10446 37998 10498
rect 38050 10446 38062 10498
rect 13694 10434 13746 10446
rect 26462 10434 26514 10446
rect 36766 10434 36818 10446
rect 23662 10386 23714 10398
rect 23662 10322 23714 10334
rect 33182 10386 33234 10398
rect 43150 10386 43202 10398
rect 39218 10334 39230 10386
rect 39282 10334 39294 10386
rect 33182 10322 33234 10334
rect 43150 10322 43202 10334
rect 43598 10386 43650 10398
rect 43598 10322 43650 10334
rect 44046 10386 44098 10398
rect 44046 10322 44098 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 21870 10050 21922 10062
rect 21870 9986 21922 9998
rect 22206 10050 22258 10062
rect 22206 9986 22258 9998
rect 26126 10050 26178 10062
rect 26126 9986 26178 9998
rect 26462 10050 26514 10062
rect 26462 9986 26514 9998
rect 16270 9938 16322 9950
rect 16270 9874 16322 9886
rect 17166 9938 17218 9950
rect 17166 9874 17218 9886
rect 18174 9938 18226 9950
rect 18174 9874 18226 9886
rect 25006 9938 25058 9950
rect 25006 9874 25058 9886
rect 25902 9938 25954 9950
rect 31838 9938 31890 9950
rect 31266 9886 31278 9938
rect 31330 9886 31342 9938
rect 25902 9874 25954 9886
rect 31838 9874 31890 9886
rect 34190 9938 34242 9950
rect 39230 9938 39282 9950
rect 46734 9938 46786 9950
rect 34850 9886 34862 9938
rect 34914 9886 34926 9938
rect 44258 9886 44270 9938
rect 44322 9886 44334 9938
rect 34190 9874 34242 9886
rect 39230 9874 39282 9886
rect 46734 9874 46786 9886
rect 16606 9826 16658 9838
rect 14354 9774 14366 9826
rect 14418 9774 14430 9826
rect 15586 9774 15598 9826
rect 15650 9774 15662 9826
rect 16606 9762 16658 9774
rect 18398 9826 18450 9838
rect 18398 9762 18450 9774
rect 19854 9826 19906 9838
rect 19854 9762 19906 9774
rect 20190 9826 20242 9838
rect 20190 9762 20242 9774
rect 26910 9826 26962 9838
rect 37998 9826 38050 9838
rect 29810 9774 29822 9826
rect 29874 9774 29886 9826
rect 34962 9774 34974 9826
rect 35026 9774 35038 9826
rect 26910 9762 26962 9774
rect 37998 9762 38050 9774
rect 38670 9826 38722 9838
rect 42814 9826 42866 9838
rect 40786 9774 40798 9826
rect 40850 9774 40862 9826
rect 42130 9774 42142 9826
rect 42194 9774 42206 9826
rect 43474 9774 43486 9826
rect 43538 9774 43550 9826
rect 46946 9774 46958 9826
rect 47010 9774 47022 9826
rect 38670 9762 38722 9774
rect 42814 9762 42866 9774
rect 14590 9714 14642 9726
rect 19630 9714 19682 9726
rect 15810 9662 15822 9714
rect 15874 9662 15886 9714
rect 18722 9662 18734 9714
rect 18786 9662 18798 9714
rect 14590 9650 14642 9662
rect 19630 9650 19682 9662
rect 21646 9714 21698 9726
rect 21646 9650 21698 9662
rect 27022 9714 27074 9726
rect 27022 9650 27074 9662
rect 27582 9714 27634 9726
rect 34526 9714 34578 9726
rect 30706 9662 30718 9714
rect 30770 9662 30782 9714
rect 27582 9650 27634 9662
rect 34526 9650 34578 9662
rect 37438 9714 37490 9726
rect 37438 9650 37490 9662
rect 38110 9714 38162 9726
rect 38110 9650 38162 9662
rect 38334 9714 38386 9726
rect 39330 9662 39342 9714
rect 39394 9662 39406 9714
rect 48066 9662 48078 9714
rect 48130 9662 48142 9714
rect 38334 9650 38386 9662
rect 20078 9602 20130 9614
rect 15474 9550 15486 9602
rect 15538 9550 15550 9602
rect 20078 9538 20130 9550
rect 27246 9602 27298 9614
rect 31726 9602 31778 9614
rect 29474 9550 29486 9602
rect 29538 9550 29550 9602
rect 40898 9550 40910 9602
rect 40962 9550 40974 9602
rect 27246 9538 27298 9550
rect 31726 9538 31778 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 31278 9266 31330 9278
rect 31278 9202 31330 9214
rect 31390 9266 31442 9278
rect 31390 9202 31442 9214
rect 38670 9266 38722 9278
rect 38670 9202 38722 9214
rect 42926 9266 42978 9278
rect 42926 9202 42978 9214
rect 43934 9266 43986 9278
rect 43934 9202 43986 9214
rect 44158 9266 44210 9278
rect 44158 9202 44210 9214
rect 14366 9154 14418 9166
rect 14366 9090 14418 9102
rect 14926 9154 14978 9166
rect 31166 9154 31218 9166
rect 15698 9102 15710 9154
rect 15762 9102 15774 9154
rect 14926 9090 14978 9102
rect 31166 9090 31218 9102
rect 34750 9154 34802 9166
rect 34750 9090 34802 9102
rect 14254 9042 14306 9054
rect 31838 9042 31890 9054
rect 37214 9042 37266 9054
rect 38446 9042 38498 9054
rect 13906 8990 13918 9042
rect 13970 8990 13982 9042
rect 15026 8990 15038 9042
rect 15090 8990 15102 9042
rect 15586 8990 15598 9042
rect 15650 8990 15662 9042
rect 35074 8990 35086 9042
rect 35138 8990 35150 9042
rect 37650 8990 37662 9042
rect 37714 8990 37726 9042
rect 14254 8978 14306 8990
rect 31838 8978 31890 8990
rect 37214 8978 37266 8990
rect 38446 8978 38498 8990
rect 42702 9042 42754 9054
rect 42702 8978 42754 8990
rect 43374 9042 43426 9054
rect 43374 8978 43426 8990
rect 43486 9042 43538 9054
rect 43486 8978 43538 8990
rect 44046 9042 44098 9054
rect 44046 8978 44098 8990
rect 34862 8930 34914 8942
rect 15922 8878 15934 8930
rect 15986 8878 15998 8930
rect 34862 8866 34914 8878
rect 38110 8930 38162 8942
rect 38110 8866 38162 8878
rect 42814 8930 42866 8942
rect 42814 8866 42866 8878
rect 38782 8818 38834 8830
rect 38782 8754 38834 8766
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 35086 8482 35138 8494
rect 35086 8418 35138 8430
rect 23550 8370 23602 8382
rect 15138 8318 15150 8370
rect 15202 8318 15214 8370
rect 16594 8318 16606 8370
rect 16658 8318 16670 8370
rect 18050 8318 18062 8370
rect 18114 8318 18126 8370
rect 18722 8318 18734 8370
rect 18786 8318 18798 8370
rect 20738 8318 20750 8370
rect 20802 8318 20814 8370
rect 21858 8318 21870 8370
rect 21922 8318 21934 8370
rect 31714 8318 31726 8370
rect 31778 8318 31790 8370
rect 41682 8318 41694 8370
rect 41746 8318 41758 8370
rect 23550 8306 23602 8318
rect 15710 8258 15762 8270
rect 17726 8258 17778 8270
rect 22318 8258 22370 8270
rect 14802 8206 14814 8258
rect 14866 8206 14878 8258
rect 16482 8206 16494 8258
rect 16546 8206 16558 8258
rect 18610 8206 18622 8258
rect 18674 8206 18686 8258
rect 21746 8206 21758 8258
rect 21810 8206 21822 8258
rect 15710 8194 15762 8206
rect 17726 8194 17778 8206
rect 22318 8194 22370 8206
rect 23774 8258 23826 8270
rect 23774 8194 23826 8206
rect 27358 8258 27410 8270
rect 34190 8258 34242 8270
rect 31490 8206 31502 8258
rect 31554 8206 31566 8258
rect 27358 8194 27410 8206
rect 34190 8194 34242 8206
rect 34750 8258 34802 8270
rect 35074 8206 35086 8258
rect 35138 8206 35150 8258
rect 40114 8206 40126 8258
rect 40178 8206 40190 8258
rect 34750 8194 34802 8206
rect 17390 8146 17442 8158
rect 17390 8082 17442 8094
rect 17950 8146 18002 8158
rect 17950 8082 18002 8094
rect 19518 8146 19570 8158
rect 19518 8082 19570 8094
rect 20414 8146 20466 8158
rect 20414 8082 20466 8094
rect 32174 8146 32226 8158
rect 32174 8082 32226 8094
rect 34526 8146 34578 8158
rect 34526 8082 34578 8094
rect 35422 8146 35474 8158
rect 41122 8094 41134 8146
rect 41186 8094 41198 8146
rect 35422 8082 35474 8094
rect 20638 8034 20690 8046
rect 27806 8034 27858 8046
rect 24098 7982 24110 8034
rect 24162 7982 24174 8034
rect 20638 7970 20690 7982
rect 27806 7970 27858 7982
rect 27918 8034 27970 8046
rect 27918 7970 27970 7982
rect 28030 8034 28082 8046
rect 28030 7970 28082 7982
rect 34638 8034 34690 8046
rect 39890 7982 39902 8034
rect 39954 7982 39966 8034
rect 34638 7970 34690 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 18398 7698 18450 7710
rect 31838 7698 31890 7710
rect 28690 7646 28702 7698
rect 28754 7646 28766 7698
rect 18398 7634 18450 7646
rect 31838 7634 31890 7646
rect 33406 7698 33458 7710
rect 33406 7634 33458 7646
rect 33518 7698 33570 7710
rect 33518 7634 33570 7646
rect 42030 7698 42082 7710
rect 42030 7634 42082 7646
rect 42142 7698 42194 7710
rect 42142 7634 42194 7646
rect 18622 7586 18674 7598
rect 18622 7522 18674 7534
rect 20974 7586 21026 7598
rect 20974 7522 21026 7534
rect 21310 7586 21362 7598
rect 21310 7522 21362 7534
rect 21870 7586 21922 7598
rect 32062 7586 32114 7598
rect 26338 7534 26350 7586
rect 26402 7534 26414 7586
rect 21870 7522 21922 7534
rect 32062 7522 32114 7534
rect 21646 7474 21698 7486
rect 26910 7474 26962 7486
rect 28142 7474 28194 7486
rect 20290 7422 20302 7474
rect 20354 7422 20366 7474
rect 23762 7422 23774 7474
rect 23826 7422 23838 7474
rect 25218 7422 25230 7474
rect 25282 7422 25294 7474
rect 25778 7422 25790 7474
rect 25842 7422 25854 7474
rect 27346 7422 27358 7474
rect 27410 7422 27422 7474
rect 21646 7410 21698 7422
rect 26910 7410 26962 7422
rect 28142 7410 28194 7422
rect 28366 7474 28418 7486
rect 28366 7410 28418 7422
rect 32174 7474 32226 7486
rect 32174 7410 32226 7422
rect 32958 7474 33010 7486
rect 32958 7410 33010 7422
rect 33630 7474 33682 7486
rect 33630 7410 33682 7422
rect 41470 7474 41522 7486
rect 41470 7410 41522 7422
rect 41918 7474 41970 7486
rect 41918 7410 41970 7422
rect 21758 7362 21810 7374
rect 27806 7362 27858 7374
rect 18386 7310 18398 7362
rect 18450 7310 18462 7362
rect 20514 7310 20526 7362
rect 20578 7310 20590 7362
rect 23874 7310 23886 7362
rect 23938 7310 23950 7362
rect 25666 7310 25678 7362
rect 25730 7310 25742 7362
rect 21758 7298 21810 7310
rect 27806 7298 27858 7310
rect 24546 7198 24558 7250
rect 24610 7198 24622 7250
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 13694 6914 13746 6926
rect 13694 6850 13746 6862
rect 23998 6914 24050 6926
rect 23998 6850 24050 6862
rect 27246 6914 27298 6926
rect 27246 6850 27298 6862
rect 27582 6914 27634 6926
rect 27582 6850 27634 6862
rect 23774 6802 23826 6814
rect 23774 6738 23826 6750
rect 26574 6802 26626 6814
rect 26574 6738 26626 6750
rect 27806 6802 27858 6814
rect 27806 6738 27858 6750
rect 33854 6802 33906 6814
rect 33854 6738 33906 6750
rect 34526 6802 34578 6814
rect 34526 6738 34578 6750
rect 39566 6802 39618 6814
rect 39566 6738 39618 6750
rect 13470 6690 13522 6702
rect 13470 6626 13522 6638
rect 15934 6690 15986 6702
rect 15934 6626 15986 6638
rect 16382 6690 16434 6702
rect 18734 6690 18786 6702
rect 29710 6690 29762 6702
rect 31278 6690 31330 6702
rect 18162 6638 18174 6690
rect 18226 6638 18238 6690
rect 24322 6638 24334 6690
rect 24386 6638 24398 6690
rect 30146 6638 30158 6690
rect 30210 6638 30222 6690
rect 16382 6626 16434 6638
rect 18734 6626 18786 6638
rect 29710 6626 29762 6638
rect 31278 6626 31330 6638
rect 31614 6690 31666 6702
rect 31614 6626 31666 6638
rect 31838 6690 31890 6702
rect 34414 6690 34466 6702
rect 42254 6690 42306 6702
rect 46734 6690 46786 6702
rect 32386 6638 32398 6690
rect 32450 6638 32462 6690
rect 37650 6638 37662 6690
rect 37714 6638 37726 6690
rect 38546 6638 38558 6690
rect 38610 6638 38622 6690
rect 41122 6638 41134 6690
rect 41186 6638 41198 6690
rect 42578 6638 42590 6690
rect 42642 6638 42654 6690
rect 46946 6638 46958 6690
rect 47010 6638 47022 6690
rect 31838 6626 31890 6638
rect 34414 6626 34466 6638
rect 42254 6626 42306 6638
rect 46734 6626 46786 6638
rect 31390 6578 31442 6590
rect 34638 6578 34690 6590
rect 33394 6526 33406 6578
rect 33458 6526 33470 6578
rect 31390 6514 31442 6526
rect 34638 6514 34690 6526
rect 35310 6578 35362 6590
rect 35310 6514 35362 6526
rect 35646 6578 35698 6590
rect 35646 6514 35698 6526
rect 35870 6578 35922 6590
rect 42142 6578 42194 6590
rect 37314 6526 37326 6578
rect 37378 6526 37390 6578
rect 39890 6526 39902 6578
rect 39954 6526 39966 6578
rect 41458 6526 41470 6578
rect 41522 6526 41534 6578
rect 48066 6526 48078 6578
rect 48130 6526 48142 6578
rect 35870 6514 35922 6526
rect 42142 6514 42194 6526
rect 15710 6466 15762 6478
rect 14018 6414 14030 6466
rect 14082 6414 14094 6466
rect 15710 6402 15762 6414
rect 15822 6466 15874 6478
rect 15822 6402 15874 6414
rect 18510 6466 18562 6478
rect 18510 6402 18562 6414
rect 18622 6466 18674 6478
rect 18622 6402 18674 6414
rect 29598 6466 29650 6478
rect 29598 6402 29650 6414
rect 29822 6466 29874 6478
rect 29822 6402 29874 6414
rect 35422 6466 35474 6478
rect 35422 6402 35474 6414
rect 36430 6466 36482 6478
rect 38882 6414 38894 6466
rect 38946 6414 38958 6466
rect 36430 6402 36482 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 16494 6130 16546 6142
rect 16494 6066 16546 6078
rect 20302 6130 20354 6142
rect 33182 6130 33234 6142
rect 38894 6130 38946 6142
rect 30258 6078 30270 6130
rect 30322 6078 30334 6130
rect 35522 6078 35534 6130
rect 35586 6078 35598 6130
rect 20302 6066 20354 6078
rect 33182 6066 33234 6078
rect 38894 6066 38946 6078
rect 39566 6130 39618 6142
rect 39566 6066 39618 6078
rect 41358 6130 41410 6142
rect 41358 6066 41410 6078
rect 16718 6018 16770 6030
rect 13570 5966 13582 6018
rect 13634 5966 13646 6018
rect 16718 5954 16770 5966
rect 16830 6018 16882 6030
rect 16830 5954 16882 5966
rect 18398 6018 18450 6030
rect 18398 5954 18450 5966
rect 20862 6018 20914 6030
rect 20862 5954 20914 5966
rect 26238 6018 26290 6030
rect 32510 6018 32562 6030
rect 39118 6018 39170 6030
rect 28690 5966 28702 6018
rect 28754 5966 28766 6018
rect 33842 5966 33854 6018
rect 33906 5966 33918 6018
rect 26238 5954 26290 5966
rect 32510 5954 32562 5966
rect 39118 5954 39170 5966
rect 41582 6018 41634 6030
rect 41582 5954 41634 5966
rect 43038 6018 43090 6030
rect 43038 5954 43090 5966
rect 14254 5906 14306 5918
rect 16270 5906 16322 5918
rect 18734 5906 18786 5918
rect 13458 5854 13470 5906
rect 13522 5854 13534 5906
rect 15586 5854 15598 5906
rect 15650 5854 15662 5906
rect 17714 5854 17726 5906
rect 17778 5854 17790 5906
rect 14254 5842 14306 5854
rect 16270 5842 16322 5854
rect 18734 5842 18786 5854
rect 18958 5906 19010 5918
rect 18958 5842 19010 5854
rect 19182 5906 19234 5918
rect 19182 5842 19234 5854
rect 20414 5906 20466 5918
rect 20414 5842 20466 5854
rect 20638 5906 20690 5918
rect 20638 5842 20690 5854
rect 20974 5906 21026 5918
rect 22878 5906 22930 5918
rect 36094 5906 36146 5918
rect 37550 5906 37602 5918
rect 39342 5906 39394 5918
rect 22306 5854 22318 5906
rect 22370 5854 22382 5906
rect 25666 5854 25678 5906
rect 25730 5854 25742 5906
rect 29250 5854 29262 5906
rect 29314 5854 29326 5906
rect 29922 5854 29934 5906
rect 29986 5854 29998 5906
rect 31938 5854 31950 5906
rect 32002 5854 32014 5906
rect 35298 5854 35310 5906
rect 35362 5854 35374 5906
rect 36642 5854 36654 5906
rect 36706 5854 36718 5906
rect 37874 5854 37886 5906
rect 37938 5854 37950 5906
rect 20974 5842 21026 5854
rect 22878 5842 22930 5854
rect 36094 5842 36146 5854
rect 37550 5842 37602 5854
rect 39342 5842 39394 5854
rect 39678 5906 39730 5918
rect 39678 5842 39730 5854
rect 41694 5906 41746 5918
rect 41694 5842 41746 5854
rect 42142 5906 42194 5918
rect 42354 5854 42366 5906
rect 42418 5854 42430 5906
rect 42142 5842 42194 5854
rect 22990 5794 23042 5806
rect 37438 5794 37490 5806
rect 15810 5742 15822 5794
rect 15874 5742 15886 5794
rect 17602 5742 17614 5794
rect 17666 5742 17678 5794
rect 25330 5742 25342 5794
rect 25394 5742 25406 5794
rect 32162 5742 32174 5794
rect 32226 5742 32238 5794
rect 33618 5742 33630 5794
rect 33682 5742 33694 5794
rect 36866 5742 36878 5794
rect 36930 5742 36942 5794
rect 22990 5730 23042 5742
rect 37438 5730 37490 5742
rect 14590 5682 14642 5694
rect 14590 5618 14642 5630
rect 19630 5682 19682 5694
rect 19630 5618 19682 5630
rect 20302 5682 20354 5694
rect 20302 5618 20354 5630
rect 38782 5682 38834 5694
rect 38782 5618 38834 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 18958 5346 19010 5358
rect 24994 5294 25006 5346
rect 25058 5294 25070 5346
rect 34962 5294 34974 5346
rect 35026 5294 35038 5346
rect 18958 5282 19010 5294
rect 15038 5234 15090 5246
rect 14578 5182 14590 5234
rect 14642 5182 14654 5234
rect 15038 5170 15090 5182
rect 15934 5234 15986 5246
rect 15934 5170 15986 5182
rect 18734 5234 18786 5246
rect 26014 5234 26066 5246
rect 20514 5182 20526 5234
rect 20578 5182 20590 5234
rect 21522 5182 21534 5234
rect 21586 5182 21598 5234
rect 23090 5182 23102 5234
rect 23154 5182 23166 5234
rect 18734 5170 18786 5182
rect 26014 5170 26066 5182
rect 29486 5234 29538 5246
rect 37214 5234 37266 5246
rect 35522 5182 35534 5234
rect 35586 5182 35598 5234
rect 29486 5170 29538 5182
rect 37214 5170 37266 5182
rect 38894 5234 38946 5246
rect 38894 5170 38946 5182
rect 40910 5234 40962 5246
rect 40910 5170 40962 5182
rect 46622 5234 46674 5246
rect 46622 5170 46674 5182
rect 20750 5122 20802 5134
rect 22430 5122 22482 5134
rect 37774 5122 37826 5134
rect 14354 5070 14366 5122
rect 14418 5070 14430 5122
rect 17266 5070 17278 5122
rect 17330 5070 17342 5122
rect 19282 5070 19294 5122
rect 19346 5070 19358 5122
rect 19842 5070 19854 5122
rect 19906 5070 19918 5122
rect 21746 5070 21758 5122
rect 21810 5070 21822 5122
rect 23314 5070 23326 5122
rect 23378 5070 23390 5122
rect 24322 5070 24334 5122
rect 24386 5070 24398 5122
rect 27570 5070 27582 5122
rect 27634 5070 27646 5122
rect 30594 5070 30606 5122
rect 30658 5070 30670 5122
rect 31490 5070 31502 5122
rect 31554 5070 31566 5122
rect 35634 5070 35646 5122
rect 35698 5070 35710 5122
rect 20750 5058 20802 5070
rect 22430 5058 22482 5070
rect 37774 5058 37826 5070
rect 37998 5122 38050 5134
rect 37998 5058 38050 5070
rect 38334 5122 38386 5134
rect 46958 5122 47010 5134
rect 40450 5070 40462 5122
rect 40514 5070 40526 5122
rect 38334 5058 38386 5070
rect 46958 5058 47010 5070
rect 47742 5122 47794 5134
rect 47742 5058 47794 5070
rect 17950 5010 18002 5022
rect 28030 5010 28082 5022
rect 16146 4958 16158 5010
rect 16210 4958 16222 5010
rect 26114 4958 26126 5010
rect 26178 4958 26190 5010
rect 17950 4946 18002 4958
rect 28030 4946 28082 4958
rect 29374 5010 29426 5022
rect 29374 4946 29426 4958
rect 29598 5010 29650 5022
rect 38110 5010 38162 5022
rect 30370 4958 30382 5010
rect 30434 4958 30446 5010
rect 38994 4958 39006 5010
rect 39058 4958 39070 5010
rect 29598 4946 29650 4958
rect 38110 4946 38162 4958
rect 31938 4846 31950 4898
rect 32002 4846 32014 4898
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 23662 4562 23714 4574
rect 19730 4510 19742 4562
rect 19794 4510 19806 4562
rect 23662 4498 23714 4510
rect 23774 4562 23826 4574
rect 23774 4498 23826 4510
rect 30046 4562 30098 4574
rect 30046 4498 30098 4510
rect 35982 4562 36034 4574
rect 35982 4498 36034 4510
rect 38670 4562 38722 4574
rect 38670 4498 38722 4510
rect 38894 4562 38946 4574
rect 38894 4498 38946 4510
rect 39566 4562 39618 4574
rect 39566 4498 39618 4510
rect 14702 4450 14754 4462
rect 14702 4386 14754 4398
rect 22094 4450 22146 4462
rect 29934 4450 29986 4462
rect 25890 4398 25902 4450
rect 25954 4398 25966 4450
rect 22094 4386 22146 4398
rect 29934 4386 29986 4398
rect 30494 4450 30546 4462
rect 30494 4386 30546 4398
rect 35870 4450 35922 4462
rect 35870 4386 35922 4398
rect 46622 4450 46674 4462
rect 46622 4386 46674 4398
rect 14366 4338 14418 4350
rect 14018 4286 14030 4338
rect 14082 4286 14094 4338
rect 14366 4274 14418 4286
rect 22318 4338 22370 4350
rect 22318 4274 22370 4286
rect 23102 4338 23154 4350
rect 23102 4274 23154 4286
rect 23550 4338 23602 4350
rect 27470 4338 27522 4350
rect 27010 4286 27022 4338
rect 27074 4286 27086 4338
rect 23550 4274 23602 4286
rect 27470 4274 27522 4286
rect 30606 4338 30658 4350
rect 30606 4274 30658 4286
rect 38782 4338 38834 4350
rect 39678 4338 39730 4350
rect 39218 4286 39230 4338
rect 39282 4286 39294 4338
rect 46946 4286 46958 4338
rect 47010 4286 47022 4338
rect 38782 4274 38834 4286
rect 39678 4274 39730 4286
rect 13470 4226 13522 4238
rect 13470 4162 13522 4174
rect 18958 4226 19010 4238
rect 18958 4162 19010 4174
rect 19182 4226 19234 4238
rect 19182 4162 19234 4174
rect 22654 4226 22706 4238
rect 25330 4174 25342 4226
rect 25394 4174 25406 4226
rect 48066 4174 48078 4226
rect 48130 4174 48142 4226
rect 22654 4162 22706 4174
rect 13694 4114 13746 4126
rect 13694 4050 13746 4062
rect 19406 4114 19458 4126
rect 19406 4050 19458 4062
rect 30046 4114 30098 4126
rect 30046 4050 30098 4062
rect 36094 4114 36146 4126
rect 36094 4050 36146 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 45278 3666 45330 3678
rect 22978 3614 22990 3666
rect 23042 3614 23054 3666
rect 40226 3614 40238 3666
rect 40290 3614 40302 3666
rect 44034 3614 44046 3666
rect 44098 3614 44110 3666
rect 45278 3602 45330 3614
rect 26910 3554 26962 3566
rect 45614 3554 45666 3566
rect 27346 3502 27358 3554
rect 27410 3502 27422 3554
rect 31378 3502 31390 3554
rect 31442 3502 31454 3554
rect 26910 3490 26962 3502
rect 45614 3490 45666 3502
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 2942 3442 2994 3454
rect 2942 3378 2994 3390
rect 3278 3442 3330 3454
rect 3278 3378 3330 3390
rect 6750 3442 6802 3454
rect 6750 3378 6802 3390
rect 6974 3442 7026 3454
rect 10782 3442 10834 3454
rect 7298 3390 7310 3442
rect 7362 3390 7374 3442
rect 6974 3378 7026 3390
rect 10782 3378 10834 3390
rect 11006 3442 11058 3454
rect 11006 3378 11058 3390
rect 11342 3442 11394 3454
rect 11342 3378 11394 3390
rect 14814 3442 14866 3454
rect 14814 3378 14866 3390
rect 15038 3442 15090 3454
rect 15038 3378 15090 3390
rect 15374 3442 15426 3454
rect 15374 3378 15426 3390
rect 18846 3442 18898 3454
rect 18846 3378 18898 3390
rect 19070 3442 19122 3454
rect 19070 3378 19122 3390
rect 19406 3442 19458 3454
rect 19406 3378 19458 3390
rect 23438 3442 23490 3454
rect 23438 3378 23490 3390
rect 23886 3442 23938 3454
rect 23886 3378 23938 3390
rect 28478 3442 28530 3454
rect 28478 3378 28530 3390
rect 30942 3442 30994 3454
rect 30942 3378 30994 3390
rect 39342 3442 39394 3454
rect 39342 3378 39394 3390
rect 39790 3442 39842 3454
rect 39790 3378 39842 3390
rect 43150 3442 43202 3454
rect 43150 3378 43202 3390
rect 43598 3442 43650 3454
rect 43598 3378 43650 3390
rect 46398 3442 46450 3454
rect 46398 3378 46450 3390
rect 31154 3278 31166 3330
rect 31218 3278 31230 3330
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 16830 76974 16882 77026
rect 17950 76974 18002 77026
rect 18622 76974 18674 77026
rect 19182 76974 19234 77026
rect 20414 76974 20466 77026
rect 21534 76974 21586 77026
rect 22206 76974 22258 77026
rect 23102 76974 23154 77026
rect 25790 76974 25842 77026
rect 26350 76974 26402 77026
rect 43710 76974 43762 77026
rect 44270 76974 44322 77026
rect 44718 76974 44770 77026
rect 45502 76974 45554 77026
rect 46062 76974 46114 77026
rect 46510 76974 46562 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 10222 76638 10274 76690
rect 11790 76638 11842 76690
rect 21534 76638 21586 76690
rect 30382 76638 30434 76690
rect 32622 76638 32674 76690
rect 37550 76638 37602 76690
rect 42926 76638 42978 76690
rect 44270 76638 44322 76690
rect 44718 76638 44770 76690
rect 46062 76638 46114 76690
rect 46510 76638 46562 76690
rect 48190 76638 48242 76690
rect 2494 76526 2546 76578
rect 7870 76526 7922 76578
rect 17950 76526 18002 76578
rect 19182 76526 19234 76578
rect 26350 76526 26402 76578
rect 36094 76526 36146 76578
rect 41470 76526 41522 76578
rect 3278 76414 3330 76466
rect 3726 76414 3778 76466
rect 6974 76414 7026 76466
rect 8766 76414 8818 76466
rect 10894 76414 10946 76466
rect 12462 76414 12514 76466
rect 13470 76414 13522 76466
rect 15150 76414 15202 76466
rect 17054 76414 17106 76466
rect 20078 76414 20130 76466
rect 20750 76414 20802 76466
rect 22430 76414 22482 76466
rect 27246 76414 27298 76466
rect 28814 76414 28866 76466
rect 31166 76414 31218 76466
rect 33406 76414 33458 76466
rect 35086 76414 35138 76466
rect 36990 76414 37042 76466
rect 38782 76414 38834 76466
rect 40798 76414 40850 76466
rect 42366 76414 42418 76466
rect 43710 76414 43762 76466
rect 4398 76302 4450 76354
rect 6190 76302 6242 76354
rect 13918 76302 13970 76354
rect 15598 76302 15650 76354
rect 22094 76302 22146 76354
rect 23102 76302 23154 76354
rect 29262 76302 29314 76354
rect 36542 76302 36594 76354
rect 38334 76302 38386 76354
rect 42030 76302 42082 76354
rect 45502 76302 45554 76354
rect 34302 76190 34354 76242
rect 40014 76190 40066 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 3614 75742 3666 75794
rect 19070 75742 19122 75794
rect 24446 75742 24498 75794
rect 34750 75742 34802 75794
rect 39118 75742 39170 75794
rect 2606 75630 2658 75682
rect 3166 75630 3218 75682
rect 9102 75630 9154 75682
rect 20526 75630 20578 75682
rect 25454 75630 25506 75682
rect 29262 75630 29314 75682
rect 31502 75630 31554 75682
rect 31950 75630 32002 75682
rect 1710 75518 1762 75570
rect 2270 75518 2322 75570
rect 15934 75518 15986 75570
rect 16270 75518 16322 75570
rect 32622 75518 32674 75570
rect 48190 75518 48242 75570
rect 13694 75406 13746 75458
rect 17054 75406 17106 75458
rect 26014 75406 26066 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 33294 75070 33346 75122
rect 33518 75070 33570 75122
rect 4062 74958 4114 75010
rect 5406 74958 5458 75010
rect 6638 74958 6690 75010
rect 14702 74958 14754 75010
rect 25230 74958 25282 75010
rect 4846 74846 4898 74898
rect 5854 74846 5906 74898
rect 10670 74846 10722 74898
rect 14030 74846 14082 74898
rect 17390 74846 17442 74898
rect 23550 74846 23602 74898
rect 23998 74846 24050 74898
rect 24670 74846 24722 74898
rect 25454 74846 25506 74898
rect 26014 74846 26066 74898
rect 31950 74846 32002 74898
rect 1934 74734 1986 74786
rect 8766 74734 8818 74786
rect 9662 74734 9714 74786
rect 11342 74734 11394 74786
rect 13470 74734 13522 74786
rect 16830 74734 16882 74786
rect 18174 74734 18226 74786
rect 20302 74734 20354 74786
rect 20638 74734 20690 74786
rect 22766 74734 22818 74786
rect 26686 74734 26738 74786
rect 28814 74734 28866 74786
rect 29150 74734 29202 74786
rect 31278 74734 31330 74786
rect 33966 74734 34018 74786
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 1822 74174 1874 74226
rect 12014 74174 12066 74226
rect 13470 74174 13522 74226
rect 15598 74174 15650 74226
rect 20190 74174 20242 74226
rect 22318 74174 22370 74226
rect 22766 74174 22818 74226
rect 23886 74174 23938 74226
rect 26014 74174 26066 74226
rect 32398 74174 32450 74226
rect 3950 74062 4002 74114
rect 9102 74062 9154 74114
rect 16382 74062 16434 74114
rect 17614 74062 17666 74114
rect 18174 74062 18226 74114
rect 23214 74062 23266 74114
rect 26574 74062 26626 74114
rect 29598 74062 29650 74114
rect 33294 74062 33346 74114
rect 3390 73950 3442 74002
rect 4734 73950 4786 74002
rect 5742 73950 5794 74002
rect 9886 73950 9938 74002
rect 12462 73950 12514 74002
rect 16830 73950 16882 74002
rect 18846 73950 18898 74002
rect 19406 73950 19458 74002
rect 19742 73950 19794 74002
rect 20750 73950 20802 74002
rect 26350 73950 26402 74002
rect 27246 73950 27298 74002
rect 27582 73950 27634 74002
rect 28254 73950 28306 74002
rect 28590 73950 28642 74002
rect 30270 73950 30322 74002
rect 33070 73950 33122 74002
rect 4174 73838 4226 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 10334 73502 10386 73554
rect 23102 73502 23154 73554
rect 27694 73502 27746 73554
rect 29150 73502 29202 73554
rect 30606 73502 30658 73554
rect 9550 73390 9602 73442
rect 25454 73390 25506 73442
rect 48190 73390 48242 73442
rect 1710 73278 1762 73330
rect 4062 73278 4114 73330
rect 9886 73278 9938 73330
rect 10670 73278 10722 73330
rect 13806 73278 13858 73330
rect 18622 73278 18674 73330
rect 19182 73278 19234 73330
rect 20302 73278 20354 73330
rect 20638 73278 20690 73330
rect 21982 73278 22034 73330
rect 22430 73278 22482 73330
rect 23886 73278 23938 73330
rect 24334 73278 24386 73330
rect 25678 73278 25730 73330
rect 28030 73278 28082 73330
rect 30830 73278 30882 73330
rect 2270 73166 2322 73218
rect 4846 73166 4898 73218
rect 6974 73166 7026 73218
rect 7422 73166 7474 73218
rect 9102 73166 9154 73218
rect 11118 73166 11170 73218
rect 14478 73166 14530 73218
rect 16606 73166 16658 73218
rect 17950 73166 18002 73218
rect 19294 73166 19346 73218
rect 21310 73166 21362 73218
rect 22654 73166 22706 73218
rect 23662 73166 23714 73218
rect 26238 73166 26290 73218
rect 26686 73166 26738 73218
rect 28478 73166 28530 73218
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 10670 72718 10722 72770
rect 11006 72718 11058 72770
rect 1822 72606 1874 72658
rect 8318 72606 8370 72658
rect 10446 72606 10498 72658
rect 10894 72606 10946 72658
rect 17166 72606 17218 72658
rect 18174 72606 18226 72658
rect 18958 72606 19010 72658
rect 20638 72606 20690 72658
rect 22430 72606 22482 72658
rect 25678 72606 25730 72658
rect 30494 72606 30546 72658
rect 33182 72606 33234 72658
rect 5854 72494 5906 72546
rect 7534 72494 7586 72546
rect 18734 72494 18786 72546
rect 20302 72494 20354 72546
rect 22206 72494 22258 72546
rect 23998 72494 24050 72546
rect 24558 72494 24610 72546
rect 31166 72494 31218 72546
rect 31390 72494 31442 72546
rect 32510 72494 32562 72546
rect 33070 72494 33122 72546
rect 33854 72494 33906 72546
rect 34078 72494 34130 72546
rect 5630 72382 5682 72434
rect 6526 72382 6578 72434
rect 19406 72382 19458 72434
rect 19742 72382 19794 72434
rect 21646 72382 21698 72434
rect 22878 72382 22930 72434
rect 25118 72382 25170 72434
rect 33518 72382 33570 72434
rect 17054 72270 17106 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 25342 71934 25394 71986
rect 31166 71934 31218 71986
rect 31950 71934 32002 71986
rect 18734 71822 18786 71874
rect 20750 71822 20802 71874
rect 29822 71822 29874 71874
rect 30494 71822 30546 71874
rect 31390 71822 31442 71874
rect 32174 71822 32226 71874
rect 32286 71822 32338 71874
rect 19742 71710 19794 71762
rect 21870 71710 21922 71762
rect 22654 71710 22706 71762
rect 24334 71710 24386 71762
rect 30046 71710 30098 71762
rect 30718 71710 30770 71762
rect 33854 71710 33906 71762
rect 35086 71710 35138 71762
rect 35646 71710 35698 71762
rect 35870 71710 35922 71762
rect 37102 71710 37154 71762
rect 37550 71710 37602 71762
rect 37774 71710 37826 71762
rect 18510 71598 18562 71650
rect 22766 71598 22818 71650
rect 23774 71598 23826 71650
rect 30270 71598 30322 71650
rect 31054 71598 31106 71650
rect 33182 71598 33234 71650
rect 34078 71598 34130 71650
rect 35758 71598 35810 71650
rect 37326 71598 37378 71650
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 19854 71150 19906 71202
rect 32510 71150 32562 71202
rect 35870 71150 35922 71202
rect 6302 71038 6354 71090
rect 9214 71038 9266 71090
rect 12798 71038 12850 71090
rect 16606 71038 16658 71090
rect 18958 71038 19010 71090
rect 23102 71038 23154 71090
rect 26462 71038 26514 71090
rect 31390 71038 31442 71090
rect 8430 70926 8482 70978
rect 9998 70926 10050 70978
rect 13694 70926 13746 70978
rect 17838 70926 17890 70978
rect 18286 70926 18338 70978
rect 19630 70926 19682 70978
rect 20078 70926 20130 70978
rect 22430 70926 22482 70978
rect 24558 70926 24610 70978
rect 26574 70926 26626 70978
rect 26910 70926 26962 70978
rect 29934 70926 29986 70978
rect 30942 70926 30994 70978
rect 32958 70926 33010 70978
rect 33182 70926 33234 70978
rect 33406 70926 33458 70978
rect 33966 70926 34018 70978
rect 34862 70926 34914 70978
rect 35982 70926 36034 70978
rect 37998 70926 38050 70978
rect 38558 70926 38610 70978
rect 2270 70814 2322 70866
rect 8206 70814 8258 70866
rect 10670 70814 10722 70866
rect 14478 70814 14530 70866
rect 19406 70814 19458 70866
rect 20526 70814 20578 70866
rect 23550 70814 23602 70866
rect 25006 70814 25058 70866
rect 29486 70814 29538 70866
rect 36990 70814 37042 70866
rect 1710 70702 1762 70754
rect 6190 70702 6242 70754
rect 6974 70702 7026 70754
rect 7422 70702 7474 70754
rect 8654 70702 8706 70754
rect 8766 70702 8818 70754
rect 17166 70702 17218 70754
rect 21422 70702 21474 70754
rect 28702 70702 28754 70754
rect 39118 70702 39170 70754
rect 48190 70702 48242 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 1822 70366 1874 70418
rect 7646 70366 7698 70418
rect 10446 70366 10498 70418
rect 22430 70366 22482 70418
rect 25902 70366 25954 70418
rect 34974 70366 35026 70418
rect 35086 70366 35138 70418
rect 38894 70366 38946 70418
rect 8766 70254 8818 70306
rect 8990 70254 9042 70306
rect 18398 70254 18450 70306
rect 19742 70254 19794 70306
rect 20190 70254 20242 70306
rect 24558 70254 24610 70306
rect 26014 70254 26066 70306
rect 26462 70254 26514 70306
rect 28478 70254 28530 70306
rect 30046 70254 30098 70306
rect 33966 70254 34018 70306
rect 35534 70254 35586 70306
rect 37774 70254 37826 70306
rect 39006 70254 39058 70306
rect 7198 70142 7250 70194
rect 8206 70142 8258 70194
rect 10222 70142 10274 70194
rect 12462 70142 12514 70194
rect 17726 70142 17778 70194
rect 18286 70142 18338 70194
rect 19070 70142 19122 70194
rect 21310 70142 21362 70194
rect 21870 70142 21922 70194
rect 23662 70142 23714 70194
rect 27134 70142 27186 70194
rect 27358 70142 27410 70194
rect 29038 70142 29090 70194
rect 30494 70142 30546 70194
rect 30942 70142 30994 70194
rect 32958 70142 33010 70194
rect 33742 70142 33794 70194
rect 36878 70142 36930 70194
rect 37662 70142 37714 70194
rect 39566 70142 39618 70194
rect 4286 70030 4338 70082
rect 6414 70030 6466 70082
rect 8654 70030 8706 70082
rect 9774 70030 9826 70082
rect 13134 70030 13186 70082
rect 15262 70030 15314 70082
rect 16830 70030 16882 70082
rect 19294 70030 19346 70082
rect 20638 70030 20690 70082
rect 21982 70030 22034 70082
rect 23550 70030 23602 70082
rect 25454 70030 25506 70082
rect 29374 70030 29426 70082
rect 33630 70030 33682 70082
rect 8430 69918 8482 69970
rect 25790 69918 25842 69970
rect 35198 69918 35250 69970
rect 38782 69918 38834 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 22542 69582 22594 69634
rect 22766 69582 22818 69634
rect 23438 69582 23490 69634
rect 27806 69582 27858 69634
rect 29374 69582 29426 69634
rect 33406 69582 33458 69634
rect 36430 69582 36482 69634
rect 38446 69582 38498 69634
rect 12798 69470 12850 69522
rect 17054 69470 17106 69522
rect 17502 69470 17554 69522
rect 17726 69470 17778 69522
rect 18734 69470 18786 69522
rect 25006 69470 25058 69522
rect 25902 69470 25954 69522
rect 28030 69470 28082 69522
rect 29710 69470 29762 69522
rect 35646 69470 35698 69522
rect 37998 69470 38050 69522
rect 39118 69470 39170 69522
rect 41806 69470 41858 69522
rect 6190 69358 6242 69410
rect 6414 69358 6466 69410
rect 8430 69358 8482 69410
rect 8766 69358 8818 69410
rect 9998 69358 10050 69410
rect 14142 69358 14194 69410
rect 22318 69358 22370 69410
rect 22990 69358 23042 69410
rect 25678 69358 25730 69410
rect 26574 69358 26626 69410
rect 26798 69358 26850 69410
rect 33406 69358 33458 69410
rect 37102 69358 37154 69410
rect 37326 69358 37378 69410
rect 39230 69358 39282 69410
rect 42254 69358 42306 69410
rect 42702 69358 42754 69410
rect 6638 69246 6690 69298
rect 7982 69246 8034 69298
rect 10670 69246 10722 69298
rect 14926 69246 14978 69298
rect 27134 69246 27186 69298
rect 27470 69246 27522 69298
rect 29598 69246 29650 69298
rect 33070 69246 33122 69298
rect 36318 69246 36370 69298
rect 5854 69134 5906 69186
rect 7086 69134 7138 69186
rect 24222 69134 24274 69186
rect 24670 69134 24722 69186
rect 26686 69134 26738 69186
rect 35198 69134 35250 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 27134 68798 27186 68850
rect 33742 68798 33794 68850
rect 6414 68686 6466 68738
rect 8094 68674 8146 68726
rect 23438 68686 23490 68738
rect 25454 68686 25506 68738
rect 34302 68686 34354 68738
rect 48190 68686 48242 68738
rect 1822 68574 1874 68626
rect 5854 68574 5906 68626
rect 6078 68574 6130 68626
rect 8318 68574 8370 68626
rect 9550 68574 9602 68626
rect 23886 68574 23938 68626
rect 24334 68574 24386 68626
rect 26126 68574 26178 68626
rect 33630 68574 33682 68626
rect 34190 68574 34242 68626
rect 38670 68574 38722 68626
rect 39566 68574 39618 68626
rect 2270 68462 2322 68514
rect 5966 68462 6018 68514
rect 7310 68462 7362 68514
rect 7982 68462 8034 68514
rect 9998 68462 10050 68514
rect 26238 68462 26290 68514
rect 27918 68462 27970 68514
rect 35198 68462 35250 68514
rect 35758 68462 35810 68514
rect 39118 68462 39170 68514
rect 40014 68462 40066 68514
rect 35086 68350 35138 68402
rect 38782 68350 38834 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 24334 68014 24386 68066
rect 24782 68014 24834 68066
rect 1822 67902 1874 67954
rect 6638 67902 6690 67954
rect 7646 67902 7698 67954
rect 8206 67902 8258 67954
rect 20750 67902 20802 67954
rect 24782 67902 24834 67954
rect 29150 67902 29202 67954
rect 34078 67902 34130 67954
rect 39790 67902 39842 67954
rect 40462 67902 40514 67954
rect 7198 67790 7250 67842
rect 10110 67790 10162 67842
rect 17390 67790 17442 67842
rect 17950 67790 18002 67842
rect 26238 67790 26290 67842
rect 26462 67790 26514 67842
rect 26798 67790 26850 67842
rect 27022 67790 27074 67842
rect 27358 67790 27410 67842
rect 29822 67790 29874 67842
rect 30046 67790 30098 67842
rect 32398 67790 32450 67842
rect 32958 67790 33010 67842
rect 34414 67790 34466 67842
rect 35758 67790 35810 67842
rect 39118 67790 39170 67842
rect 39342 67790 39394 67842
rect 39678 67790 39730 67842
rect 40574 67790 40626 67842
rect 43150 67790 43202 67842
rect 7534 67678 7586 67730
rect 10334 67678 10386 67730
rect 18622 67678 18674 67730
rect 33070 67678 33122 67730
rect 33406 67678 33458 67730
rect 40910 67678 40962 67730
rect 43598 67678 43650 67730
rect 43822 67678 43874 67730
rect 7758 67566 7810 67618
rect 15262 67566 15314 67618
rect 17390 67566 17442 67618
rect 26350 67566 26402 67618
rect 27246 67566 27298 67618
rect 27918 67566 27970 67618
rect 28366 67566 28418 67618
rect 30718 67566 30770 67618
rect 31054 67566 31106 67618
rect 31726 67566 31778 67618
rect 43486 67566 43538 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 14590 67230 14642 67282
rect 36206 67230 36258 67282
rect 39230 67230 39282 67282
rect 6750 67118 6802 67170
rect 18622 67118 18674 67170
rect 23326 67118 23378 67170
rect 30830 67118 30882 67170
rect 33182 67118 33234 67170
rect 33406 67118 33458 67170
rect 34078 67118 34130 67170
rect 36318 67118 36370 67170
rect 41022 67118 41074 67170
rect 42926 67118 42978 67170
rect 7086 67006 7138 67058
rect 9886 67006 9938 67058
rect 13918 67006 13970 67058
rect 14478 67006 14530 67058
rect 14814 67006 14866 67058
rect 15038 67006 15090 67058
rect 18286 67006 18338 67058
rect 20638 67006 20690 67058
rect 26686 67006 26738 67058
rect 27694 67006 27746 67058
rect 28366 67006 28418 67058
rect 29150 67006 29202 67058
rect 30270 67006 30322 67058
rect 30718 67006 30770 67058
rect 33070 67006 33122 67058
rect 35310 67006 35362 67058
rect 35646 67006 35698 67058
rect 36094 67006 36146 67058
rect 39006 67006 39058 67058
rect 39118 67006 39170 67058
rect 39454 67006 39506 67058
rect 41918 67006 41970 67058
rect 43374 67006 43426 67058
rect 44382 67006 44434 67058
rect 44606 67006 44658 67058
rect 10558 66894 10610 66946
rect 12686 66894 12738 66946
rect 15486 66894 15538 66946
rect 15934 66894 15986 66946
rect 20750 66894 20802 66946
rect 22990 66894 23042 66946
rect 25454 66894 25506 66946
rect 26574 66894 26626 66946
rect 30830 66894 30882 66946
rect 31838 66894 31890 66946
rect 41358 66894 41410 66946
rect 43262 66894 43314 66946
rect 14478 66782 14530 66834
rect 26238 66782 26290 66834
rect 29374 66782 29426 66834
rect 44270 66782 44322 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 12238 66446 12290 66498
rect 14142 66446 14194 66498
rect 14702 66446 14754 66498
rect 35646 66446 35698 66498
rect 37550 66446 37602 66498
rect 6526 66334 6578 66386
rect 19070 66334 19122 66386
rect 24558 66334 24610 66386
rect 27358 66334 27410 66386
rect 30158 66334 30210 66386
rect 32174 66334 32226 66386
rect 32510 66334 32562 66386
rect 34190 66334 34242 66386
rect 36094 66334 36146 66386
rect 38558 66334 38610 66386
rect 39342 66334 39394 66386
rect 41358 66334 41410 66386
rect 41918 66334 41970 66386
rect 1822 66222 1874 66274
rect 2270 66222 2322 66274
rect 9438 66222 9490 66274
rect 14478 66222 14530 66274
rect 15038 66222 15090 66274
rect 15262 66222 15314 66274
rect 16270 66222 16322 66274
rect 21646 66222 21698 66274
rect 29486 66222 29538 66274
rect 29934 66222 29986 66274
rect 30606 66222 30658 66274
rect 32062 66222 32114 66274
rect 32846 66222 32898 66274
rect 33406 66222 33458 66274
rect 33742 66222 33794 66274
rect 34302 66222 34354 66274
rect 35870 66222 35922 66274
rect 38446 66222 38498 66274
rect 39230 66222 39282 66274
rect 42254 66222 42306 66274
rect 42590 66222 42642 66274
rect 5966 66110 6018 66162
rect 8654 66110 8706 66162
rect 11902 66110 11954 66162
rect 12238 66110 12290 66162
rect 12350 66110 12402 66162
rect 13806 66110 13858 66162
rect 15710 66110 15762 66162
rect 16942 66110 16994 66162
rect 22430 66110 22482 66162
rect 34414 66110 34466 66162
rect 37550 66110 37602 66162
rect 37662 66110 37714 66162
rect 39566 66110 39618 66162
rect 42366 66110 42418 66162
rect 5630 65998 5682 66050
rect 13022 65998 13074 66050
rect 14030 65998 14082 66050
rect 14926 65998 14978 66050
rect 15598 65998 15650 66050
rect 26462 65998 26514 66050
rect 26798 65998 26850 66050
rect 27806 65998 27858 66050
rect 31054 65998 31106 66050
rect 40574 65998 40626 66050
rect 41022 65998 41074 66050
rect 41246 65998 41298 66050
rect 41470 65998 41522 66050
rect 48190 65998 48242 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 1822 65662 1874 65714
rect 13694 65662 13746 65714
rect 14814 65662 14866 65714
rect 15598 65662 15650 65714
rect 38334 65662 38386 65714
rect 39230 65662 39282 65714
rect 39454 65662 39506 65714
rect 5070 65550 5122 65602
rect 7646 65550 7698 65602
rect 7758 65550 7810 65602
rect 12462 65550 12514 65602
rect 13918 65550 13970 65602
rect 14142 65550 14194 65602
rect 15262 65550 15314 65602
rect 16494 65550 16546 65602
rect 18958 65550 19010 65602
rect 20862 65550 20914 65602
rect 20974 65550 21026 65602
rect 24670 65550 24722 65602
rect 32286 65550 32338 65602
rect 34078 65550 34130 65602
rect 35870 65550 35922 65602
rect 38446 65550 38498 65602
rect 39678 65550 39730 65602
rect 40238 65550 40290 65602
rect 41134 65550 41186 65602
rect 41918 65550 41970 65602
rect 4398 65438 4450 65490
rect 8318 65438 8370 65490
rect 11118 65438 11170 65490
rect 11342 65438 11394 65490
rect 11566 65438 11618 65490
rect 11790 65438 11842 65490
rect 12014 65438 12066 65490
rect 12238 65438 12290 65490
rect 12574 65438 12626 65490
rect 13582 65438 13634 65490
rect 14702 65438 14754 65490
rect 15038 65438 15090 65490
rect 15934 65438 15986 65490
rect 20190 65438 20242 65490
rect 20750 65438 20802 65490
rect 21310 65438 21362 65490
rect 22094 65438 22146 65490
rect 30606 65438 30658 65490
rect 32398 65438 32450 65490
rect 33630 65438 33682 65490
rect 36094 65438 36146 65490
rect 36766 65438 36818 65490
rect 37438 65438 37490 65490
rect 37662 65438 37714 65490
rect 38670 65438 38722 65490
rect 40014 65438 40066 65490
rect 40350 65438 40402 65490
rect 42366 65438 42418 65490
rect 7198 65326 7250 65378
rect 8654 65326 8706 65378
rect 10110 65326 10162 65378
rect 10558 65326 10610 65378
rect 10894 65326 10946 65378
rect 16382 65326 16434 65378
rect 18622 65326 18674 65378
rect 19854 65326 19906 65378
rect 24222 65326 24274 65378
rect 30494 65326 30546 65378
rect 33182 65326 33234 65378
rect 36430 65326 36482 65378
rect 39566 65326 39618 65378
rect 41246 65326 41298 65378
rect 42814 65326 42866 65378
rect 7646 65214 7698 65266
rect 8430 65214 8482 65266
rect 8990 65214 9042 65266
rect 13694 65214 13746 65266
rect 14814 65214 14866 65266
rect 16270 65214 16322 65266
rect 18846 65214 18898 65266
rect 20414 65214 20466 65266
rect 24558 65214 24610 65266
rect 30158 65214 30210 65266
rect 32510 65214 32562 65266
rect 40910 65214 40962 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 5966 64878 6018 64930
rect 8430 64878 8482 64930
rect 9326 64878 9378 64930
rect 9886 64878 9938 64930
rect 13918 64878 13970 64930
rect 14254 64878 14306 64930
rect 17838 64878 17890 64930
rect 20414 64878 20466 64930
rect 35758 64878 35810 64930
rect 6190 64766 6242 64818
rect 8878 64766 8930 64818
rect 11342 64766 11394 64818
rect 15934 64766 15986 64818
rect 25342 64766 25394 64818
rect 26126 64766 26178 64818
rect 29822 64766 29874 64818
rect 34414 64766 34466 64818
rect 35422 64766 35474 64818
rect 37550 64766 37602 64818
rect 37886 64766 37938 64818
rect 38222 64766 38274 64818
rect 6526 64654 6578 64706
rect 8990 64654 9042 64706
rect 9550 64654 9602 64706
rect 9886 64654 9938 64706
rect 11118 64654 11170 64706
rect 12014 64654 12066 64706
rect 12350 64654 12402 64706
rect 12910 64654 12962 64706
rect 14254 64654 14306 64706
rect 14926 64654 14978 64706
rect 17614 64654 17666 64706
rect 19070 64654 19122 64706
rect 19294 64654 19346 64706
rect 20414 64654 20466 64706
rect 21310 64654 21362 64706
rect 21646 64654 21698 64706
rect 22094 64654 22146 64706
rect 25902 64654 25954 64706
rect 33742 64654 33794 64706
rect 34638 64654 34690 64706
rect 38558 64654 38610 64706
rect 40014 64654 40066 64706
rect 40686 64654 40738 64706
rect 7982 64542 8034 64594
rect 8318 64542 8370 64594
rect 8766 64542 8818 64594
rect 10222 64542 10274 64594
rect 10782 64542 10834 64594
rect 10894 64542 10946 64594
rect 11566 64542 11618 64594
rect 11790 64542 11842 64594
rect 12574 64542 12626 64594
rect 14590 64542 14642 64594
rect 17278 64542 17330 64594
rect 18174 64542 18226 64594
rect 18398 64542 18450 64594
rect 19518 64542 19570 64594
rect 19742 64542 19794 64594
rect 20078 64542 20130 64594
rect 21870 64542 21922 64594
rect 35198 64542 35250 64594
rect 41246 64542 41298 64594
rect 7198 64430 7250 64482
rect 10558 64430 10610 64482
rect 12238 64430 12290 64482
rect 12798 64430 12850 64482
rect 13694 64430 13746 64482
rect 15486 64430 15538 64482
rect 16942 64430 16994 64482
rect 17614 64430 17666 64482
rect 18958 64430 19010 64482
rect 21758 64430 21810 64482
rect 30270 64430 30322 64482
rect 31166 64430 31218 64482
rect 39678 64430 39730 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 8990 64094 9042 64146
rect 10334 64094 10386 64146
rect 11006 64094 11058 64146
rect 11230 64094 11282 64146
rect 12014 64094 12066 64146
rect 13022 64094 13074 64146
rect 38446 64094 38498 64146
rect 39342 64094 39394 64146
rect 39790 64094 39842 64146
rect 43038 64094 43090 64146
rect 10782 63982 10834 64034
rect 11790 63982 11842 64034
rect 13918 63982 13970 64034
rect 14142 63982 14194 64034
rect 14590 63982 14642 64034
rect 19630 63982 19682 64034
rect 26238 63982 26290 64034
rect 36654 63982 36706 64034
rect 39902 63982 39954 64034
rect 48190 63982 48242 64034
rect 1822 63870 1874 63922
rect 2270 63870 2322 63922
rect 9774 63870 9826 63922
rect 11342 63870 11394 63922
rect 11678 63870 11730 63922
rect 13470 63870 13522 63922
rect 22766 63870 22818 63922
rect 23214 63870 23266 63922
rect 25454 63870 25506 63922
rect 25678 63870 25730 63922
rect 26014 63870 26066 63922
rect 26686 63870 26738 63922
rect 29598 63870 29650 63922
rect 35646 63870 35698 63922
rect 37886 63870 37938 63922
rect 38782 63870 38834 63922
rect 44942 63870 44994 63922
rect 45950 63870 46002 63922
rect 12574 63758 12626 63810
rect 13806 63758 13858 63810
rect 25790 63758 25842 63810
rect 26574 63758 26626 63810
rect 27694 63758 27746 63810
rect 28926 63758 28978 63810
rect 29262 63758 29314 63810
rect 29374 63758 29426 63810
rect 30046 63758 30098 63810
rect 30270 63758 30322 63810
rect 31502 63758 31554 63810
rect 31950 63758 32002 63810
rect 35198 63758 35250 63810
rect 36094 63758 36146 63810
rect 36430 63758 36482 63810
rect 36766 63758 36818 63810
rect 39006 63758 39058 63810
rect 43150 63758 43202 63810
rect 45838 63758 45890 63810
rect 30494 63646 30546 63698
rect 30942 63646 30994 63698
rect 38110 63646 38162 63698
rect 39678 63646 39730 63698
rect 44270 63646 44322 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 17838 63310 17890 63362
rect 18846 63310 18898 63362
rect 19182 63310 19234 63362
rect 19966 63310 20018 63362
rect 27022 63310 27074 63362
rect 31950 63310 32002 63362
rect 32286 63310 32338 63362
rect 34414 63310 34466 63362
rect 35758 63310 35810 63362
rect 42926 63310 42978 63362
rect 1822 63198 1874 63250
rect 6638 63198 6690 63250
rect 17726 63198 17778 63250
rect 20302 63198 20354 63250
rect 25678 63198 25730 63250
rect 29374 63198 29426 63250
rect 34302 63198 34354 63250
rect 42254 63198 42306 63250
rect 43262 63198 43314 63250
rect 44046 63198 44098 63250
rect 46846 63198 46898 63250
rect 17278 63086 17330 63138
rect 17502 63086 17554 63138
rect 18398 63086 18450 63138
rect 18846 63086 18898 63138
rect 26350 63086 26402 63138
rect 26574 63086 26626 63138
rect 27358 63086 27410 63138
rect 27582 63086 27634 63138
rect 31726 63086 31778 63138
rect 34190 63086 34242 63138
rect 35422 63086 35474 63138
rect 43934 63086 43986 63138
rect 45390 63086 45442 63138
rect 45614 63086 45666 63138
rect 46622 63086 46674 63138
rect 14030 62974 14082 63026
rect 14254 62974 14306 63026
rect 14590 62974 14642 63026
rect 18174 62974 18226 63026
rect 25342 62974 25394 63026
rect 29486 62974 29538 63026
rect 31166 62974 31218 63026
rect 35198 62974 35250 63026
rect 6302 62862 6354 62914
rect 16382 62862 16434 62914
rect 16830 62862 16882 62914
rect 19742 62862 19794 62914
rect 20190 62862 20242 62914
rect 28030 62862 28082 62914
rect 28478 62862 28530 62914
rect 31054 62862 31106 62914
rect 42702 62862 42754 62914
rect 42814 62862 42866 62914
rect 45950 62862 46002 62914
rect 46286 62862 46338 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 4622 62526 4674 62578
rect 11118 62526 11170 62578
rect 13134 62526 13186 62578
rect 14702 62526 14754 62578
rect 15262 62526 15314 62578
rect 15598 62526 15650 62578
rect 17502 62526 17554 62578
rect 18174 62526 18226 62578
rect 19406 62526 19458 62578
rect 36766 62526 36818 62578
rect 44046 62526 44098 62578
rect 45278 62526 45330 62578
rect 45726 62526 45778 62578
rect 45950 62526 46002 62578
rect 6414 62414 6466 62466
rect 10670 62414 10722 62466
rect 16270 62414 16322 62466
rect 16606 62414 16658 62466
rect 27022 62414 27074 62466
rect 28030 62414 28082 62466
rect 42478 62414 42530 62466
rect 4958 62302 5010 62354
rect 5854 62302 5906 62354
rect 6302 62302 6354 62354
rect 6638 62302 6690 62354
rect 6974 62302 7026 62354
rect 7758 62302 7810 62354
rect 8430 62302 8482 62354
rect 10446 62302 10498 62354
rect 14926 62302 14978 62354
rect 15934 62302 15986 62354
rect 17278 62302 17330 62354
rect 17614 62302 17666 62354
rect 17950 62302 18002 62354
rect 18286 62302 18338 62354
rect 21870 62302 21922 62354
rect 29150 62302 29202 62354
rect 30270 62302 30322 62354
rect 31390 62302 31442 62354
rect 33182 62302 33234 62354
rect 36990 62302 37042 62354
rect 41582 62302 41634 62354
rect 41694 62302 41746 62354
rect 41806 62302 41858 62354
rect 42254 62302 42306 62354
rect 42926 62302 42978 62354
rect 43710 62302 43762 62354
rect 44046 62302 44098 62354
rect 44270 62302 44322 62354
rect 44942 62302 44994 62354
rect 46286 62302 46338 62354
rect 5742 62190 5794 62242
rect 7310 62190 7362 62242
rect 8990 62190 9042 62242
rect 14254 62190 14306 62242
rect 18846 62190 18898 62242
rect 22542 62190 22594 62242
rect 24670 62190 24722 62242
rect 26686 62190 26738 62242
rect 32174 62190 32226 62242
rect 43374 62190 43426 62242
rect 44718 62190 44770 62242
rect 45838 62190 45890 62242
rect 27246 62078 27298 62130
rect 27582 62078 27634 62130
rect 29374 62078 29426 62130
rect 36654 62078 36706 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 22766 61742 22818 61794
rect 29486 61742 29538 61794
rect 37886 61742 37938 61794
rect 40350 61742 40402 61794
rect 44830 61742 44882 61794
rect 5070 61630 5122 61682
rect 7310 61630 7362 61682
rect 18286 61630 18338 61682
rect 21870 61630 21922 61682
rect 27134 61630 27186 61682
rect 29934 61630 29986 61682
rect 32734 61630 32786 61682
rect 42478 61630 42530 61682
rect 2158 61518 2210 61570
rect 6302 61518 6354 61570
rect 10110 61518 10162 61570
rect 11230 61518 11282 61570
rect 12686 61518 12738 61570
rect 13694 61518 13746 61570
rect 15486 61518 15538 61570
rect 18958 61518 19010 61570
rect 20078 61518 20130 61570
rect 21646 61518 21698 61570
rect 22094 61518 22146 61570
rect 27470 61518 27522 61570
rect 29598 61518 29650 61570
rect 32846 61518 32898 61570
rect 37214 61518 37266 61570
rect 37550 61518 37602 61570
rect 38110 61518 38162 61570
rect 38782 61518 38834 61570
rect 41022 61518 41074 61570
rect 42030 61518 42082 61570
rect 42814 61518 42866 61570
rect 43150 61518 43202 61570
rect 2942 61406 2994 61458
rect 5742 61406 5794 61458
rect 5854 61406 5906 61458
rect 9438 61406 9490 61458
rect 11790 61406 11842 61458
rect 13022 61406 13074 61458
rect 13470 61406 13522 61458
rect 14030 61406 14082 61458
rect 14366 61406 14418 61458
rect 14702 61406 14754 61458
rect 16158 61406 16210 61458
rect 18622 61406 18674 61458
rect 19182 61406 19234 61458
rect 19518 61406 19570 61458
rect 19742 61406 19794 61458
rect 19854 61406 19906 61458
rect 20526 61406 20578 61458
rect 22318 61406 22370 61458
rect 22654 61406 22706 61458
rect 31614 61406 31666 61458
rect 31950 61406 32002 61458
rect 32622 61406 32674 61458
rect 33182 61406 33234 61458
rect 33742 61406 33794 61458
rect 37102 61406 37154 61458
rect 37774 61406 37826 61458
rect 43038 61406 43090 61458
rect 44942 61406 44994 61458
rect 6078 61294 6130 61346
rect 6862 61294 6914 61346
rect 10894 61294 10946 61346
rect 11342 61294 11394 61346
rect 11566 61294 11618 61346
rect 12126 61294 12178 61346
rect 12798 61294 12850 61346
rect 13582 61294 13634 61346
rect 18734 61294 18786 61346
rect 19294 61294 19346 61346
rect 20190 61294 20242 61346
rect 20414 61294 20466 61346
rect 22766 61294 22818 61346
rect 24894 61294 24946 61346
rect 27806 61294 27858 61346
rect 33406 61294 33458 61346
rect 33630 61294 33682 61346
rect 34190 61294 34242 61346
rect 48190 61294 48242 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 4062 60958 4114 61010
rect 8654 60958 8706 61010
rect 14814 60958 14866 61010
rect 18062 60958 18114 61010
rect 29822 60958 29874 61010
rect 31390 60958 31442 61010
rect 31502 60958 31554 61010
rect 32510 60958 32562 61010
rect 33406 60958 33458 61010
rect 37102 60958 37154 61010
rect 37214 60958 37266 61010
rect 38446 60958 38498 61010
rect 41022 60958 41074 61010
rect 41918 60958 41970 61010
rect 4398 60846 4450 60898
rect 6638 60846 6690 60898
rect 12014 60846 12066 60898
rect 15934 60846 15986 60898
rect 16270 60846 16322 60898
rect 25230 60846 25282 60898
rect 31950 60846 32002 60898
rect 34862 60846 34914 60898
rect 35758 60846 35810 60898
rect 36318 60846 36370 60898
rect 36766 60846 36818 60898
rect 40014 60846 40066 60898
rect 41358 60846 41410 60898
rect 1710 60734 1762 60786
rect 5518 60734 5570 60786
rect 6414 60734 6466 60786
rect 6974 60734 7026 60786
rect 7870 60734 7922 60786
rect 8430 60734 8482 60786
rect 9662 60734 9714 60786
rect 11230 60734 11282 60786
rect 15598 60734 15650 60786
rect 16606 60734 16658 60786
rect 16942 60734 16994 60786
rect 17838 60734 17890 60786
rect 18510 60734 18562 60786
rect 21758 60734 21810 60786
rect 25566 60734 25618 60786
rect 29486 60734 29538 60786
rect 32958 60734 33010 60786
rect 33294 60734 33346 60786
rect 33518 60734 33570 60786
rect 33966 60734 34018 60786
rect 34750 60734 34802 60786
rect 34974 60734 35026 60786
rect 35310 60734 35362 60786
rect 35646 60734 35698 60786
rect 35982 60734 36034 60786
rect 36206 60734 36258 60786
rect 36990 60734 37042 60786
rect 37326 60734 37378 60786
rect 38670 60734 38722 60786
rect 39454 60734 39506 60786
rect 40910 60734 40962 60786
rect 41134 60734 41186 60786
rect 2270 60622 2322 60674
rect 5294 60622 5346 60674
rect 5966 60622 6018 60674
rect 14142 60622 14194 60674
rect 15262 60622 15314 60674
rect 16718 60622 16770 60674
rect 19182 60622 19234 60674
rect 21310 60622 21362 60674
rect 22430 60622 22482 60674
rect 24558 60622 24610 60674
rect 28926 60622 28978 60674
rect 29262 60622 29314 60674
rect 32174 60622 32226 60674
rect 33742 60622 33794 60674
rect 34526 60622 34578 60674
rect 41806 60622 41858 60674
rect 6302 60510 6354 60562
rect 31614 60510 31666 60562
rect 34190 60510 34242 60562
rect 34526 60510 34578 60562
rect 36318 60510 36370 60562
rect 42142 60510 42194 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 22766 60174 22818 60226
rect 31614 60174 31666 60226
rect 38222 60174 38274 60226
rect 39790 60174 39842 60226
rect 40126 60174 40178 60226
rect 40686 60174 40738 60226
rect 41022 60174 41074 60226
rect 1822 60062 1874 60114
rect 6750 60062 6802 60114
rect 7870 60062 7922 60114
rect 17614 60062 17666 60114
rect 20078 60062 20130 60114
rect 21870 60062 21922 60114
rect 23326 60062 23378 60114
rect 28590 60062 28642 60114
rect 32510 60062 32562 60114
rect 32846 60062 32898 60114
rect 39566 60062 39618 60114
rect 40462 60062 40514 60114
rect 6414 59950 6466 60002
rect 6862 59950 6914 60002
rect 10670 59950 10722 60002
rect 16942 59950 16994 60002
rect 19854 59950 19906 60002
rect 20190 59950 20242 60002
rect 21646 59950 21698 60002
rect 22094 59950 22146 60002
rect 24670 59950 24722 60002
rect 24894 59950 24946 60002
rect 25342 59950 25394 60002
rect 25678 59950 25730 60002
rect 26462 59950 26514 60002
rect 33182 59950 33234 60002
rect 33406 59950 33458 60002
rect 33630 59950 33682 60002
rect 33854 59950 33906 60002
rect 34862 59950 34914 60002
rect 37438 59950 37490 60002
rect 38334 59950 38386 60002
rect 38894 59950 38946 60002
rect 9998 59838 10050 59890
rect 17166 59838 17218 59890
rect 20526 59838 20578 59890
rect 22318 59838 22370 59890
rect 22654 59838 22706 59890
rect 22766 59838 22818 59890
rect 25118 59838 25170 59890
rect 31726 59838 31778 59890
rect 32174 59838 32226 59890
rect 32958 59838 33010 59890
rect 34190 59838 34242 59890
rect 35198 59838 35250 59890
rect 37662 59838 37714 59890
rect 6190 59726 6242 59778
rect 18286 59726 18338 59778
rect 31278 59726 31330 59778
rect 31614 59726 31666 59778
rect 32398 59726 32450 59778
rect 32622 59726 32674 59778
rect 34078 59726 34130 59778
rect 35982 59726 36034 59778
rect 36318 59726 36370 59778
rect 37102 59726 37154 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 7310 59390 7362 59442
rect 8094 59390 8146 59442
rect 21870 59390 21922 59442
rect 24222 59390 24274 59442
rect 25342 59390 25394 59442
rect 25566 59390 25618 59442
rect 37102 59390 37154 59442
rect 37774 59390 37826 59442
rect 18062 59278 18114 59330
rect 23998 59278 24050 59330
rect 31278 59278 31330 59330
rect 45838 59278 45890 59330
rect 8318 59166 8370 59218
rect 9550 59166 9602 59218
rect 17950 59166 18002 59218
rect 19630 59166 19682 59218
rect 20638 59166 20690 59218
rect 21422 59166 21474 59218
rect 23886 59166 23938 59218
rect 24558 59166 24610 59218
rect 25678 59166 25730 59218
rect 27134 59166 27186 59218
rect 31054 59166 31106 59218
rect 33182 59166 33234 59218
rect 34078 59166 34130 59218
rect 35646 59166 35698 59218
rect 36430 59166 36482 59218
rect 36878 59166 36930 59218
rect 36990 59166 37042 59218
rect 37214 59166 37266 59218
rect 37326 59166 37378 59218
rect 38110 59166 38162 59218
rect 38558 59166 38610 59218
rect 46286 59166 46338 59218
rect 5966 59054 6018 59106
rect 6526 59054 6578 59106
rect 6862 59054 6914 59106
rect 7870 59054 7922 59106
rect 9102 59054 9154 59106
rect 9998 59054 10050 59106
rect 10558 59054 10610 59106
rect 17726 59054 17778 59106
rect 23102 59054 23154 59106
rect 23550 59054 23602 59106
rect 26238 59054 26290 59106
rect 27806 59054 27858 59106
rect 29934 59054 29986 59106
rect 30606 59054 30658 59106
rect 33518 59054 33570 59106
rect 35982 59054 36034 59106
rect 39006 59054 39058 59106
rect 39566 59054 39618 59106
rect 39902 59054 39954 59106
rect 46174 59054 46226 59106
rect 5630 58942 5682 58994
rect 5966 58942 6018 58994
rect 6750 58942 6802 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 17950 58606 18002 58658
rect 22206 58606 22258 58658
rect 22766 58606 22818 58658
rect 26910 58606 26962 58658
rect 31950 58606 32002 58658
rect 6302 58494 6354 58546
rect 16382 58494 16434 58546
rect 17502 58494 17554 58546
rect 17614 58494 17666 58546
rect 18846 58494 18898 58546
rect 22206 58494 22258 58546
rect 29822 58494 29874 58546
rect 31390 58494 31442 58546
rect 43598 58494 43650 58546
rect 44830 58494 44882 58546
rect 45166 58494 45218 58546
rect 6638 58382 6690 58434
rect 6862 58382 6914 58434
rect 7422 58382 7474 58434
rect 8766 58382 8818 58434
rect 9102 58382 9154 58434
rect 13470 58382 13522 58434
rect 18062 58382 18114 58434
rect 24110 58382 24162 58434
rect 24670 58382 24722 58434
rect 25790 58382 25842 58434
rect 26238 58382 26290 58434
rect 26350 58382 26402 58434
rect 30158 58382 30210 58434
rect 30718 58382 30770 58434
rect 31278 58382 31330 58434
rect 39790 58382 39842 58434
rect 43150 58382 43202 58434
rect 43486 58382 43538 58434
rect 45278 58382 45330 58434
rect 46958 58382 47010 58434
rect 1710 58270 1762 58322
rect 2494 58270 2546 58322
rect 5966 58270 6018 58322
rect 6078 58270 6130 58322
rect 6414 58270 6466 58322
rect 8318 58270 8370 58322
rect 8430 58270 8482 58322
rect 9438 58270 9490 58322
rect 9550 58270 9602 58322
rect 14254 58270 14306 58322
rect 18958 58270 19010 58322
rect 2046 58158 2098 58210
rect 5742 58158 5794 58210
rect 7534 58158 7586 58210
rect 8094 58158 8146 58210
rect 8878 58158 8930 58210
rect 9214 58158 9266 58210
rect 9774 58158 9826 58210
rect 9998 58158 10050 58210
rect 10110 58214 10162 58266
rect 19182 58270 19234 58322
rect 23102 58270 23154 58322
rect 24222 58270 24274 58322
rect 24446 58270 24498 58322
rect 27022 58270 27074 58322
rect 29262 58270 29314 58322
rect 37886 58270 37938 58322
rect 38894 58270 38946 58322
rect 40126 58270 40178 58322
rect 43934 58270 43986 58322
rect 46398 58270 46450 58322
rect 46510 58270 46562 58322
rect 48078 58270 48130 58322
rect 10558 58158 10610 58210
rect 11006 58158 11058 58210
rect 11454 58158 11506 58210
rect 18622 58158 18674 58210
rect 22654 58158 22706 58210
rect 23886 58158 23938 58210
rect 25006 58158 25058 58210
rect 25566 58158 25618 58210
rect 26126 58158 26178 58210
rect 26910 58158 26962 58210
rect 28590 58158 28642 58210
rect 39230 58158 39282 58210
rect 40014 58158 40066 58210
rect 40574 58158 40626 58210
rect 41134 58158 41186 58210
rect 44046 58158 44098 58210
rect 44270 58158 44322 58210
rect 46734 58158 46786 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 7646 57822 7698 57874
rect 9662 57822 9714 57874
rect 14366 57822 14418 57874
rect 18174 57822 18226 57874
rect 18734 57822 18786 57874
rect 24446 57822 24498 57874
rect 25566 57822 25618 57874
rect 25790 57822 25842 57874
rect 33742 57822 33794 57874
rect 38894 57822 38946 57874
rect 45614 57822 45666 57874
rect 45838 57822 45890 57874
rect 46174 57822 46226 57874
rect 3166 57710 3218 57762
rect 5854 57710 5906 57762
rect 8766 57710 8818 57762
rect 9886 57710 9938 57762
rect 10558 57710 10610 57762
rect 15822 57710 15874 57762
rect 16718 57710 16770 57762
rect 17502 57710 17554 57762
rect 20638 57710 20690 57762
rect 23774 57710 23826 57762
rect 28366 57710 28418 57762
rect 31278 57710 31330 57762
rect 33966 57710 34018 57762
rect 38334 57710 38386 57762
rect 39118 57710 39170 57762
rect 43486 57710 43538 57762
rect 45166 57710 45218 57762
rect 46846 57710 46898 57762
rect 3502 57598 3554 57650
rect 3950 57598 4002 57650
rect 4622 57598 4674 57650
rect 6414 57598 6466 57650
rect 6750 57598 6802 57650
rect 7086 57598 7138 57650
rect 9438 57598 9490 57650
rect 10110 57598 10162 57650
rect 10894 57598 10946 57650
rect 14142 57598 14194 57650
rect 14590 57598 14642 57650
rect 14702 57598 14754 57650
rect 15486 57598 15538 57650
rect 16494 57598 16546 57650
rect 16830 57598 16882 57650
rect 17614 57598 17666 57650
rect 17950 57598 18002 57650
rect 19966 57598 20018 57650
rect 20190 57598 20242 57650
rect 20526 57598 20578 57650
rect 22206 57598 22258 57650
rect 24558 57598 24610 57650
rect 25454 57598 25506 57650
rect 26014 57598 26066 57650
rect 26238 57598 26290 57650
rect 28142 57598 28194 57650
rect 29710 57598 29762 57650
rect 30158 57598 30210 57650
rect 34078 57598 34130 57650
rect 38670 57598 38722 57650
rect 39230 57598 39282 57650
rect 39678 57598 39730 57650
rect 42926 57598 42978 57650
rect 44494 57598 44546 57650
rect 45502 57598 45554 57650
rect 46062 57598 46114 57650
rect 6078 57486 6130 57538
rect 6638 57486 6690 57538
rect 8094 57486 8146 57538
rect 8766 57486 8818 57538
rect 11678 57486 11730 57538
rect 13806 57486 13858 57538
rect 19406 57486 19458 57538
rect 28926 57486 28978 57538
rect 29598 57486 29650 57538
rect 31054 57486 31106 57538
rect 33518 57486 33570 57538
rect 40126 57486 40178 57538
rect 43038 57486 43090 57538
rect 44270 57486 44322 57538
rect 8542 57374 8594 57426
rect 17502 57374 17554 57426
rect 18286 57374 18338 57426
rect 18622 57374 18674 57426
rect 18958 57374 19010 57426
rect 19182 57374 19234 57426
rect 19518 57374 19570 57426
rect 19854 57374 19906 57426
rect 30718 57374 30770 57426
rect 46174 57374 46226 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 15710 57038 15762 57090
rect 21758 57038 21810 57090
rect 22430 57038 22482 57090
rect 42142 57038 42194 57090
rect 2718 56926 2770 56978
rect 4846 56926 4898 56978
rect 12126 56926 12178 56978
rect 15262 56926 15314 56978
rect 22094 56926 22146 56978
rect 31278 56926 31330 56978
rect 36430 56926 36482 56978
rect 1934 56814 1986 56866
rect 6190 56814 6242 56866
rect 6638 56814 6690 56866
rect 7422 56814 7474 56866
rect 7646 56814 7698 56866
rect 7982 56814 8034 56866
rect 8990 56814 9042 56866
rect 9214 56814 9266 56866
rect 9662 56814 9714 56866
rect 9886 56814 9938 56866
rect 12574 56814 12626 56866
rect 16830 56814 16882 56866
rect 18846 56814 18898 56866
rect 19294 56814 19346 56866
rect 20078 56814 20130 56866
rect 22766 56814 22818 56866
rect 23886 56814 23938 56866
rect 25454 56814 25506 56866
rect 27358 56814 27410 56866
rect 28254 56814 28306 56866
rect 29262 56814 29314 56866
rect 30382 56814 30434 56866
rect 30942 56814 30994 56866
rect 35758 56814 35810 56866
rect 36318 56814 36370 56866
rect 40462 56814 40514 56866
rect 40798 56814 40850 56866
rect 41470 56814 41522 56866
rect 43374 56814 43426 56866
rect 43598 56814 43650 56866
rect 43934 56814 43986 56866
rect 44830 56814 44882 56866
rect 45166 56814 45218 56866
rect 5966 56702 6018 56754
rect 7870 56702 7922 56754
rect 11454 56702 11506 56754
rect 11790 56702 11842 56754
rect 12014 56702 12066 56754
rect 12350 56702 12402 56754
rect 13358 56702 13410 56754
rect 13582 56702 13634 56754
rect 13694 56702 13746 56754
rect 15710 56702 15762 56754
rect 15822 56702 15874 56754
rect 17502 56702 17554 56754
rect 21982 56702 22034 56754
rect 24110 56702 24162 56754
rect 27582 56702 27634 56754
rect 28142 56702 28194 56754
rect 30046 56702 30098 56754
rect 30158 56702 30210 56754
rect 30606 56702 30658 56754
rect 36990 56702 37042 56754
rect 43038 56702 43090 56754
rect 43710 56702 43762 56754
rect 6638 56590 6690 56642
rect 8430 56590 8482 56642
rect 9550 56590 9602 56642
rect 10334 56590 10386 56642
rect 11118 56590 11170 56642
rect 11566 56590 11618 56642
rect 19182 56590 19234 56642
rect 21422 56590 21474 56642
rect 22542 56590 22594 56642
rect 23214 56590 23266 56642
rect 26126 56590 26178 56642
rect 27918 56590 27970 56642
rect 29710 56590 29762 56642
rect 30718 56590 30770 56642
rect 31726 56590 31778 56642
rect 32846 56590 32898 56642
rect 33070 56590 33122 56642
rect 33406 56590 33458 56642
rect 37102 56590 37154 56642
rect 37326 56590 37378 56642
rect 38894 56590 38946 56642
rect 43150 56590 43202 56642
rect 44942 56590 44994 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 7086 56254 7138 56306
rect 10446 56254 10498 56306
rect 14142 56254 14194 56306
rect 16942 56254 16994 56306
rect 18958 56254 19010 56306
rect 24446 56254 24498 56306
rect 25342 56254 25394 56306
rect 28478 56254 28530 56306
rect 34974 56254 35026 56306
rect 37102 56254 37154 56306
rect 41246 56254 41298 56306
rect 2046 56142 2098 56194
rect 7758 56142 7810 56194
rect 11566 56142 11618 56194
rect 12126 56142 12178 56194
rect 13470 56142 13522 56194
rect 13918 56142 13970 56194
rect 17502 56142 17554 56194
rect 20638 56142 20690 56194
rect 24670 56142 24722 56194
rect 25230 56142 25282 56194
rect 26462 56142 26514 56194
rect 28702 56142 28754 56194
rect 33518 56142 33570 56194
rect 36654 56142 36706 56194
rect 37214 56142 37266 56194
rect 41022 56142 41074 56194
rect 42030 56142 42082 56194
rect 1710 56030 1762 56082
rect 10670 56030 10722 56082
rect 11454 56030 11506 56082
rect 11790 56030 11842 56082
rect 13806 56030 13858 56082
rect 17614 56030 17666 56082
rect 20190 56030 20242 56082
rect 20526 56030 20578 56082
rect 22206 56030 22258 56082
rect 24558 56030 24610 56082
rect 25566 56030 25618 56082
rect 27694 56030 27746 56082
rect 29038 56030 29090 56082
rect 34638 56030 34690 56082
rect 36206 56030 36258 56082
rect 37998 56030 38050 56082
rect 40910 56030 40962 56082
rect 47070 56030 47122 56082
rect 2494 55918 2546 55970
rect 5070 55918 5122 55970
rect 6190 55918 6242 55970
rect 6526 55918 6578 55970
rect 9662 55918 9714 55970
rect 18398 55918 18450 55970
rect 19630 55918 19682 55970
rect 26126 55918 26178 55970
rect 30158 55918 30210 55970
rect 30606 55918 30658 55970
rect 33294 55918 33346 55970
rect 35870 55918 35922 55970
rect 38222 55918 38274 55970
rect 38670 55918 38722 55970
rect 41582 55918 41634 55970
rect 46734 55918 46786 55970
rect 48078 55918 48130 55970
rect 8318 55806 8370 55858
rect 17502 55806 17554 55858
rect 18734 55806 18786 55858
rect 19070 55806 19122 55858
rect 37102 55806 37154 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 13582 55470 13634 55522
rect 35758 55470 35810 55522
rect 6078 55358 6130 55410
rect 12910 55358 12962 55410
rect 21534 55358 21586 55410
rect 26014 55358 26066 55410
rect 28030 55358 28082 55410
rect 39342 55358 39394 55410
rect 45614 55358 45666 55410
rect 7758 55246 7810 55298
rect 10110 55246 10162 55298
rect 13694 55246 13746 55298
rect 16046 55246 16098 55298
rect 16942 55246 16994 55298
rect 18622 55246 18674 55298
rect 19294 55246 19346 55298
rect 20078 55246 20130 55298
rect 22318 55246 22370 55298
rect 23102 55246 23154 55298
rect 23550 55246 23602 55298
rect 25454 55246 25506 55298
rect 27358 55246 27410 55298
rect 33294 55246 33346 55298
rect 33518 55246 33570 55298
rect 34414 55246 34466 55298
rect 37998 55246 38050 55298
rect 40798 55246 40850 55298
rect 45838 55246 45890 55298
rect 46846 55246 46898 55298
rect 47070 55246 47122 55298
rect 10782 55134 10834 55186
rect 15934 55134 15986 55186
rect 17502 55134 17554 55186
rect 24110 55134 24162 55186
rect 27582 55134 27634 55186
rect 34190 55134 34242 55186
rect 35870 55134 35922 55186
rect 37438 55134 37490 55186
rect 39118 55134 39170 55186
rect 43934 55134 43986 55186
rect 13582 55022 13634 55074
rect 15710 55022 15762 55074
rect 19182 55022 19234 55074
rect 22766 55022 22818 55074
rect 22990 55022 23042 55074
rect 33854 55022 33906 55074
rect 34750 55022 34802 55074
rect 35758 55022 35810 55074
rect 40574 55022 40626 55074
rect 40686 55022 40738 55074
rect 41022 55022 41074 55074
rect 44046 55022 44098 55074
rect 44158 55022 44210 55074
rect 46174 55022 46226 55074
rect 46510 55022 46562 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 8542 54686 8594 54738
rect 11902 54686 11954 54738
rect 13022 54686 13074 54738
rect 13470 54686 13522 54738
rect 17950 54686 18002 54738
rect 18174 54686 18226 54738
rect 22430 54686 22482 54738
rect 23326 54686 23378 54738
rect 27582 54686 27634 54738
rect 33518 54686 33570 54738
rect 33742 54686 33794 54738
rect 33966 54686 34018 54738
rect 34078 54686 34130 54738
rect 34190 54686 34242 54738
rect 40798 54686 40850 54738
rect 44158 54686 44210 54738
rect 1710 54574 1762 54626
rect 6190 54574 6242 54626
rect 10334 54574 10386 54626
rect 11790 54574 11842 54626
rect 12126 54574 12178 54626
rect 12350 54574 12402 54626
rect 13582 54574 13634 54626
rect 17614 54574 17666 54626
rect 18622 54574 18674 54626
rect 24334 54574 24386 54626
rect 26238 54574 26290 54626
rect 27134 54574 27186 54626
rect 38782 54574 38834 54626
rect 39230 54574 39282 54626
rect 41022 54574 41074 54626
rect 43262 54574 43314 54626
rect 43598 54574 43650 54626
rect 46846 54574 46898 54626
rect 1934 54462 1986 54514
rect 5854 54462 5906 54514
rect 6078 54462 6130 54514
rect 8094 54462 8146 54514
rect 13246 54462 13298 54514
rect 13918 54462 13970 54514
rect 17838 54462 17890 54514
rect 18510 54462 18562 54514
rect 20190 54462 20242 54514
rect 21198 54462 21250 54514
rect 21982 54462 22034 54514
rect 22990 54462 23042 54514
rect 23998 54462 24050 54514
rect 25566 54462 25618 54514
rect 25790 54462 25842 54514
rect 26014 54462 26066 54514
rect 26574 54462 26626 54514
rect 26910 54462 26962 54514
rect 27470 54462 27522 54514
rect 28478 54462 28530 54514
rect 33406 54462 33458 54514
rect 34638 54462 34690 54514
rect 38334 54462 38386 54514
rect 39454 54462 39506 54514
rect 40014 54462 40066 54514
rect 41134 54462 41186 54514
rect 42814 54462 42866 54514
rect 43150 54462 43202 54514
rect 45278 54462 45330 54514
rect 45614 54462 45666 54514
rect 46286 54462 46338 54514
rect 2494 54350 2546 54402
rect 14702 54350 14754 54402
rect 16830 54350 16882 54402
rect 25342 54350 25394 54402
rect 27022 54350 27074 54402
rect 28142 54350 28194 54402
rect 29262 54350 29314 54402
rect 31390 54350 31442 54402
rect 32286 54350 32338 54402
rect 37998 54350 38050 54402
rect 39230 54350 39282 54402
rect 43822 54350 43874 54402
rect 7086 54238 7138 54290
rect 27582 54238 27634 54290
rect 32286 54238 32338 54290
rect 32622 54238 32674 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 18622 53902 18674 53954
rect 33406 53902 33458 53954
rect 38670 53902 38722 53954
rect 41134 53902 41186 53954
rect 4622 53790 4674 53842
rect 15038 53790 15090 53842
rect 32062 53790 32114 53842
rect 38334 53790 38386 53842
rect 40686 53790 40738 53842
rect 44270 53790 44322 53842
rect 45950 53790 46002 53842
rect 1822 53678 1874 53730
rect 11230 53678 11282 53730
rect 14814 53678 14866 53730
rect 15262 53678 15314 53730
rect 21534 53678 21586 53730
rect 23102 53678 23154 53730
rect 24894 53678 24946 53730
rect 25902 53678 25954 53730
rect 26238 53678 26290 53730
rect 26574 53678 26626 53730
rect 27022 53678 27074 53730
rect 29150 53678 29202 53730
rect 29934 53678 29986 53730
rect 33518 53678 33570 53730
rect 38110 53678 38162 53730
rect 41358 53678 41410 53730
rect 41694 53678 41746 53730
rect 41918 53678 41970 53730
rect 42254 53678 42306 53730
rect 42702 53678 42754 53730
rect 43374 53678 43426 53730
rect 43822 53678 43874 53730
rect 46062 53678 46114 53730
rect 46510 53678 46562 53730
rect 46958 53678 47010 53730
rect 2494 53566 2546 53618
rect 6078 53566 6130 53618
rect 6862 53566 6914 53618
rect 10558 53566 10610 53618
rect 15486 53566 15538 53618
rect 16270 53566 16322 53618
rect 18734 53566 18786 53618
rect 21422 53566 21474 53618
rect 24670 53566 24722 53618
rect 27582 53566 27634 53618
rect 27918 53566 27970 53618
rect 32958 53566 33010 53618
rect 42926 53566 42978 53618
rect 45502 53566 45554 53618
rect 48078 53566 48130 53618
rect 5070 53454 5122 53506
rect 8318 53454 8370 53506
rect 16718 53454 16770 53506
rect 18622 53454 18674 53506
rect 25342 53454 25394 53506
rect 26238 53454 26290 53506
rect 28366 53454 28418 53506
rect 32622 53454 32674 53506
rect 33406 53454 33458 53506
rect 33966 53454 34018 53506
rect 41134 53454 41186 53506
rect 41470 53510 41522 53562
rect 42030 53454 42082 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 7534 53118 7586 53170
rect 8878 53118 8930 53170
rect 9774 53118 9826 53170
rect 11566 53118 11618 53170
rect 12014 53118 12066 53170
rect 12574 53118 12626 53170
rect 13806 53118 13858 53170
rect 14254 53118 14306 53170
rect 15598 53118 15650 53170
rect 16382 53118 16434 53170
rect 18286 53118 18338 53170
rect 19294 53118 19346 53170
rect 20750 53118 20802 53170
rect 20974 53118 21026 53170
rect 24782 53118 24834 53170
rect 32510 53118 32562 53170
rect 33966 53118 34018 53170
rect 40462 53118 40514 53170
rect 41918 53118 41970 53170
rect 42478 53118 42530 53170
rect 46734 53118 46786 53170
rect 9102 53006 9154 53058
rect 9550 53006 9602 53058
rect 10110 53006 10162 53058
rect 10558 53006 10610 53058
rect 11230 53006 11282 53058
rect 16270 53006 16322 53058
rect 21870 53006 21922 53058
rect 22654 53006 22706 53058
rect 23214 53006 23266 53058
rect 24446 53006 24498 53058
rect 24558 53006 24610 53058
rect 25678 53006 25730 53058
rect 25790 53006 25842 53058
rect 26014 53006 26066 53058
rect 28142 53006 28194 53058
rect 31390 53006 31442 53058
rect 32286 53006 32338 53058
rect 33742 53006 33794 53058
rect 35870 53006 35922 53058
rect 37438 53006 37490 53058
rect 40238 53006 40290 53058
rect 41246 53006 41298 53058
rect 41806 53006 41858 53058
rect 1710 52894 1762 52946
rect 4958 52894 5010 52946
rect 5966 52894 6018 52946
rect 6190 52894 6242 52946
rect 8766 52894 8818 52946
rect 9886 52894 9938 52946
rect 10334 52894 10386 52946
rect 10670 52894 10722 52946
rect 11902 52894 11954 52946
rect 12238 52894 12290 52946
rect 14142 52894 14194 52946
rect 14478 52894 14530 52946
rect 15262 52894 15314 52946
rect 15710 52894 15762 52946
rect 15822 52894 15874 52946
rect 16606 52894 16658 52946
rect 18510 52894 18562 52946
rect 18958 52894 19010 52946
rect 20638 52894 20690 52946
rect 21982 52894 22034 52946
rect 22430 52894 22482 52946
rect 23550 52894 23602 52946
rect 26910 52894 26962 52946
rect 27470 52894 27522 52946
rect 31054 52894 31106 52946
rect 32174 52894 32226 52946
rect 33630 52894 33682 52946
rect 36318 52894 36370 52946
rect 40126 52894 40178 52946
rect 41022 52894 41074 52946
rect 42142 52894 42194 52946
rect 2494 52782 2546 52834
rect 4622 52782 4674 52834
rect 6750 52782 6802 52834
rect 8094 52782 8146 52834
rect 8430 52782 8482 52834
rect 21422 52782 21474 52834
rect 23998 52782 24050 52834
rect 25454 52782 25506 52834
rect 30270 52782 30322 52834
rect 30718 52782 30770 52834
rect 34302 52782 34354 52834
rect 36766 52782 36818 52834
rect 37550 52782 37602 52834
rect 42926 52782 42978 52834
rect 43374 52782 43426 52834
rect 5406 52670 5458 52722
rect 21870 52670 21922 52722
rect 26238 52670 26290 52722
rect 37214 52670 37266 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 4958 52334 5010 52386
rect 18846 52334 18898 52386
rect 21982 52334 22034 52386
rect 34974 52334 35026 52386
rect 36094 52334 36146 52386
rect 41694 52334 41746 52386
rect 6190 52222 6242 52274
rect 6638 52222 6690 52274
rect 9214 52222 9266 52274
rect 11006 52222 11058 52274
rect 15598 52222 15650 52274
rect 17726 52222 17778 52274
rect 21646 52222 21698 52274
rect 22878 52222 22930 52274
rect 23438 52222 23490 52274
rect 32286 52222 32338 52274
rect 37998 52222 38050 52274
rect 39566 52222 39618 52274
rect 40350 52222 40402 52274
rect 4174 52110 4226 52162
rect 5630 52110 5682 52162
rect 7198 52110 7250 52162
rect 8318 52110 8370 52162
rect 9102 52110 9154 52162
rect 10222 52110 10274 52162
rect 12238 52110 12290 52162
rect 12574 52110 12626 52162
rect 12686 52110 12738 52162
rect 13358 52110 13410 52162
rect 13694 52110 13746 52162
rect 14814 52110 14866 52162
rect 19182 52110 19234 52162
rect 19854 52110 19906 52162
rect 21422 52110 21474 52162
rect 22318 52110 22370 52162
rect 23662 52110 23714 52162
rect 25006 52110 25058 52162
rect 25342 52110 25394 52162
rect 26686 52110 26738 52162
rect 28478 52110 28530 52162
rect 29262 52110 29314 52162
rect 31726 52110 31778 52162
rect 32846 52110 32898 52162
rect 35086 52110 35138 52162
rect 35534 52110 35586 52162
rect 35758 52110 35810 52162
rect 37662 52110 37714 52162
rect 37886 52110 37938 52162
rect 39118 52110 39170 52162
rect 41022 52110 41074 52162
rect 2382 51998 2434 52050
rect 2718 51998 2770 52050
rect 3614 51998 3666 52050
rect 4846 51998 4898 52050
rect 4958 51998 5010 52050
rect 6526 51998 6578 52050
rect 6750 51998 6802 52050
rect 13582 51998 13634 52050
rect 18846 51998 18898 52050
rect 18958 51998 19010 52050
rect 19518 51998 19570 52050
rect 20414 51998 20466 52050
rect 27134 51998 27186 52050
rect 32622 51998 32674 52050
rect 41806 51998 41858 52050
rect 42142 51998 42194 52050
rect 4062 51886 4114 51938
rect 12350 51886 12402 51938
rect 19406 51886 19458 51938
rect 26910 51886 26962 51938
rect 34638 51886 34690 51938
rect 34974 51886 35026 51938
rect 37662 51886 37714 51938
rect 41694 51886 41746 51938
rect 42254 51886 42306 51938
rect 42478 51886 42530 51938
rect 42814 51886 42866 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 9774 51550 9826 51602
rect 20862 51550 20914 51602
rect 22318 51550 22370 51602
rect 22542 51550 22594 51602
rect 22766 51550 22818 51602
rect 23886 51550 23938 51602
rect 24222 51550 24274 51602
rect 35534 51550 35586 51602
rect 38894 51550 38946 51602
rect 40910 51550 40962 51602
rect 46622 51550 46674 51602
rect 4174 51438 4226 51490
rect 7310 51438 7362 51490
rect 11790 51438 11842 51490
rect 20526 51438 20578 51490
rect 20638 51438 20690 51490
rect 41246 51438 41298 51490
rect 43822 51438 43874 51490
rect 44046 51438 44098 51490
rect 4734 51326 4786 51378
rect 5630 51326 5682 51378
rect 6302 51326 6354 51378
rect 8318 51326 8370 51378
rect 8766 51326 8818 51378
rect 11006 51326 11058 51378
rect 22206 51326 22258 51378
rect 25790 51326 25842 51378
rect 26910 51326 26962 51378
rect 28030 51326 28082 51378
rect 28254 51326 28306 51378
rect 29038 51326 29090 51378
rect 30718 51326 30770 51378
rect 35422 51326 35474 51378
rect 39118 51326 39170 51378
rect 42590 51326 42642 51378
rect 46958 51326 47010 51378
rect 2382 51214 2434 51266
rect 3166 51214 3218 51266
rect 8430 51214 8482 51266
rect 10334 51214 10386 51266
rect 13918 51214 13970 51266
rect 18958 51214 19010 51266
rect 23214 51214 23266 51266
rect 28926 51214 28978 51266
rect 30270 51214 30322 51266
rect 33630 51214 33682 51266
rect 36318 51214 36370 51266
rect 41694 51214 41746 51266
rect 42702 51214 42754 51266
rect 43934 51214 43986 51266
rect 48078 51214 48130 51266
rect 8878 51102 8930 51154
rect 26798 51102 26850 51154
rect 28814 51102 28866 51154
rect 35534 51102 35586 51154
rect 42926 51102 42978 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 21310 50766 21362 50818
rect 33294 50766 33346 50818
rect 35982 50766 36034 50818
rect 3726 50654 3778 50706
rect 6526 50654 6578 50706
rect 15374 50654 15426 50706
rect 18174 50654 18226 50706
rect 20078 50654 20130 50706
rect 23438 50654 23490 50706
rect 29822 50654 29874 50706
rect 33966 50654 34018 50706
rect 35310 50654 35362 50706
rect 43038 50654 43090 50706
rect 46062 50654 46114 50706
rect 47630 50654 47682 50706
rect 2494 50542 2546 50594
rect 4510 50542 4562 50594
rect 5630 50542 5682 50594
rect 7534 50542 7586 50594
rect 9774 50542 9826 50594
rect 19070 50542 19122 50594
rect 22206 50542 22258 50594
rect 23662 50542 23714 50594
rect 25006 50542 25058 50594
rect 25342 50542 25394 50594
rect 26686 50542 26738 50594
rect 28366 50542 28418 50594
rect 29374 50542 29426 50594
rect 30270 50542 30322 50594
rect 32510 50542 32562 50594
rect 34302 50542 34354 50594
rect 35758 50542 35810 50594
rect 37886 50542 37938 50594
rect 38334 50542 38386 50594
rect 42814 50542 42866 50594
rect 43486 50542 43538 50594
rect 43934 50542 43986 50594
rect 45950 50542 46002 50594
rect 47406 50542 47458 50594
rect 2158 50430 2210 50482
rect 2830 50430 2882 50482
rect 4286 50430 4338 50482
rect 4958 50430 5010 50482
rect 7646 50430 7698 50482
rect 10222 50430 10274 50482
rect 21422 50430 21474 50482
rect 21646 50430 21698 50482
rect 27134 50430 27186 50482
rect 29038 50430 29090 50482
rect 29262 50430 29314 50482
rect 31054 50430 31106 50482
rect 32734 50430 32786 50482
rect 33294 50430 33346 50482
rect 33406 50430 33458 50482
rect 34750 50430 34802 50482
rect 43150 50430 43202 50482
rect 44270 50430 44322 50482
rect 1934 50318 1986 50370
rect 2046 50318 2098 50370
rect 11118 50318 11170 50370
rect 18622 50318 18674 50370
rect 20750 50318 20802 50370
rect 28590 50318 28642 50370
rect 31390 50318 31442 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 2606 49982 2658 50034
rect 3838 49982 3890 50034
rect 7870 49982 7922 50034
rect 12238 49982 12290 50034
rect 13470 49982 13522 50034
rect 15822 49982 15874 50034
rect 6862 49870 6914 49922
rect 8542 49870 8594 49922
rect 11006 49870 11058 49922
rect 12350 49870 12402 49922
rect 16270 49870 16322 49922
rect 16382 49926 16434 49978
rect 17838 49982 17890 50034
rect 17950 49982 18002 50034
rect 18510 49982 18562 50034
rect 18846 49982 18898 50034
rect 19406 49982 19458 50034
rect 25566 49982 25618 50034
rect 26238 49982 26290 50034
rect 19630 49870 19682 49922
rect 21870 49870 21922 49922
rect 25230 49870 25282 49922
rect 25902 49870 25954 49922
rect 26014 49870 26066 49922
rect 26574 49870 26626 49922
rect 33182 49926 33234 49978
rect 35758 49982 35810 50034
rect 39902 49982 39954 50034
rect 41582 49982 41634 50034
rect 33406 49870 33458 49922
rect 34302 49870 34354 49922
rect 35982 49870 36034 49922
rect 39566 49870 39618 49922
rect 40910 49870 40962 49922
rect 41022 49870 41074 49922
rect 47742 49870 47794 49922
rect 2158 49758 2210 49810
rect 2382 49758 2434 49810
rect 2606 49758 2658 49810
rect 2942 49758 2994 49810
rect 6638 49758 6690 49810
rect 7758 49758 7810 49810
rect 11118 49758 11170 49810
rect 13806 49758 13858 49810
rect 15150 49758 15202 49810
rect 15598 49758 15650 49810
rect 19182 49758 19234 49810
rect 19742 49758 19794 49810
rect 20750 49758 20802 49810
rect 21198 49758 21250 49810
rect 22206 49758 22258 49810
rect 23438 49758 23490 49810
rect 26462 49758 26514 49810
rect 26798 49758 26850 49810
rect 27134 49758 27186 49810
rect 27806 49758 27858 49810
rect 31614 49758 31666 49810
rect 33070 49758 33122 49810
rect 33742 49758 33794 49810
rect 34526 49758 34578 49810
rect 36094 49758 36146 49810
rect 40126 49758 40178 49810
rect 43262 49758 43314 49810
rect 43710 49758 43762 49810
rect 46174 49758 46226 49810
rect 47518 49758 47570 49810
rect 1934 49646 1986 49698
rect 3390 49646 3442 49698
rect 4510 49646 4562 49698
rect 4958 49646 5010 49698
rect 5518 49646 5570 49698
rect 10558 49646 10610 49698
rect 14254 49646 14306 49698
rect 14814 49646 14866 49698
rect 20302 49646 20354 49698
rect 23774 49646 23826 49698
rect 24670 49646 24722 49698
rect 28590 49646 28642 49698
rect 30718 49646 30770 49698
rect 31390 49646 31442 49698
rect 36542 49646 36594 49698
rect 44158 49646 44210 49698
rect 45950 49646 46002 49698
rect 11006 49534 11058 49586
rect 12238 49534 12290 49586
rect 14814 49534 14866 49586
rect 15150 49534 15202 49586
rect 16270 49534 16322 49586
rect 18062 49534 18114 49586
rect 31950 49534 32002 49586
rect 34862 49534 34914 49586
rect 41022 49534 41074 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 46062 49198 46114 49250
rect 12686 49086 12738 49138
rect 18398 49086 18450 49138
rect 21758 49086 21810 49138
rect 22654 49086 22706 49138
rect 32062 49086 32114 49138
rect 35870 49086 35922 49138
rect 38894 49086 38946 49138
rect 40462 49086 40514 49138
rect 40798 49086 40850 49138
rect 44270 49086 44322 49138
rect 46398 49086 46450 49138
rect 1710 48974 1762 49026
rect 7198 48974 7250 49026
rect 7646 48974 7698 49026
rect 8990 48974 9042 49026
rect 9886 48974 9938 49026
rect 10558 48974 10610 49026
rect 13582 48974 13634 49026
rect 14142 48974 14194 49026
rect 15038 48974 15090 49026
rect 15710 48974 15762 49026
rect 16158 48974 16210 49026
rect 17054 48974 17106 49026
rect 17726 48974 17778 49026
rect 18622 48974 18674 49026
rect 19070 48974 19122 49026
rect 20750 48974 20802 49026
rect 21422 48974 21474 49026
rect 22206 48974 22258 49026
rect 23326 48974 23378 49026
rect 25230 48974 25282 49026
rect 26910 48974 26962 49026
rect 29150 48974 29202 49026
rect 35086 48974 35138 49026
rect 36094 48974 36146 49026
rect 39230 48974 39282 49026
rect 40014 48974 40066 49026
rect 43822 48974 43874 49026
rect 44158 48974 44210 49026
rect 46174 48974 46226 49026
rect 46958 48974 47010 49026
rect 2494 48862 2546 48914
rect 7534 48862 7586 48914
rect 13806 48862 13858 48914
rect 14478 48862 14530 48914
rect 14702 48862 14754 48914
rect 15262 48862 15314 48914
rect 19518 48862 19570 48914
rect 23214 48862 23266 48914
rect 27358 48862 27410 48914
rect 29934 48862 29986 48914
rect 32398 48862 32450 48914
rect 32958 48862 33010 48914
rect 33630 48862 33682 48914
rect 35534 48862 35586 48914
rect 35646 48862 35698 48914
rect 37998 48862 38050 48914
rect 39566 48862 39618 48914
rect 40126 48862 40178 48914
rect 40910 48862 40962 48914
rect 41582 48862 41634 48914
rect 4734 48750 4786 48802
rect 14254 48750 14306 48802
rect 14814 48750 14866 48802
rect 20190 48750 20242 48802
rect 25790 48750 25842 48802
rect 27806 48750 27858 48802
rect 33294 48750 33346 48802
rect 34862 48750 34914 48802
rect 35310 48750 35362 48802
rect 36430 48750 36482 48802
rect 37662 48750 37714 48802
rect 37886 48750 37938 48802
rect 40350 48750 40402 48802
rect 40462 48750 40514 48802
rect 41134 48750 41186 48802
rect 41358 48750 41410 48802
rect 47742 48750 47794 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 2494 48414 2546 48466
rect 4846 48414 4898 48466
rect 6078 48414 6130 48466
rect 8990 48414 9042 48466
rect 9550 48414 9602 48466
rect 10782 48414 10834 48466
rect 12238 48414 12290 48466
rect 24334 48414 24386 48466
rect 25342 48414 25394 48466
rect 28478 48414 28530 48466
rect 31838 48414 31890 48466
rect 34414 48414 34466 48466
rect 41022 48414 41074 48466
rect 41246 48414 41298 48466
rect 46174 48414 46226 48466
rect 46734 48414 46786 48466
rect 47182 48414 47234 48466
rect 2158 48302 2210 48354
rect 3614 48302 3666 48354
rect 4398 48302 4450 48354
rect 6414 48302 6466 48354
rect 11006 48302 11058 48354
rect 12574 48302 12626 48354
rect 14142 48302 14194 48354
rect 17838 48302 17890 48354
rect 17950 48302 18002 48354
rect 26462 48302 26514 48354
rect 37886 48302 37938 48354
rect 38222 48302 38274 48354
rect 43038 48302 43090 48354
rect 44382 48302 44434 48354
rect 44494 48302 44546 48354
rect 47406 48302 47458 48354
rect 47742 48302 47794 48354
rect 2494 48190 2546 48242
rect 2718 48190 2770 48242
rect 3390 48190 3442 48242
rect 4286 48190 4338 48242
rect 6638 48190 6690 48242
rect 8206 48190 8258 48242
rect 10670 48190 10722 48242
rect 11230 48190 11282 48242
rect 13470 48190 13522 48242
rect 23662 48190 23714 48242
rect 23998 48190 24050 48242
rect 24334 48190 24386 48242
rect 24558 48190 24610 48242
rect 25230 48190 25282 48242
rect 25454 48190 25506 48242
rect 25790 48190 25842 48242
rect 26798 48190 26850 48242
rect 28254 48190 28306 48242
rect 28590 48190 28642 48242
rect 31502 48190 31554 48242
rect 34526 48190 34578 48242
rect 35198 48190 35250 48242
rect 37214 48190 37266 48242
rect 38670 48190 38722 48242
rect 39566 48190 39618 48242
rect 40910 48190 40962 48242
rect 42590 48190 42642 48242
rect 42814 48190 42866 48242
rect 44718 48190 44770 48242
rect 9998 48078 10050 48130
rect 11342 48078 11394 48130
rect 11678 48078 11730 48130
rect 16270 48078 16322 48130
rect 18622 48078 18674 48130
rect 34974 48078 35026 48130
rect 35870 48078 35922 48130
rect 37102 48078 37154 48130
rect 38558 48078 38610 48130
rect 40126 48078 40178 48130
rect 2606 47966 2658 48018
rect 42702 48078 42754 48130
rect 45390 48078 45442 48130
rect 45614 48078 45666 48130
rect 11678 47966 11730 48018
rect 18062 47966 18114 48018
rect 34414 47966 34466 48018
rect 45838 47966 45890 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 2158 47630 2210 47682
rect 2494 47630 2546 47682
rect 20302 47630 20354 47682
rect 32958 47630 33010 47682
rect 43486 47630 43538 47682
rect 3838 47518 3890 47570
rect 19742 47518 19794 47570
rect 23774 47518 23826 47570
rect 25678 47518 25730 47570
rect 26574 47518 26626 47570
rect 33630 47518 33682 47570
rect 34414 47518 34466 47570
rect 41918 47518 41970 47570
rect 2494 47406 2546 47458
rect 2942 47406 2994 47458
rect 4846 47406 4898 47458
rect 7646 47406 7698 47458
rect 10558 47406 10610 47458
rect 11006 47406 11058 47458
rect 14590 47406 14642 47458
rect 15150 47406 15202 47458
rect 20414 47406 20466 47458
rect 21310 47406 21362 47458
rect 4174 47294 4226 47346
rect 4398 47294 4450 47346
rect 22990 47350 23042 47402
rect 24334 47406 24386 47458
rect 24670 47406 24722 47458
rect 25342 47406 25394 47458
rect 33854 47406 33906 47458
rect 34750 47406 34802 47458
rect 34974 47406 35026 47458
rect 37214 47406 37266 47458
rect 37438 47406 37490 47458
rect 40238 47406 40290 47458
rect 41806 47406 41858 47458
rect 42814 47406 42866 47458
rect 4958 47294 5010 47346
rect 7982 47294 8034 47346
rect 14366 47294 14418 47346
rect 15374 47294 15426 47346
rect 22430 47294 22482 47346
rect 23102 47294 23154 47346
rect 25006 47294 25058 47346
rect 25118 47294 25170 47346
rect 32958 47294 33010 47346
rect 33070 47294 33122 47346
rect 37662 47294 37714 47346
rect 39902 47294 39954 47346
rect 40014 47294 40066 47346
rect 40462 47294 40514 47346
rect 4286 47182 4338 47234
rect 5182 47182 5234 47234
rect 7646 47182 7698 47234
rect 20302 47182 20354 47234
rect 23326 47182 23378 47234
rect 24222 47182 24274 47234
rect 24558 47182 24610 47234
rect 26126 47182 26178 47234
rect 34862 47182 34914 47234
rect 35198 47182 35250 47234
rect 37326 47182 37378 47234
rect 38446 47182 38498 47234
rect 38782 47182 38834 47234
rect 39678 47182 39730 47234
rect 40574 47182 40626 47234
rect 40798 47182 40850 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 7534 46846 7586 46898
rect 8318 46846 8370 46898
rect 9886 46846 9938 46898
rect 11678 46846 11730 46898
rect 13470 46846 13522 46898
rect 14142 46846 14194 46898
rect 17502 46846 17554 46898
rect 18062 46846 18114 46898
rect 20638 46846 20690 46898
rect 23326 46846 23378 46898
rect 23886 46846 23938 46898
rect 26238 46846 26290 46898
rect 34974 46846 35026 46898
rect 35086 46846 35138 46898
rect 42590 46846 42642 46898
rect 46622 46846 46674 46898
rect 3502 46734 3554 46786
rect 5406 46734 5458 46786
rect 5742 46734 5794 46786
rect 6078 46734 6130 46786
rect 8878 46734 8930 46786
rect 9550 46734 9602 46786
rect 10558 46734 10610 46786
rect 11230 46734 11282 46786
rect 13806 46734 13858 46786
rect 22990 46734 23042 46786
rect 23102 46734 23154 46786
rect 24222 46734 24274 46786
rect 24334 46734 24386 46786
rect 30718 46734 30770 46786
rect 33742 46734 33794 46786
rect 33854 46734 33906 46786
rect 44494 46734 44546 46786
rect 3838 46622 3890 46674
rect 4846 46622 4898 46674
rect 10222 46622 10274 46674
rect 17390 46622 17442 46674
rect 18286 46622 18338 46674
rect 20750 46622 20802 46674
rect 23550 46622 23602 46674
rect 24558 46622 24610 46674
rect 25118 46622 25170 46674
rect 25566 46622 25618 46674
rect 25678 46622 25730 46674
rect 26126 46622 26178 46674
rect 26798 46622 26850 46674
rect 34414 46622 34466 46674
rect 34750 46622 34802 46674
rect 42254 46622 42306 46674
rect 43822 46622 43874 46674
rect 46958 46622 47010 46674
rect 7982 46510 8034 46562
rect 18958 46510 19010 46562
rect 21198 46510 21250 46562
rect 22206 46510 22258 46562
rect 22654 46510 22706 46562
rect 25342 46510 25394 46562
rect 27470 46510 27522 46562
rect 29598 46510 29650 46562
rect 31278 46510 31330 46562
rect 38110 46510 38162 46562
rect 40126 46510 40178 46562
rect 42030 46510 42082 46562
rect 44046 46510 44098 46562
rect 48078 46510 48130 46562
rect 11230 46398 11282 46450
rect 11678 46398 11730 46450
rect 17502 46398 17554 46450
rect 26238 46398 26290 46450
rect 30606 46398 30658 46450
rect 33742 46398 33794 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 17502 46062 17554 46114
rect 18510 46062 18562 46114
rect 42478 46062 42530 46114
rect 42814 46062 42866 46114
rect 6414 45950 6466 46002
rect 8542 45950 8594 46002
rect 11566 45950 11618 46002
rect 13582 45950 13634 46002
rect 17166 45950 17218 46002
rect 24894 45950 24946 46002
rect 39902 45950 39954 46002
rect 43710 45950 43762 46002
rect 45166 45950 45218 46002
rect 4398 45838 4450 45890
rect 4734 45838 4786 45890
rect 4958 45838 5010 45890
rect 5742 45838 5794 45890
rect 14142 45838 14194 45890
rect 14814 45838 14866 45890
rect 15374 45838 15426 45890
rect 15822 45838 15874 45890
rect 15934 45838 15986 45890
rect 16606 45838 16658 45890
rect 17838 45838 17890 45890
rect 18622 45838 18674 45890
rect 18958 45838 19010 45890
rect 20638 45838 20690 45890
rect 22318 45838 22370 45890
rect 22878 45838 22930 45890
rect 23886 45838 23938 45890
rect 24446 45838 24498 45890
rect 26910 45838 26962 45890
rect 31390 45838 31442 45890
rect 40798 45838 40850 45890
rect 42254 45838 42306 45890
rect 44046 45838 44098 45890
rect 9550 45726 9602 45778
rect 9886 45726 9938 45778
rect 10222 45726 10274 45778
rect 10558 45726 10610 45778
rect 11006 45726 11058 45778
rect 11230 45726 11282 45778
rect 11678 45726 11730 45778
rect 11902 45726 11954 45778
rect 14478 45726 14530 45778
rect 18062 45726 18114 45778
rect 20750 45726 20802 45778
rect 21534 45726 21586 45778
rect 21870 45726 21922 45778
rect 23214 45726 23266 45778
rect 23438 45726 23490 45778
rect 26238 45726 26290 45778
rect 26574 45726 26626 45778
rect 30270 45726 30322 45778
rect 30830 45726 30882 45778
rect 31054 45726 31106 45778
rect 31502 45726 31554 45778
rect 32062 45726 32114 45778
rect 40462 45726 40514 45778
rect 40574 45726 40626 45778
rect 44158 45726 44210 45778
rect 45614 45726 45666 45778
rect 46958 45726 47010 45778
rect 4846 45614 4898 45666
rect 9326 45614 9378 45666
rect 11118 45614 11170 45666
rect 12350 45614 12402 45666
rect 15150 45614 15202 45666
rect 15598 45614 15650 45666
rect 16382 45614 16434 45666
rect 19630 45614 19682 45666
rect 20190 45614 20242 45666
rect 21982 45614 22034 45666
rect 23326 45614 23378 45666
rect 29598 45614 29650 45666
rect 29934 45614 29986 45666
rect 30942 45614 30994 45666
rect 41246 45614 41298 45666
rect 44382 45614 44434 45666
rect 46846 45614 46898 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 1934 45278 1986 45330
rect 2158 45278 2210 45330
rect 14590 45278 14642 45330
rect 15262 45278 15314 45330
rect 15374 45278 15426 45330
rect 15598 45278 15650 45330
rect 18622 45278 18674 45330
rect 29934 45278 29986 45330
rect 41022 45278 41074 45330
rect 41470 45278 41522 45330
rect 3166 45166 3218 45218
rect 12238 45166 12290 45218
rect 13694 45166 13746 45218
rect 18958 45166 19010 45218
rect 20414 45166 20466 45218
rect 20750 45166 20802 45218
rect 23662 45166 23714 45218
rect 25902 45166 25954 45218
rect 27134 45166 27186 45218
rect 32062 45166 32114 45218
rect 35198 45166 35250 45218
rect 35646 45166 35698 45218
rect 35870 45166 35922 45218
rect 36206 45166 36258 45218
rect 36318 45166 36370 45218
rect 36766 45166 36818 45218
rect 38334 45166 38386 45218
rect 39902 45166 39954 45218
rect 2494 45054 2546 45106
rect 2830 45054 2882 45106
rect 7870 45054 7922 45106
rect 8318 45054 8370 45106
rect 13022 45054 13074 45106
rect 13358 45054 13410 45106
rect 15710 45054 15762 45106
rect 17502 45054 17554 45106
rect 17838 45054 17890 45106
rect 21198 45054 21250 45106
rect 23326 45054 23378 45106
rect 25230 45054 25282 45106
rect 25790 45054 25842 45106
rect 26014 45054 26066 45106
rect 26350 45054 26402 45106
rect 29822 45054 29874 45106
rect 30158 45054 30210 45106
rect 30830 45054 30882 45106
rect 31838 45054 31890 45106
rect 34750 45054 34802 45106
rect 35534 45054 35586 45106
rect 36542 45054 36594 45106
rect 36878 45110 36930 45162
rect 40238 45166 40290 45218
rect 42030 45166 42082 45218
rect 44718 45166 44770 45218
rect 44830 45166 44882 45218
rect 38670 45054 38722 45106
rect 41358 45054 41410 45106
rect 45054 45054 45106 45106
rect 3614 44942 3666 44994
rect 7534 44942 7586 44994
rect 8990 44942 9042 44994
rect 9662 44942 9714 44994
rect 10110 44942 10162 44994
rect 14142 44942 14194 44994
rect 17726 44942 17778 44994
rect 19182 44942 19234 44994
rect 19630 44942 19682 44994
rect 2830 44830 2882 44882
rect 13358 44830 13410 44882
rect 21758 44942 21810 44994
rect 22206 44942 22258 44994
rect 24670 44942 24722 44994
rect 29262 44942 29314 44994
rect 30718 44942 30770 44994
rect 31950 44942 32002 44994
rect 34302 44942 34354 44994
rect 37998 44942 38050 44994
rect 39566 44942 39618 44994
rect 45726 44942 45778 44994
rect 19518 44830 19570 44882
rect 19854 44830 19906 44882
rect 20190 44830 20242 44882
rect 24446 44830 24498 44882
rect 24670 44830 24722 44882
rect 25454 44830 25506 44882
rect 31054 44830 31106 44882
rect 36206 44830 36258 44882
rect 41470 44830 41522 44882
rect 45838 44830 45890 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 2718 44494 2770 44546
rect 13694 44494 13746 44546
rect 20078 44494 20130 44546
rect 23102 44494 23154 44546
rect 25118 44494 25170 44546
rect 43262 44494 43314 44546
rect 46622 44494 46674 44546
rect 5742 44382 5794 44434
rect 6302 44382 6354 44434
rect 14030 44382 14082 44434
rect 15934 44382 15986 44434
rect 18062 44382 18114 44434
rect 20414 44382 20466 44434
rect 23550 44382 23602 44434
rect 24670 44382 24722 44434
rect 31502 44382 31554 44434
rect 32398 44382 32450 44434
rect 34078 44382 34130 44434
rect 42702 44382 42754 44434
rect 45950 44382 46002 44434
rect 2158 44270 2210 44322
rect 2942 44270 2994 44322
rect 12910 44270 12962 44322
rect 14590 44270 14642 44322
rect 16382 44270 16434 44322
rect 16830 44270 16882 44322
rect 17838 44270 17890 44322
rect 22094 44270 22146 44322
rect 23886 44270 23938 44322
rect 24894 44270 24946 44322
rect 25342 44270 25394 44322
rect 30046 44270 30098 44322
rect 30718 44270 30770 44322
rect 30942 44270 30994 44322
rect 31838 44270 31890 44322
rect 34414 44270 34466 44322
rect 34974 44270 35026 44322
rect 37102 44270 37154 44322
rect 37326 44270 37378 44322
rect 37998 44270 38050 44322
rect 38446 44270 38498 44322
rect 38670 44270 38722 44322
rect 39678 44270 39730 44322
rect 42590 44270 42642 44322
rect 47070 44270 47122 44322
rect 2382 44158 2434 44210
rect 3278 44158 3330 44210
rect 3950 44158 4002 44210
rect 4174 44158 4226 44210
rect 6526 44158 6578 44210
rect 7198 44158 7250 44210
rect 7870 44158 7922 44210
rect 13918 44158 13970 44210
rect 14366 44158 14418 44210
rect 16270 44158 16322 44210
rect 17054 44158 17106 44210
rect 22430 44158 22482 44210
rect 22766 44158 22818 44210
rect 23998 44158 24050 44210
rect 25678 44158 25730 44210
rect 29710 44158 29762 44210
rect 31054 44158 31106 44210
rect 39342 44158 39394 44210
rect 40014 44158 40066 44210
rect 40686 44158 40738 44210
rect 41022 44158 41074 44210
rect 41134 44158 41186 44210
rect 41582 44158 41634 44210
rect 41694 44158 41746 44210
rect 46286 44158 46338 44210
rect 46510 44158 46562 44210
rect 2494 44046 2546 44098
rect 3614 44046 3666 44098
rect 4062 44046 4114 44098
rect 4734 44046 4786 44098
rect 6638 44046 6690 44098
rect 6862 44046 6914 44098
rect 7086 44046 7138 44098
rect 15262 44046 15314 44098
rect 16046 44046 16098 44098
rect 17502 44046 17554 44098
rect 20302 44046 20354 44098
rect 21758 44046 21810 44098
rect 22990 44046 23042 44098
rect 24222 44046 24274 44098
rect 25566 44046 25618 44098
rect 26238 44046 26290 44098
rect 29374 44046 29426 44098
rect 29822 44046 29874 44098
rect 40350 44046 40402 44098
rect 41358 44046 41410 44098
rect 41918 44046 41970 44098
rect 47742 44046 47794 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 3726 43710 3778 43762
rect 10894 43710 10946 43762
rect 12462 43710 12514 43762
rect 14478 43710 14530 43762
rect 18286 43710 18338 43762
rect 19518 43710 19570 43762
rect 20302 43710 20354 43762
rect 39342 43710 39394 43762
rect 39902 43710 39954 43762
rect 41022 43710 41074 43762
rect 2158 43598 2210 43650
rect 5294 43598 5346 43650
rect 5406 43598 5458 43650
rect 5854 43598 5906 43650
rect 6638 43598 6690 43650
rect 6862 43598 6914 43650
rect 8878 43598 8930 43650
rect 10222 43598 10274 43650
rect 11454 43598 11506 43650
rect 15374 43598 15426 43650
rect 15598 43598 15650 43650
rect 16382 43598 16434 43650
rect 16606 43598 16658 43650
rect 16718 43598 16770 43650
rect 18510 43598 18562 43650
rect 20190 43598 20242 43650
rect 20862 43598 20914 43650
rect 22094 43598 22146 43650
rect 23774 43598 23826 43650
rect 23998 43598 24050 43650
rect 24110 43598 24162 43650
rect 42478 43598 42530 43650
rect 42814 43598 42866 43650
rect 2382 43486 2434 43538
rect 2606 43486 2658 43538
rect 2942 43486 2994 43538
rect 4510 43486 4562 43538
rect 4622 43486 4674 43538
rect 4958 43486 5010 43538
rect 5630 43486 5682 43538
rect 6190 43486 6242 43538
rect 7086 43486 7138 43538
rect 7646 43486 7698 43538
rect 9550 43486 9602 43538
rect 9886 43486 9938 43538
rect 10558 43486 10610 43538
rect 11006 43486 11058 43538
rect 11230 43486 11282 43538
rect 11678 43486 11730 43538
rect 12014 43486 12066 43538
rect 12350 43486 12402 43538
rect 12574 43486 12626 43538
rect 12798 43486 12850 43538
rect 13694 43486 13746 43538
rect 14030 43486 14082 43538
rect 14142 43486 14194 43538
rect 14254 43486 14306 43538
rect 15934 43486 15986 43538
rect 16270 43486 16322 43538
rect 18622 43486 18674 43538
rect 19854 43486 19906 43538
rect 21310 43486 21362 43538
rect 21870 43486 21922 43538
rect 24334 43486 24386 43538
rect 25230 43486 25282 43538
rect 25566 43486 25618 43538
rect 25790 43486 25842 43538
rect 26462 43486 26514 43538
rect 37886 43486 37938 43538
rect 38110 43486 38162 43538
rect 40126 43486 40178 43538
rect 41582 43486 41634 43538
rect 42030 43486 42082 43538
rect 43038 43486 43090 43538
rect 45950 43486 46002 43538
rect 46510 43486 46562 43538
rect 46622 43486 46674 43538
rect 46846 43486 46898 43538
rect 47182 43486 47234 43538
rect 47406 43486 47458 43538
rect 2270 43374 2322 43426
rect 4846 43374 4898 43426
rect 6750 43374 6802 43426
rect 7534 43374 7586 43426
rect 8542 43374 8594 43426
rect 13246 43374 13298 43426
rect 16046 43374 16098 43426
rect 18174 43374 18226 43426
rect 18958 43374 19010 43426
rect 25342 43374 25394 43426
rect 27246 43374 27298 43426
rect 29374 43374 29426 43426
rect 45278 43374 45330 43426
rect 47070 43374 47122 43426
rect 9886 43262 9938 43314
rect 19182 43262 19234 43314
rect 38446 43262 38498 43314
rect 43374 43262 43426 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 6638 42926 6690 42978
rect 7086 42926 7138 42978
rect 8654 42926 8706 42978
rect 9886 42926 9938 42978
rect 11006 42926 11058 42978
rect 12574 42926 12626 42978
rect 13022 42926 13074 42978
rect 27022 42926 27074 42978
rect 33070 42926 33122 42978
rect 42590 42926 42642 42978
rect 8766 42814 8818 42866
rect 12798 42814 12850 42866
rect 15038 42814 15090 42866
rect 16382 42814 16434 42866
rect 34414 42814 34466 42866
rect 37550 42814 37602 42866
rect 38110 42814 38162 42866
rect 41246 42814 41298 42866
rect 41918 42814 41970 42866
rect 43038 42814 43090 42866
rect 46398 42814 46450 42866
rect 46846 42814 46898 42866
rect 3726 42702 3778 42754
rect 4398 42702 4450 42754
rect 5630 42702 5682 42754
rect 7310 42702 7362 42754
rect 9550 42702 9602 42754
rect 10334 42702 10386 42754
rect 10894 42702 10946 42754
rect 11230 42702 11282 42754
rect 11454 42702 11506 42754
rect 13806 42702 13858 42754
rect 20414 42702 20466 42754
rect 22430 42702 22482 42754
rect 24110 42702 24162 42754
rect 26238 42702 26290 42754
rect 26910 42702 26962 42754
rect 27694 42702 27746 42754
rect 33294 42702 33346 42754
rect 37438 42702 37490 42754
rect 38446 42702 38498 42754
rect 43262 42702 43314 42754
rect 46174 42702 46226 42754
rect 3166 42590 3218 42642
rect 6526 42590 6578 42642
rect 6974 42590 7026 42642
rect 7758 42590 7810 42642
rect 9102 42590 9154 42642
rect 10110 42590 10162 42642
rect 13470 42590 13522 42642
rect 20078 42590 20130 42642
rect 20302 42590 20354 42642
rect 23214 42590 23266 42642
rect 25678 42590 25730 42642
rect 27022 42590 27074 42642
rect 33966 42590 34018 42642
rect 37214 42590 37266 42642
rect 42702 42590 42754 42642
rect 4958 42478 5010 42530
rect 5742 42478 5794 42530
rect 5854 42478 5906 42530
rect 9550 42478 9602 42530
rect 11342 42478 11394 42530
rect 11902 42478 11954 42530
rect 12350 42478 12402 42530
rect 19742 42478 19794 42530
rect 21422 42478 21474 42530
rect 22094 42478 22146 42530
rect 25006 42478 25058 42530
rect 28030 42478 28082 42530
rect 32734 42478 32786 42530
rect 36318 42478 36370 42530
rect 39006 42478 39058 42530
rect 40686 42478 40738 42530
rect 42254 42478 42306 42530
rect 42478 42478 42530 42530
rect 43598 42478 43650 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 10222 42142 10274 42194
rect 10894 42142 10946 42194
rect 16494 42142 16546 42194
rect 20638 42142 20690 42194
rect 20974 42142 21026 42194
rect 33294 42142 33346 42194
rect 36654 42142 36706 42194
rect 4734 42030 4786 42082
rect 16382 42030 16434 42082
rect 24222 42030 24274 42082
rect 33406 42030 33458 42082
rect 33742 42030 33794 42082
rect 33854 42030 33906 42082
rect 34302 42030 34354 42082
rect 34414 42030 34466 42082
rect 36766 42030 36818 42082
rect 38110 42030 38162 42082
rect 41246 42030 41298 42082
rect 45726 42030 45778 42082
rect 5070 41918 5122 41970
rect 9662 41918 9714 41970
rect 16718 41918 16770 41970
rect 19630 41918 19682 41970
rect 20302 41918 20354 41970
rect 21534 41918 21586 41970
rect 23214 41918 23266 41970
rect 23662 41918 23714 41970
rect 25118 41918 25170 41970
rect 25454 41918 25506 41970
rect 25790 41918 25842 41970
rect 26686 41918 26738 41970
rect 31502 41918 31554 41970
rect 31950 41918 32002 41970
rect 33070 41918 33122 41970
rect 34078 41918 34130 41970
rect 35422 41918 35474 41970
rect 36094 41918 36146 41970
rect 37438 41918 37490 41970
rect 40014 41918 40066 41970
rect 40910 41918 40962 41970
rect 45838 41918 45890 41970
rect 5518 41806 5570 41858
rect 6190 41806 6242 41858
rect 8990 41806 9042 41858
rect 11342 41806 11394 41858
rect 11790 41806 11842 41858
rect 16046 41806 16098 41858
rect 17502 41806 17554 41858
rect 18958 41806 19010 41858
rect 19182 41806 19234 41858
rect 20078 41806 20130 41858
rect 22318 41806 22370 41858
rect 22766 41806 22818 41858
rect 24110 41806 24162 41858
rect 24670 41806 24722 41858
rect 25342 41806 25394 41858
rect 27470 41806 27522 41858
rect 29598 41806 29650 41858
rect 31054 41806 31106 41858
rect 32398 41806 32450 41858
rect 35646 41806 35698 41858
rect 37214 41806 37266 41858
rect 5070 41694 5122 41746
rect 11006 41694 11058 41746
rect 11342 41694 11394 41746
rect 11790 41694 11842 41746
rect 21310 41694 21362 41746
rect 34414 41694 34466 41746
rect 36654 41694 36706 41746
rect 45726 41694 45778 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 18958 41358 19010 41410
rect 19294 41358 19346 41410
rect 21310 41358 21362 41410
rect 21758 41358 21810 41410
rect 22430 41358 22482 41410
rect 35422 41358 35474 41410
rect 37214 41358 37266 41410
rect 45054 41358 45106 41410
rect 6750 41246 6802 41298
rect 15038 41246 15090 41298
rect 17838 41246 17890 41298
rect 21982 41246 22034 41298
rect 33070 41246 33122 41298
rect 38222 41246 38274 41298
rect 41582 41246 41634 41298
rect 15374 41134 15426 41186
rect 16382 41134 16434 41186
rect 16718 41134 16770 41186
rect 17054 41134 17106 41186
rect 17278 41134 17330 41186
rect 19630 41134 19682 41186
rect 24446 41134 24498 41186
rect 24782 41134 24834 41186
rect 30382 41134 30434 41186
rect 30942 41134 30994 41186
rect 31838 41134 31890 41186
rect 32958 41134 33010 41186
rect 33966 41134 34018 41186
rect 34414 41134 34466 41186
rect 35758 41134 35810 41186
rect 38558 41134 38610 41186
rect 39342 41134 39394 41186
rect 39790 41134 39842 41186
rect 40014 41134 40066 41186
rect 40462 41134 40514 41186
rect 40574 41134 40626 41186
rect 45390 41134 45442 41186
rect 45838 41134 45890 41186
rect 47182 41134 47234 41186
rect 2158 41022 2210 41074
rect 3166 41022 3218 41074
rect 3726 41022 3778 41074
rect 8094 41022 8146 41074
rect 15710 41022 15762 41074
rect 15934 41022 15986 41074
rect 16270 41022 16322 41074
rect 19518 41022 19570 41074
rect 20190 41022 20242 41074
rect 20414 41022 20466 41074
rect 22430 41022 22482 41074
rect 31390 41022 31442 41074
rect 33406 41022 33458 41074
rect 33742 41022 33794 41074
rect 34526 41022 34578 41074
rect 36318 41022 36370 41074
rect 37438 41022 37490 41074
rect 40686 41022 40738 41074
rect 45614 41022 45666 41074
rect 46062 41022 46114 41074
rect 46174 41022 46226 41074
rect 48078 41022 48130 41074
rect 2494 40910 2546 40962
rect 2830 40910 2882 40962
rect 7198 40910 7250 40962
rect 8206 40910 8258 40962
rect 8430 40910 8482 40962
rect 15486 40910 15538 40962
rect 16046 40910 16098 40962
rect 17054 40910 17106 40962
rect 19294 40910 19346 40962
rect 21422 40910 21474 40962
rect 22878 40910 22930 40962
rect 24558 40910 24610 40962
rect 30158 40910 30210 40962
rect 30494 40910 30546 40962
rect 30606 40910 30658 40962
rect 31614 40910 31666 40962
rect 34750 40910 34802 40962
rect 35534 40910 35586 40962
rect 35982 40910 36034 40962
rect 36206 40910 36258 40962
rect 37326 40910 37378 40962
rect 39118 40910 39170 40962
rect 39902 40910 39954 40962
rect 41134 40910 41186 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 4734 40574 4786 40626
rect 5518 40574 5570 40626
rect 9662 40574 9714 40626
rect 16382 40574 16434 40626
rect 16942 40574 16994 40626
rect 21646 40574 21698 40626
rect 23102 40574 23154 40626
rect 23662 40574 23714 40626
rect 24222 40574 24274 40626
rect 31950 40574 32002 40626
rect 32398 40574 32450 40626
rect 34078 40574 34130 40626
rect 34862 40574 34914 40626
rect 38670 40574 38722 40626
rect 39118 40574 39170 40626
rect 41134 40574 41186 40626
rect 41694 40574 41746 40626
rect 42254 40574 42306 40626
rect 42702 40574 42754 40626
rect 2494 40462 2546 40514
rect 7198 40462 7250 40514
rect 8430 40462 8482 40514
rect 11678 40462 11730 40514
rect 12910 40462 12962 40514
rect 16718 40462 16770 40514
rect 18174 40462 18226 40514
rect 21534 40462 21586 40514
rect 22094 40462 22146 40514
rect 22990 40462 23042 40514
rect 23326 40462 23378 40514
rect 23550 40462 23602 40514
rect 33070 40462 33122 40514
rect 33182 40462 33234 40514
rect 34638 40462 34690 40514
rect 40238 40462 40290 40514
rect 41582 40462 41634 40514
rect 44494 40462 44546 40514
rect 45950 40462 46002 40514
rect 1822 40350 1874 40402
rect 5742 40350 5794 40402
rect 8318 40350 8370 40402
rect 11230 40350 11282 40402
rect 12126 40350 12178 40402
rect 16606 40350 16658 40402
rect 17502 40350 17554 40402
rect 20974 40350 21026 40402
rect 22430 40350 22482 40402
rect 22654 40350 22706 40402
rect 25790 40350 25842 40402
rect 26574 40350 26626 40402
rect 30382 40350 30434 40402
rect 30830 40350 30882 40402
rect 31390 40350 31442 40402
rect 31614 40350 31666 40402
rect 34414 40350 34466 40402
rect 35422 40350 35474 40402
rect 35870 40350 35922 40402
rect 37438 40350 37490 40402
rect 38558 40350 38610 40402
rect 38894 40350 38946 40402
rect 39342 40350 39394 40402
rect 39902 40350 39954 40402
rect 41918 40350 41970 40402
rect 43710 40350 43762 40402
rect 45278 40350 45330 40402
rect 10110 40238 10162 40290
rect 15038 40238 15090 40290
rect 20302 40238 20354 40290
rect 22542 40238 22594 40290
rect 24782 40238 24834 40290
rect 28702 40238 28754 40290
rect 34974 40238 35026 40290
rect 35982 40238 36034 40290
rect 37326 40238 37378 40290
rect 43598 40238 43650 40290
rect 45054 40238 45106 40290
rect 6750 40126 6802 40178
rect 21646 40126 21698 40178
rect 23662 40126 23714 40178
rect 23998 40126 24050 40178
rect 24782 40126 24834 40178
rect 33182 40126 33234 40178
rect 36206 40126 36258 40178
rect 37886 40126 37938 40178
rect 42030 40126 42082 40178
rect 42590 40126 42642 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 6862 39790 6914 39842
rect 23102 39790 23154 39842
rect 38894 39790 38946 39842
rect 39342 39790 39394 39842
rect 44158 39790 44210 39842
rect 2494 39678 2546 39730
rect 4622 39678 4674 39730
rect 9214 39678 9266 39730
rect 11902 39678 11954 39730
rect 14254 39678 14306 39730
rect 16382 39678 16434 39730
rect 21758 39678 21810 39730
rect 32062 39678 32114 39730
rect 33630 39678 33682 39730
rect 35982 39678 36034 39730
rect 36318 39678 36370 39730
rect 38446 39678 38498 39730
rect 38894 39678 38946 39730
rect 43038 39678 43090 39730
rect 1822 39566 1874 39618
rect 7086 39566 7138 39618
rect 7422 39566 7474 39618
rect 10558 39566 10610 39618
rect 13470 39566 13522 39618
rect 16942 39566 16994 39618
rect 17278 39566 17330 39618
rect 22430 39566 22482 39618
rect 23214 39566 23266 39618
rect 23550 39566 23602 39618
rect 23886 39566 23938 39618
rect 24222 39566 24274 39618
rect 25342 39566 25394 39618
rect 25902 39566 25954 39618
rect 32286 39566 32338 39618
rect 32622 39566 32674 39618
rect 33182 39566 33234 39618
rect 33518 39566 33570 39618
rect 35086 39566 35138 39618
rect 35870 39566 35922 39618
rect 40238 39566 40290 39618
rect 40910 39566 40962 39618
rect 41582 39566 41634 39618
rect 41918 39566 41970 39618
rect 42590 39566 42642 39618
rect 43486 39566 43538 39618
rect 45054 39566 45106 39618
rect 45502 39566 45554 39618
rect 5966 39454 6018 39506
rect 7982 39454 8034 39506
rect 9214 39454 9266 39506
rect 20750 39454 20802 39506
rect 23662 39454 23714 39506
rect 26014 39454 26066 39506
rect 33966 39454 34018 39506
rect 34750 39454 34802 39506
rect 34862 39454 34914 39506
rect 39342 39454 39394 39506
rect 39678 39454 39730 39506
rect 41246 39454 41298 39506
rect 41694 39454 41746 39506
rect 43934 39454 43986 39506
rect 5630 39342 5682 39394
rect 6526 39342 6578 39394
rect 11118 39342 11170 39394
rect 17166 39342 17218 39394
rect 17838 39342 17890 39394
rect 20414 39342 20466 39394
rect 21310 39342 21362 39394
rect 22542 39342 22594 39394
rect 22766 39342 22818 39394
rect 23102 39342 23154 39394
rect 32398 39342 32450 39394
rect 37998 39342 38050 39394
rect 44046 39342 44098 39394
rect 44830 39342 44882 39394
rect 44942 39342 44994 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 2606 39006 2658 39058
rect 3950 39006 4002 39058
rect 16494 39006 16546 39058
rect 21310 39006 21362 39058
rect 21870 39006 21922 39058
rect 22318 39006 22370 39058
rect 23214 39006 23266 39058
rect 28814 39006 28866 39058
rect 34638 39006 34690 39058
rect 41470 39006 41522 39058
rect 41806 39006 41858 39058
rect 42254 39006 42306 39058
rect 42926 39006 42978 39058
rect 5406 38894 5458 38946
rect 7198 38894 7250 38946
rect 8094 38894 8146 38946
rect 11678 38894 11730 38946
rect 15486 38894 15538 38946
rect 15822 38894 15874 38946
rect 23998 38894 24050 38946
rect 25230 38894 25282 38946
rect 25566 38894 25618 38946
rect 25790 38894 25842 38946
rect 26238 38894 26290 38946
rect 26798 38894 26850 38946
rect 29598 38894 29650 38946
rect 29822 38894 29874 38946
rect 30942 38894 30994 38946
rect 42702 38894 42754 38946
rect 43710 38894 43762 38946
rect 48190 38894 48242 38946
rect 1710 38782 1762 38834
rect 2942 38782 2994 38834
rect 3390 38782 3442 38834
rect 7310 38782 7362 38834
rect 8318 38782 8370 38834
rect 12350 38782 12402 38834
rect 16270 38782 16322 38834
rect 23550 38782 23602 38834
rect 24670 38782 24722 38834
rect 26126 38782 26178 38834
rect 26462 38782 26514 38834
rect 29374 38782 29426 38834
rect 33518 38782 33570 38834
rect 35198 38782 35250 38834
rect 43374 38782 43426 38834
rect 2158 38670 2210 38722
rect 8430 38670 8482 38722
rect 9550 38670 9602 38722
rect 24222 38670 24274 38722
rect 25342 38670 25394 38722
rect 30494 38670 30546 38722
rect 33630 38670 33682 38722
rect 41022 38670 41074 38722
rect 43038 38670 43090 38722
rect 5070 38558 5122 38610
rect 5518 38558 5570 38610
rect 33406 38558 33458 38610
rect 43374 38558 43426 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 8206 38222 8258 38274
rect 20750 38222 20802 38274
rect 24894 38222 24946 38274
rect 34190 38222 34242 38274
rect 1822 38110 1874 38162
rect 8430 38110 8482 38162
rect 9662 38110 9714 38162
rect 11790 38110 11842 38162
rect 15374 38110 15426 38162
rect 17502 38110 17554 38162
rect 28478 38110 28530 38162
rect 34414 38110 34466 38162
rect 34974 38110 35026 38162
rect 38446 38110 38498 38162
rect 3838 37998 3890 38050
rect 8878 37998 8930 38050
rect 14702 37998 14754 38050
rect 18510 37998 18562 38050
rect 19630 37998 19682 38050
rect 25006 37998 25058 38050
rect 27022 37998 27074 38050
rect 27470 37998 27522 38050
rect 29598 37998 29650 38050
rect 29822 37998 29874 38050
rect 29934 37998 29986 38050
rect 38782 37998 38834 38050
rect 39902 37998 39954 38050
rect 18174 37886 18226 37938
rect 29486 37886 29538 37938
rect 30718 37886 30770 37938
rect 30830 37886 30882 37938
rect 3726 37774 3778 37826
rect 7870 37774 7922 37826
rect 24894 37774 24946 37826
rect 25566 37774 25618 37826
rect 30494 37774 30546 37826
rect 33854 37774 33906 37826
rect 38558 37774 38610 37826
rect 39230 37774 39282 37826
rect 39678 37774 39730 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 8990 37438 9042 37490
rect 18062 37438 18114 37490
rect 18286 37438 18338 37490
rect 18510 37438 18562 37490
rect 26574 37438 26626 37490
rect 27246 37438 27298 37490
rect 41918 37438 41970 37490
rect 5070 37326 5122 37378
rect 12350 37326 12402 37378
rect 19518 37326 19570 37378
rect 22654 37326 22706 37378
rect 26686 37326 26738 37378
rect 34974 37326 35026 37378
rect 38110 37326 38162 37378
rect 39566 37326 39618 37378
rect 44270 37326 44322 37378
rect 45950 37326 46002 37378
rect 4398 37214 4450 37266
rect 9550 37214 9602 37266
rect 9774 37214 9826 37266
rect 11566 37214 11618 37266
rect 15710 37214 15762 37266
rect 16270 37214 16322 37266
rect 18622 37214 18674 37266
rect 19854 37214 19906 37266
rect 20862 37214 20914 37266
rect 21982 37214 22034 37266
rect 28030 37214 28082 37266
rect 28142 37214 28194 37266
rect 29598 37214 29650 37266
rect 31278 37214 31330 37266
rect 31502 37214 31554 37266
rect 34750 37214 34802 37266
rect 38446 37214 38498 37266
rect 40910 37214 40962 37266
rect 41134 37214 41186 37266
rect 41806 37214 41858 37266
rect 42142 37214 42194 37266
rect 43374 37214 43426 37266
rect 46846 37214 46898 37266
rect 1822 37102 1874 37154
rect 7198 37102 7250 37154
rect 7646 37102 7698 37154
rect 14478 37102 14530 37154
rect 15374 37102 15426 37154
rect 19966 37102 20018 37154
rect 20414 37102 20466 37154
rect 26126 37102 26178 37154
rect 28590 37102 28642 37154
rect 29262 37102 29314 37154
rect 30158 37102 30210 37154
rect 31838 37102 31890 37154
rect 40238 37102 40290 37154
rect 43486 37102 43538 37154
rect 45390 37102 45442 37154
rect 47854 37102 47906 37154
rect 10110 36990 10162 37042
rect 26574 36990 26626 37042
rect 28478 36990 28530 37042
rect 30830 36990 30882 37042
rect 32062 36990 32114 37042
rect 32398 36990 32450 37042
rect 41470 36990 41522 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19742 36654 19794 36706
rect 22206 36654 22258 36706
rect 23102 36654 23154 36706
rect 28366 36654 28418 36706
rect 45950 36654 46002 36706
rect 2270 36542 2322 36594
rect 4398 36542 4450 36594
rect 8766 36542 8818 36594
rect 10446 36542 10498 36594
rect 12574 36542 12626 36594
rect 14254 36542 14306 36594
rect 17950 36542 18002 36594
rect 18398 36542 18450 36594
rect 19070 36542 19122 36594
rect 20302 36542 20354 36594
rect 22318 36542 22370 36594
rect 22654 36542 22706 36594
rect 23102 36542 23154 36594
rect 27806 36542 27858 36594
rect 29934 36542 29986 36594
rect 30942 36542 30994 36594
rect 46398 36542 46450 36594
rect 4510 36430 4562 36482
rect 5854 36430 5906 36482
rect 7758 36430 7810 36482
rect 7982 36430 8034 36482
rect 8318 36430 8370 36482
rect 9662 36430 9714 36482
rect 14590 36430 14642 36482
rect 23774 36430 23826 36482
rect 25678 36430 25730 36482
rect 26238 36430 26290 36482
rect 27134 36430 27186 36482
rect 28030 36430 28082 36482
rect 30046 36430 30098 36482
rect 32622 36430 32674 36482
rect 39454 36430 39506 36482
rect 39790 36430 39842 36482
rect 41246 36430 41298 36482
rect 41694 36430 41746 36482
rect 45614 36430 45666 36482
rect 46174 36430 46226 36482
rect 46846 36430 46898 36482
rect 3838 36318 3890 36370
rect 5070 36318 5122 36370
rect 17166 36318 17218 36370
rect 19742 36318 19794 36370
rect 19854 36318 19906 36370
rect 23438 36318 23490 36370
rect 30494 36318 30546 36370
rect 31166 36318 31218 36370
rect 33070 36318 33122 36370
rect 39118 36318 39170 36370
rect 39902 36318 39954 36370
rect 40014 36318 40066 36370
rect 40910 36318 40962 36370
rect 1710 36206 1762 36258
rect 4846 36206 4898 36258
rect 5182 36206 5234 36258
rect 5630 36206 5682 36258
rect 5742 36206 5794 36258
rect 6078 36206 6130 36258
rect 7422 36206 7474 36258
rect 8206 36206 8258 36258
rect 17390 36206 17442 36258
rect 24222 36206 24274 36258
rect 25006 36206 25058 36258
rect 38446 36206 38498 36258
rect 38782 36206 38834 36258
rect 40574 36206 40626 36258
rect 46622 36206 46674 36258
rect 46734 36206 46786 36258
rect 48190 36206 48242 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 17726 35870 17778 35922
rect 20974 35870 21026 35922
rect 26350 35870 26402 35922
rect 40014 35870 40066 35922
rect 40350 35870 40402 35922
rect 5294 35758 5346 35810
rect 6862 35758 6914 35810
rect 11566 35758 11618 35810
rect 17950 35758 18002 35810
rect 19742 35758 19794 35810
rect 29374 35758 29426 35810
rect 29486 35758 29538 35810
rect 29934 35758 29986 35810
rect 39678 35758 39730 35810
rect 39790 35758 39842 35810
rect 41134 35758 41186 35810
rect 42366 35758 42418 35810
rect 43038 35758 43090 35810
rect 45390 35758 45442 35810
rect 46846 35758 46898 35810
rect 1822 35646 1874 35698
rect 8094 35646 8146 35698
rect 17502 35646 17554 35698
rect 18174 35646 18226 35698
rect 18846 35646 18898 35698
rect 19182 35646 19234 35698
rect 21758 35646 21810 35698
rect 23550 35646 23602 35698
rect 27806 35646 27858 35698
rect 31054 35646 31106 35698
rect 31838 35646 31890 35698
rect 34414 35646 34466 35698
rect 36430 35646 36482 35698
rect 38110 35646 38162 35698
rect 39006 35646 39058 35698
rect 41358 35646 41410 35698
rect 42478 35646 42530 35698
rect 43374 35646 43426 35698
rect 46174 35646 46226 35698
rect 2494 35534 2546 35586
rect 4622 35534 4674 35586
rect 4958 35534 5010 35586
rect 6974 35534 7026 35586
rect 8430 35534 8482 35586
rect 11230 35534 11282 35586
rect 17838 35534 17890 35586
rect 19070 35534 19122 35586
rect 21310 35534 21362 35586
rect 23438 35534 23490 35586
rect 25902 35534 25954 35586
rect 26798 35534 26850 35586
rect 27358 35534 27410 35586
rect 28254 35534 28306 35586
rect 28702 35534 28754 35586
rect 31390 35534 31442 35586
rect 34862 35534 34914 35586
rect 38558 35534 38610 35586
rect 42366 35534 42418 35586
rect 43262 35534 43314 35586
rect 46062 35534 46114 35586
rect 8654 35422 8706 35474
rect 25790 35422 25842 35474
rect 26350 35422 26402 35474
rect 29486 35422 29538 35474
rect 30494 35422 30546 35474
rect 37214 35422 37266 35474
rect 39006 35422 39058 35474
rect 39342 35422 39394 35474
rect 41694 35422 41746 35474
rect 45502 35422 45554 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 4622 35086 4674 35138
rect 18846 35086 18898 35138
rect 20638 35086 20690 35138
rect 32174 35086 32226 35138
rect 39678 35086 39730 35138
rect 4062 34974 4114 35026
rect 5070 34974 5122 35026
rect 8878 34974 8930 35026
rect 20190 34974 20242 35026
rect 26350 34974 26402 35026
rect 28478 34974 28530 35026
rect 32286 34974 32338 35026
rect 33406 34974 33458 35026
rect 45390 34974 45442 35026
rect 2270 34862 2322 34914
rect 4286 34862 4338 34914
rect 5966 34862 6018 34914
rect 6190 34862 6242 34914
rect 8430 34862 8482 34914
rect 11566 34862 11618 34914
rect 16046 34862 16098 34914
rect 17838 34862 17890 34914
rect 18510 34862 18562 34914
rect 18958 34862 19010 34914
rect 20414 34862 20466 34914
rect 21646 34862 21698 34914
rect 21982 34862 22034 34914
rect 22318 34862 22370 34914
rect 22766 34862 22818 34914
rect 23438 34862 23490 34914
rect 24222 34862 24274 34914
rect 24894 34862 24946 34914
rect 25790 34862 25842 34914
rect 27022 34862 27074 34914
rect 31166 34862 31218 34914
rect 31838 34862 31890 34914
rect 32062 34862 32114 34914
rect 33294 34862 33346 34914
rect 34974 34862 35026 34914
rect 37774 34862 37826 34914
rect 38446 34862 38498 34914
rect 39230 34862 39282 34914
rect 41246 34862 41298 34914
rect 41470 34862 41522 34914
rect 42030 34862 42082 34914
rect 42478 34862 42530 34914
rect 42926 34862 42978 34914
rect 45166 34862 45218 34914
rect 2494 34750 2546 34802
rect 3838 34750 3890 34802
rect 6638 34750 6690 34802
rect 6862 34750 6914 34802
rect 7534 34750 7586 34802
rect 7758 34750 7810 34802
rect 16718 34750 16770 34802
rect 17950 34750 18002 34802
rect 21310 34750 21362 34802
rect 21422 34750 21474 34802
rect 27918 34750 27970 34802
rect 29822 34750 29874 34802
rect 30830 34750 30882 34802
rect 35646 34750 35698 34802
rect 36094 34750 36146 34802
rect 36206 34750 36258 34802
rect 40910 34750 40962 34802
rect 41022 34750 41074 34802
rect 43374 34750 43426 34802
rect 45838 34750 45890 34802
rect 5742 34638 5794 34690
rect 7982 34638 8034 34690
rect 8094 34638 8146 34690
rect 9326 34638 9378 34690
rect 9774 34638 9826 34690
rect 11902 34638 11954 34690
rect 15486 34638 15538 34690
rect 16382 34638 16434 34690
rect 17390 34638 17442 34690
rect 29262 34638 29314 34690
rect 34750 34638 34802 34690
rect 35310 34638 35362 34690
rect 35534 34638 35586 34690
rect 35870 34638 35922 34690
rect 37102 34638 37154 34690
rect 40350 34638 40402 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2718 34302 2770 34354
rect 4286 34302 4338 34354
rect 4622 34302 4674 34354
rect 9102 34302 9154 34354
rect 17726 34302 17778 34354
rect 21422 34302 21474 34354
rect 24558 34302 24610 34354
rect 27022 34302 27074 34354
rect 29038 34302 29090 34354
rect 29486 34302 29538 34354
rect 40238 34302 40290 34354
rect 43598 34302 43650 34354
rect 44830 34302 44882 34354
rect 45502 34302 45554 34354
rect 47742 34302 47794 34354
rect 5182 34190 5234 34242
rect 5742 34190 5794 34242
rect 8542 34190 8594 34242
rect 13918 34190 13970 34242
rect 15934 34190 15986 34242
rect 16494 34190 16546 34242
rect 22094 34190 22146 34242
rect 23662 34190 23714 34242
rect 34190 34190 34242 34242
rect 34638 34190 34690 34242
rect 35198 34190 35250 34242
rect 35870 34190 35922 34242
rect 38110 34190 38162 34242
rect 45054 34190 45106 34242
rect 45726 34190 45778 34242
rect 46622 34190 46674 34242
rect 47182 34190 47234 34242
rect 48190 34190 48242 34242
rect 1710 34078 1762 34130
rect 2270 34078 2322 34130
rect 5070 34078 5122 34130
rect 6526 34078 6578 34130
rect 6862 34078 6914 34130
rect 12014 34078 12066 34130
rect 12462 34078 12514 34130
rect 14702 34078 14754 34130
rect 16270 34078 16322 34130
rect 16830 34078 16882 34130
rect 17390 34078 17442 34130
rect 18846 34078 18898 34130
rect 25454 34078 25506 34130
rect 27918 34078 27970 34130
rect 33294 34078 33346 34130
rect 36878 34078 36930 34130
rect 37774 34078 37826 34130
rect 41022 34078 41074 34130
rect 42926 34078 42978 34130
rect 43262 34078 43314 34130
rect 43486 34078 43538 34130
rect 44270 34078 44322 34130
rect 44494 34078 44546 34130
rect 44718 34078 44770 34130
rect 45278 34078 45330 34130
rect 2718 33966 2770 34018
rect 3390 33966 3442 34018
rect 6190 33966 6242 34018
rect 7982 33966 8034 34018
rect 13582 33966 13634 34018
rect 16382 33966 16434 34018
rect 19294 33966 19346 34018
rect 22318 33966 22370 34018
rect 25566 33966 25618 34018
rect 26574 33966 26626 34018
rect 28254 33966 28306 34018
rect 28590 33966 28642 34018
rect 33406 33966 33458 34018
rect 34750 33966 34802 34018
rect 39678 33966 39730 34018
rect 41694 33966 41746 34018
rect 45390 33966 45442 34018
rect 2942 33854 2994 33906
rect 8430 33854 8482 33906
rect 8878 33854 8930 33906
rect 9102 33854 9154 33906
rect 25902 33854 25954 33906
rect 34862 33854 34914 33906
rect 35310 33854 35362 33906
rect 42702 33854 42754 33906
rect 46510 33854 46562 33906
rect 46846 33854 46898 33906
rect 47294 33854 47346 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 2158 33518 2210 33570
rect 12686 33518 12738 33570
rect 13806 33518 13858 33570
rect 14142 33518 14194 33570
rect 19630 33518 19682 33570
rect 19966 33518 20018 33570
rect 2494 33406 2546 33458
rect 2942 33406 2994 33458
rect 3390 33406 3442 33458
rect 3838 33406 3890 33458
rect 14702 33406 14754 33458
rect 18174 33406 18226 33458
rect 25342 33406 25394 33458
rect 27470 33406 27522 33458
rect 37102 33406 37154 33458
rect 37998 33406 38050 33458
rect 44270 33406 44322 33458
rect 1934 33294 1986 33346
rect 5966 33294 6018 33346
rect 6750 33294 6802 33346
rect 7086 33294 7138 33346
rect 9550 33294 9602 33346
rect 12238 33294 12290 33346
rect 12574 33294 12626 33346
rect 14926 33294 14978 33346
rect 21310 33294 21362 33346
rect 24558 33294 24610 33346
rect 29934 33294 29986 33346
rect 30382 33294 30434 33346
rect 33854 33294 33906 33346
rect 34414 33294 34466 33346
rect 34750 33294 34802 33346
rect 37438 33294 37490 33346
rect 38446 33294 38498 33346
rect 38782 33294 38834 33346
rect 41246 33294 41298 33346
rect 42702 33294 42754 33346
rect 43374 33294 43426 33346
rect 43598 33294 43650 33346
rect 46174 33294 46226 33346
rect 46734 33294 46786 33346
rect 47070 33294 47122 33346
rect 2382 33182 2434 33234
rect 5742 33182 5794 33234
rect 6638 33182 6690 33234
rect 9326 33182 9378 33234
rect 9886 33182 9938 33234
rect 10334 33182 10386 33234
rect 12686 33182 12738 33234
rect 13582 33182 13634 33234
rect 14814 33182 14866 33234
rect 16270 33182 16322 33234
rect 18734 33182 18786 33234
rect 21534 33182 21586 33234
rect 21982 33182 22034 33234
rect 38334 33182 38386 33234
rect 39790 33182 39842 33234
rect 41022 33182 41074 33234
rect 41358 33182 41410 33234
rect 9550 33070 9602 33122
rect 10222 33070 10274 33122
rect 10446 33070 10498 33122
rect 10670 33070 10722 33122
rect 17166 33070 17218 33122
rect 18398 33070 18450 33122
rect 19406 33070 19458 33122
rect 19854 33070 19906 33122
rect 34750 33070 34802 33122
rect 40126 33070 40178 33122
rect 42478 33070 42530 33122
rect 42814 33070 42866 33122
rect 42926 33070 42978 33122
rect 45726 33070 45778 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 1822 32734 1874 32786
rect 4286 32734 4338 32786
rect 4734 32734 4786 32786
rect 8654 32734 8706 32786
rect 9886 32734 9938 32786
rect 12126 32734 12178 32786
rect 14366 32734 14418 32786
rect 19630 32734 19682 32786
rect 21086 32734 21138 32786
rect 22094 32734 22146 32786
rect 28254 32734 28306 32786
rect 34974 32734 35026 32786
rect 38558 32734 38610 32786
rect 39566 32734 39618 32786
rect 41694 32734 41746 32786
rect 3166 32622 3218 32674
rect 8206 32622 8258 32674
rect 9550 32622 9602 32674
rect 11006 32622 11058 32674
rect 15822 32622 15874 32674
rect 17390 32622 17442 32674
rect 19966 32622 20018 32674
rect 20414 32622 20466 32674
rect 20526 32622 20578 32674
rect 30718 32622 30770 32674
rect 33518 32622 33570 32674
rect 37214 32622 37266 32674
rect 38222 32622 38274 32674
rect 38446 32622 38498 32674
rect 39790 32622 39842 32674
rect 40350 32622 40402 32674
rect 40910 32622 40962 32674
rect 41246 32622 41298 32674
rect 46062 32622 46114 32674
rect 48190 32622 48242 32674
rect 2494 32510 2546 32562
rect 2718 32510 2770 32562
rect 2942 32510 2994 32562
rect 5630 32510 5682 32562
rect 6302 32510 6354 32562
rect 7198 32510 7250 32562
rect 7758 32510 7810 32562
rect 12350 32510 12402 32562
rect 13806 32510 13858 32562
rect 14030 32510 14082 32562
rect 17614 32510 17666 32562
rect 18846 32510 18898 32562
rect 21870 32510 21922 32562
rect 22542 32510 22594 32562
rect 22766 32510 22818 32562
rect 23102 32510 23154 32562
rect 25230 32510 25282 32562
rect 31054 32510 31106 32562
rect 32062 32510 32114 32562
rect 33854 32510 33906 32562
rect 34862 32510 34914 32562
rect 37438 32510 37490 32562
rect 38894 32510 38946 32562
rect 47294 32510 47346 32562
rect 3054 32398 3106 32450
rect 3838 32398 3890 32450
rect 5070 32398 5122 32450
rect 6526 32398 6578 32450
rect 7422 32398 7474 32450
rect 18510 32398 18562 32450
rect 21982 32398 22034 32450
rect 22878 32398 22930 32450
rect 24670 32398 24722 32450
rect 26014 32398 26066 32450
rect 30046 32398 30098 32450
rect 31950 32398 32002 32450
rect 47070 32398 47122 32450
rect 5966 32286 6018 32338
rect 11230 32286 11282 32338
rect 11566 32286 11618 32338
rect 16046 32286 16098 32338
rect 16382 32286 16434 32338
rect 18958 32286 19010 32338
rect 20414 32286 20466 32338
rect 31726 32286 31778 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 2718 31950 2770 32002
rect 11454 31950 11506 32002
rect 42702 31950 42754 32002
rect 6414 31838 6466 31890
rect 7310 31838 7362 31890
rect 15710 31838 15762 31890
rect 23326 31838 23378 31890
rect 29262 31838 29314 31890
rect 31726 31838 31778 31890
rect 35646 31838 35698 31890
rect 41134 31838 41186 31890
rect 41358 31838 41410 31890
rect 42254 31838 42306 31890
rect 2158 31726 2210 31778
rect 2494 31726 2546 31778
rect 2830 31726 2882 31778
rect 3838 31726 3890 31778
rect 6638 31726 6690 31778
rect 7422 31726 7474 31778
rect 9326 31726 9378 31778
rect 10670 31726 10722 31778
rect 10894 31726 10946 31778
rect 14590 31726 14642 31778
rect 14926 31726 14978 31778
rect 17390 31726 17442 31778
rect 22094 31726 22146 31778
rect 22654 31726 22706 31778
rect 23550 31726 23602 31778
rect 30718 31726 30770 31778
rect 34414 31726 34466 31778
rect 35534 31726 35586 31778
rect 1934 31614 1986 31666
rect 4846 31614 4898 31666
rect 7758 31614 7810 31666
rect 9550 31614 9602 31666
rect 11118 31614 11170 31666
rect 16046 31614 16098 31666
rect 18398 31614 18450 31666
rect 23886 31614 23938 31666
rect 28590 31614 28642 31666
rect 29486 31614 29538 31666
rect 33294 31614 33346 31666
rect 34526 31614 34578 31666
rect 35982 31614 36034 31666
rect 39790 31614 39842 31666
rect 42590 31614 42642 31666
rect 2606 31502 2658 31554
rect 3278 31502 3330 31554
rect 4622 31502 4674 31554
rect 4958 31502 5010 31554
rect 5182 31502 5234 31554
rect 5966 31502 6018 31554
rect 9998 31502 10050 31554
rect 11902 31502 11954 31554
rect 12238 31502 12290 31554
rect 23774 31502 23826 31554
rect 32958 31502 33010 31554
rect 34750 31502 34802 31554
rect 40686 31502 40738 31554
rect 41694 31502 41746 31554
rect 48190 31502 48242 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 23326 31166 23378 31218
rect 25790 31166 25842 31218
rect 27246 31166 27298 31218
rect 6862 31054 6914 31106
rect 7870 31054 7922 31106
rect 8094 31054 8146 31106
rect 10894 31054 10946 31106
rect 11230 31054 11282 31106
rect 17502 31054 17554 31106
rect 20750 31054 20802 31106
rect 21422 31054 21474 31106
rect 27470 31054 27522 31106
rect 29934 31054 29986 31106
rect 32062 31054 32114 31106
rect 34414 31054 34466 31106
rect 42478 31054 42530 31106
rect 1710 30942 1762 30994
rect 5518 30942 5570 30994
rect 6414 30942 6466 30994
rect 8318 30942 8370 30994
rect 8430 30942 8482 30994
rect 9662 30942 9714 30994
rect 9886 30942 9938 30994
rect 12238 30942 12290 30994
rect 13246 30942 13298 30994
rect 14030 30942 14082 30994
rect 14366 30942 14418 30994
rect 14926 30942 14978 30994
rect 16158 30942 16210 30994
rect 17390 30942 17442 30994
rect 18286 30942 18338 30994
rect 20078 30942 20130 30994
rect 21198 30942 21250 30994
rect 23550 30942 23602 30994
rect 25566 30942 25618 30994
rect 28478 30942 28530 30994
rect 28814 30942 28866 30994
rect 29038 30942 29090 30994
rect 30830 30942 30882 30994
rect 31838 30942 31890 30994
rect 36206 30942 36258 30994
rect 36542 30942 36594 30994
rect 37550 30942 37602 30994
rect 37886 30942 37938 30994
rect 38558 30942 38610 30994
rect 41582 30942 41634 30994
rect 41806 30942 41858 30994
rect 2494 30830 2546 30882
rect 4622 30830 4674 30882
rect 4958 30830 5010 30882
rect 10558 30830 10610 30882
rect 11790 30830 11842 30882
rect 15374 30830 15426 30882
rect 16718 30830 16770 30882
rect 18062 30830 18114 30882
rect 20526 30830 20578 30882
rect 40910 30830 40962 30882
rect 42590 30830 42642 30882
rect 8878 30718 8930 30770
rect 16382 30718 16434 30770
rect 29150 30718 29202 30770
rect 34526 30718 34578 30770
rect 35310 30718 35362 30770
rect 42254 30718 42306 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 4510 30270 4562 30322
rect 6638 30270 6690 30322
rect 14142 30270 14194 30322
rect 15150 30270 15202 30322
rect 16046 30270 16098 30322
rect 16382 30270 16434 30322
rect 16606 30270 16658 30322
rect 18062 30270 18114 30322
rect 20750 30270 20802 30322
rect 29934 30270 29986 30322
rect 1934 30158 1986 30210
rect 2942 30158 2994 30210
rect 4398 30158 4450 30210
rect 5182 30158 5234 30210
rect 6526 30158 6578 30210
rect 8542 30158 8594 30210
rect 10110 30158 10162 30210
rect 12126 30158 12178 30210
rect 12910 30158 12962 30210
rect 2606 30046 2658 30098
rect 4286 30046 4338 30098
rect 7758 30046 7810 30098
rect 8094 30046 8146 30098
rect 11342 30046 11394 30098
rect 12574 30046 12626 30098
rect 12686 30046 12738 30098
rect 14478 30102 14530 30154
rect 14814 30158 14866 30210
rect 15598 30158 15650 30210
rect 16718 30158 16770 30210
rect 19406 30158 19458 30210
rect 21422 30158 21474 30210
rect 23550 30158 23602 30210
rect 27246 30158 27298 30210
rect 27582 30158 27634 30210
rect 28254 30158 28306 30210
rect 28478 30158 28530 30210
rect 31950 30158 32002 30210
rect 32622 30158 32674 30210
rect 33070 30158 33122 30210
rect 35422 30158 35474 30210
rect 36990 30158 37042 30210
rect 37102 30158 37154 30210
rect 37438 30158 37490 30210
rect 40350 30158 40402 30210
rect 41134 30158 41186 30210
rect 41806 30158 41858 30210
rect 42366 30158 42418 30210
rect 17278 30046 17330 30098
rect 17390 30046 17442 30098
rect 18174 30046 18226 30098
rect 21758 30046 21810 30098
rect 22654 30046 22706 30098
rect 23214 30046 23266 30098
rect 29262 30046 29314 30098
rect 29374 30046 29426 30098
rect 32062 30046 32114 30098
rect 35870 30046 35922 30098
rect 36094 30046 36146 30098
rect 40574 30046 40626 30098
rect 40686 30046 40738 30098
rect 41582 30046 41634 30098
rect 43934 30046 43986 30098
rect 2270 29934 2322 29986
rect 3502 29934 3554 29986
rect 5742 29934 5794 29986
rect 9662 29934 9714 29986
rect 14590 29934 14642 29986
rect 17614 29934 17666 29986
rect 21870 29934 21922 29986
rect 22766 29934 22818 29986
rect 29038 29934 29090 29986
rect 35982 29934 36034 29986
rect 38446 29934 38498 29986
rect 40014 29934 40066 29986
rect 42478 29934 42530 29986
rect 44046 29934 44098 29986
rect 44270 29934 44322 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5406 29598 5458 29650
rect 5966 29598 6018 29650
rect 7534 29598 7586 29650
rect 7982 29598 8034 29650
rect 8990 29598 9042 29650
rect 12014 29598 12066 29650
rect 12574 29598 12626 29650
rect 20638 29598 20690 29650
rect 24670 29598 24722 29650
rect 30046 29598 30098 29650
rect 39566 29598 39618 29650
rect 40350 29598 40402 29650
rect 41246 29598 41298 29650
rect 47518 29598 47570 29650
rect 5630 29486 5682 29538
rect 5742 29486 5794 29538
rect 11230 29486 11282 29538
rect 14702 29486 14754 29538
rect 14814 29486 14866 29538
rect 18622 29486 18674 29538
rect 18846 29486 18898 29538
rect 21758 29486 21810 29538
rect 27358 29486 27410 29538
rect 28254 29486 28306 29538
rect 32510 29486 32562 29538
rect 36430 29486 36482 29538
rect 38334 29486 38386 29538
rect 39118 29486 39170 29538
rect 41358 29486 41410 29538
rect 42590 29486 42642 29538
rect 43374 29486 43426 29538
rect 45278 29486 45330 29538
rect 45950 29486 46002 29538
rect 1710 29374 1762 29426
rect 2270 29374 2322 29426
rect 9550 29374 9602 29426
rect 9774 29374 9826 29426
rect 10446 29374 10498 29426
rect 10670 29374 10722 29426
rect 10894 29374 10946 29426
rect 11902 29374 11954 29426
rect 12238 29374 12290 29426
rect 22094 29374 22146 29426
rect 25454 29374 25506 29426
rect 26798 29374 26850 29426
rect 29710 29374 29762 29426
rect 31614 29374 31666 29426
rect 31950 29374 32002 29426
rect 37326 29374 37378 29426
rect 40910 29374 40962 29426
rect 41470 29374 41522 29426
rect 42702 29374 42754 29426
rect 43934 29374 43986 29426
rect 44606 29374 44658 29426
rect 47182 29374 47234 29426
rect 4846 29262 4898 29314
rect 15374 29262 15426 29314
rect 18846 29262 18898 29314
rect 25902 29262 25954 29314
rect 28030 29262 28082 29314
rect 35870 29262 35922 29314
rect 45726 29262 45778 29314
rect 9998 29150 10050 29202
rect 14814 29150 14866 29202
rect 39006 29150 39058 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 10782 28814 10834 28866
rect 27582 28814 27634 28866
rect 33742 28814 33794 28866
rect 35534 28814 35586 28866
rect 39454 28814 39506 28866
rect 40462 28814 40514 28866
rect 47070 28814 47122 28866
rect 2494 28702 2546 28754
rect 4622 28702 4674 28754
rect 12014 28702 12066 28754
rect 17054 28702 17106 28754
rect 18510 28702 18562 28754
rect 20190 28702 20242 28754
rect 24222 28702 24274 28754
rect 27022 28702 27074 28754
rect 27470 28702 27522 28754
rect 38670 28702 38722 28754
rect 40238 28702 40290 28754
rect 41246 28702 41298 28754
rect 43486 28702 43538 28754
rect 43710 28702 43762 28754
rect 45278 28702 45330 28754
rect 46622 28702 46674 28754
rect 1710 28590 1762 28642
rect 5070 28590 5122 28642
rect 5742 28590 5794 28642
rect 9550 28590 9602 28642
rect 11230 28590 11282 28642
rect 14590 28590 14642 28642
rect 18846 28590 18898 28642
rect 18958 28590 19010 28642
rect 19182 28590 19234 28642
rect 19294 28590 19346 28642
rect 19854 28590 19906 28642
rect 20414 28590 20466 28642
rect 21534 28590 21586 28642
rect 22654 28590 22706 28642
rect 25454 28590 25506 28642
rect 25790 28590 25842 28642
rect 27582 28590 27634 28642
rect 28702 28590 28754 28642
rect 38558 28590 38610 28642
rect 44718 28590 44770 28642
rect 46734 28590 46786 28642
rect 10110 28478 10162 28530
rect 10670 28478 10722 28530
rect 10782 28478 10834 28530
rect 11566 28478 11618 28530
rect 14702 28478 14754 28530
rect 16494 28478 16546 28530
rect 16606 28478 16658 28530
rect 22094 28478 22146 28530
rect 22430 28478 22482 28530
rect 32622 28478 32674 28530
rect 33630 28478 33682 28530
rect 33742 28478 33794 28530
rect 35198 28478 35250 28530
rect 35422 28478 35474 28530
rect 35870 28478 35922 28530
rect 35982 28478 36034 28530
rect 37326 28478 37378 28530
rect 37662 28478 37714 28530
rect 39006 28478 39058 28530
rect 39342 28478 39394 28530
rect 45166 28478 45218 28530
rect 45390 28478 45442 28530
rect 48190 28478 48242 28530
rect 5742 28366 5794 28418
rect 9774 28366 9826 28418
rect 14926 28366 14978 28418
rect 16270 28366 16322 28418
rect 32734 28366 32786 28418
rect 32958 28366 33010 28418
rect 36206 28366 36258 28418
rect 39454 28366 39506 28418
rect 40798 28366 40850 28418
rect 43710 28366 43762 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 2494 28030 2546 28082
rect 3390 28030 3442 28082
rect 8542 28030 8594 28082
rect 11566 28030 11618 28082
rect 12350 28030 12402 28082
rect 12574 28030 12626 28082
rect 25902 28030 25954 28082
rect 33182 28030 33234 28082
rect 40238 28030 40290 28082
rect 46510 28030 46562 28082
rect 8878 27918 8930 27970
rect 8990 27918 9042 27970
rect 10110 27918 10162 27970
rect 11342 27918 11394 27970
rect 11678 27918 11730 27970
rect 14478 27918 14530 27970
rect 20414 27918 20466 27970
rect 20638 27918 20690 27970
rect 21534 27918 21586 27970
rect 23102 27918 23154 27970
rect 25678 27918 25730 27970
rect 26014 27918 26066 27970
rect 27582 27918 27634 27970
rect 29710 27918 29762 27970
rect 33070 27918 33122 27970
rect 33966 27918 34018 27970
rect 36094 27918 36146 27970
rect 37550 27918 37602 27970
rect 39790 27918 39842 27970
rect 2270 27806 2322 27858
rect 2942 27806 2994 27858
rect 8654 27806 8706 27858
rect 9886 27806 9938 27858
rect 10446 27806 10498 27858
rect 11006 27806 11058 27858
rect 11790 27806 11842 27858
rect 12014 27806 12066 27858
rect 12910 27806 12962 27858
rect 14814 27806 14866 27858
rect 15822 27806 15874 27858
rect 16494 27806 16546 27858
rect 19070 27806 19122 27858
rect 19406 27806 19458 27858
rect 21870 27806 21922 27858
rect 26126 27806 26178 27858
rect 28030 27806 28082 27858
rect 28478 27806 28530 27858
rect 30158 27806 30210 27858
rect 34974 27806 35026 27858
rect 35758 27806 35810 27858
rect 38558 27806 38610 27858
rect 40350 27806 40402 27858
rect 46622 27806 46674 27858
rect 1822 27694 1874 27746
rect 12462 27694 12514 27746
rect 15710 27694 15762 27746
rect 19854 27694 19906 27746
rect 20526 27694 20578 27746
rect 23438 27694 23490 27746
rect 23774 27694 23826 27746
rect 30606 27694 30658 27746
rect 36990 27694 37042 27746
rect 16382 27582 16434 27634
rect 18062 27582 18114 27634
rect 23998 27582 24050 27634
rect 24334 27582 24386 27634
rect 33182 27582 33234 27634
rect 40238 27582 40290 27634
rect 46510 27582 46562 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 18398 27246 18450 27298
rect 19182 27246 19234 27298
rect 19854 27246 19906 27298
rect 21870 27246 21922 27298
rect 35310 27246 35362 27298
rect 37662 27246 37714 27298
rect 37998 27246 38050 27298
rect 41246 27246 41298 27298
rect 2158 27134 2210 27186
rect 6750 27134 6802 27186
rect 8878 27134 8930 27186
rect 12910 27134 12962 27186
rect 17726 27134 17778 27186
rect 19406 27134 19458 27186
rect 19966 27134 20018 27186
rect 20638 27134 20690 27186
rect 22766 27134 22818 27186
rect 25566 27134 25618 27186
rect 31054 27134 31106 27186
rect 31950 27134 32002 27186
rect 35534 27134 35586 27186
rect 1822 27022 1874 27074
rect 3278 27022 3330 27074
rect 8430 27022 8482 27074
rect 12350 27022 12402 27074
rect 12798 27022 12850 27074
rect 13582 27022 13634 27074
rect 13806 27022 13858 27074
rect 15934 27022 15986 27074
rect 17054 27022 17106 27074
rect 17614 27022 17666 27074
rect 20750 27022 20802 27074
rect 21646 27022 21698 27074
rect 24222 27022 24274 27074
rect 28254 27022 28306 27074
rect 30830 27022 30882 27074
rect 31614 27022 31666 27074
rect 32622 27022 32674 27074
rect 33406 27022 33458 27074
rect 35422 27022 35474 27074
rect 36206 27022 36258 27074
rect 37438 27022 37490 27074
rect 39006 27022 39058 27074
rect 39902 27022 39954 27074
rect 2606 26910 2658 26962
rect 2942 26910 2994 26962
rect 3614 26910 3666 26962
rect 4062 26910 4114 26962
rect 5854 26910 5906 26962
rect 7758 26910 7810 26962
rect 8206 26910 8258 26962
rect 10334 26910 10386 26962
rect 10670 26910 10722 26962
rect 11006 26910 11058 26962
rect 12126 26910 12178 26962
rect 14478 26910 14530 26962
rect 16942 26910 16994 26962
rect 22990 26910 23042 26962
rect 28142 26910 28194 26962
rect 30270 26910 30322 26962
rect 33854 26910 33906 26962
rect 38782 26910 38834 26962
rect 45614 26910 45666 26962
rect 45726 26910 45778 26962
rect 6190 26798 6242 26850
rect 9998 26798 10050 26850
rect 12574 26798 12626 26850
rect 16158 26798 16210 26850
rect 22206 26798 22258 26850
rect 27694 26798 27746 26850
rect 27918 26798 27970 26850
rect 45950 26798 46002 26850
rect 48190 26798 48242 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 13806 26462 13858 26514
rect 14478 26462 14530 26514
rect 22094 26462 22146 26514
rect 30942 26462 30994 26514
rect 31054 26462 31106 26514
rect 31614 26462 31666 26514
rect 31838 26462 31890 26514
rect 38334 26462 38386 26514
rect 2718 26350 2770 26402
rect 6414 26350 6466 26402
rect 10110 26350 10162 26402
rect 10894 26350 10946 26402
rect 12462 26350 12514 26402
rect 12686 26350 12738 26402
rect 14142 26350 14194 26402
rect 16270 26350 16322 26402
rect 18958 26350 19010 26402
rect 20862 26350 20914 26402
rect 28926 26350 28978 26402
rect 31502 26350 31554 26402
rect 33070 26350 33122 26402
rect 45166 26350 45218 26402
rect 47406 26350 47458 26402
rect 2046 26238 2098 26290
rect 5630 26238 5682 26290
rect 8990 26238 9042 26290
rect 9886 26238 9938 26290
rect 13246 26238 13298 26290
rect 13470 26238 13522 26290
rect 15262 26238 15314 26290
rect 20190 26238 20242 26290
rect 22430 26238 22482 26290
rect 23102 26238 23154 26290
rect 23438 26238 23490 26290
rect 23774 26238 23826 26290
rect 23998 26238 24050 26290
rect 27694 26238 27746 26290
rect 28142 26238 28194 26290
rect 28478 26238 28530 26290
rect 29038 26238 29090 26290
rect 29150 26238 29202 26290
rect 33518 26238 33570 26290
rect 43710 26238 43762 26290
rect 46286 26238 46338 26290
rect 4846 26126 4898 26178
rect 5294 26126 5346 26178
rect 8542 26126 8594 26178
rect 10558 26126 10610 26178
rect 15150 26126 15202 26178
rect 18510 26126 18562 26178
rect 27134 26126 27186 26178
rect 33854 26126 33906 26178
rect 43374 26126 43426 26178
rect 44158 26126 44210 26178
rect 44830 26126 44882 26178
rect 15822 26014 15874 26066
rect 16494 26014 16546 26066
rect 16830 26014 16882 26066
rect 24110 26014 24162 26066
rect 27470 26014 27522 26066
rect 31166 26014 31218 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 14254 25678 14306 25730
rect 25790 25678 25842 25730
rect 4286 25566 4338 25618
rect 5070 25566 5122 25618
rect 7758 25566 7810 25618
rect 9998 25566 10050 25618
rect 11790 25566 11842 25618
rect 15822 25566 15874 25618
rect 16606 25566 16658 25618
rect 18398 25566 18450 25618
rect 27582 25566 27634 25618
rect 32286 25566 32338 25618
rect 34078 25566 34130 25618
rect 37214 25566 37266 25618
rect 43710 25566 43762 25618
rect 45390 25566 45442 25618
rect 45838 25566 45890 25618
rect 4622 25454 4674 25506
rect 5630 25454 5682 25506
rect 5854 25454 5906 25506
rect 6302 25454 6354 25506
rect 7422 25454 7474 25506
rect 8094 25454 8146 25506
rect 8542 25454 8594 25506
rect 9102 25454 9154 25506
rect 12126 25454 12178 25506
rect 14142 25454 14194 25506
rect 14702 25454 14754 25506
rect 16158 25454 16210 25506
rect 16942 25454 16994 25506
rect 18286 25454 18338 25506
rect 20750 25454 20802 25506
rect 21534 25454 21586 25506
rect 23326 25454 23378 25506
rect 25230 25454 25282 25506
rect 25454 25454 25506 25506
rect 28030 25454 28082 25506
rect 28590 25454 28642 25506
rect 32174 25454 32226 25506
rect 41022 25454 41074 25506
rect 41694 25454 41746 25506
rect 42814 25454 42866 25506
rect 43150 25454 43202 25506
rect 45166 25454 45218 25506
rect 46398 25454 46450 25506
rect 14814 25342 14866 25394
rect 15038 25342 15090 25394
rect 19070 25342 19122 25394
rect 20414 25342 20466 25394
rect 21422 25342 21474 25394
rect 23102 25342 23154 25394
rect 27918 25342 27970 25394
rect 32622 25342 32674 25394
rect 40574 25342 40626 25394
rect 46286 25342 46338 25394
rect 12238 25230 12290 25282
rect 12462 25230 12514 25282
rect 14254 25230 14306 25282
rect 17278 25230 17330 25282
rect 21198 25230 21250 25282
rect 26462 25230 26514 25282
rect 29262 25230 29314 25282
rect 33966 25230 34018 25282
rect 42142 25230 42194 25282
rect 46062 25230 46114 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 5294 24894 5346 24946
rect 6862 24894 6914 24946
rect 11118 24894 11170 24946
rect 18174 24894 18226 24946
rect 18398 24894 18450 24946
rect 18958 24894 19010 24946
rect 21310 24894 21362 24946
rect 23550 24894 23602 24946
rect 28702 24894 28754 24946
rect 32398 24894 32450 24946
rect 36878 24894 36930 24946
rect 37886 24894 37938 24946
rect 38446 24894 38498 24946
rect 39118 24894 39170 24946
rect 39566 24894 39618 24946
rect 4734 24782 4786 24834
rect 5182 24782 5234 24834
rect 5854 24782 5906 24834
rect 6750 24782 6802 24834
rect 12798 24782 12850 24834
rect 14702 24782 14754 24834
rect 19630 24782 19682 24834
rect 20862 24782 20914 24834
rect 25230 24782 25282 24834
rect 27134 24782 27186 24834
rect 28814 24782 28866 24834
rect 31950 24782 32002 24834
rect 32286 24782 32338 24834
rect 37438 24782 37490 24834
rect 37998 24782 38050 24834
rect 39454 24782 39506 24834
rect 40014 24782 40066 24834
rect 42254 24782 42306 24834
rect 43038 24782 43090 24834
rect 4846 24670 4898 24722
rect 6078 24670 6130 24722
rect 7086 24670 7138 24722
rect 7310 24670 7362 24722
rect 8318 24670 8370 24722
rect 10782 24670 10834 24722
rect 14366 24670 14418 24722
rect 18062 24670 18114 24722
rect 19406 24670 19458 24722
rect 20078 24670 20130 24722
rect 20302 24670 20354 24722
rect 22990 24670 23042 24722
rect 23214 24670 23266 24722
rect 25454 24670 25506 24722
rect 25902 24670 25954 24722
rect 27582 24670 27634 24722
rect 31502 24670 31554 24722
rect 31838 24670 31890 24722
rect 32622 24670 32674 24722
rect 32958 24670 33010 24722
rect 33966 24670 34018 24722
rect 35422 24670 35474 24722
rect 37214 24670 37266 24722
rect 39790 24670 39842 24722
rect 40350 24670 40402 24722
rect 42478 24670 42530 24722
rect 42926 24670 42978 24722
rect 43822 24670 43874 24722
rect 44046 24670 44098 24722
rect 44382 24670 44434 24722
rect 44718 24670 44770 24722
rect 45054 24670 45106 24722
rect 45390 24670 45442 24722
rect 8206 24558 8258 24610
rect 14590 24558 14642 24610
rect 19070 24558 19122 24610
rect 19854 24558 19906 24610
rect 29486 24558 29538 24610
rect 29934 24558 29986 24610
rect 33630 24558 33682 24610
rect 34974 24558 35026 24610
rect 35870 24558 35922 24610
rect 43150 24558 43202 24610
rect 45166 24558 45218 24610
rect 4734 24446 4786 24498
rect 5294 24446 5346 24498
rect 8318 24446 8370 24498
rect 13806 24446 13858 24498
rect 18734 24446 18786 24498
rect 33742 24446 33794 24498
rect 37886 24446 37938 24498
rect 40350 24446 40402 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 43710 24110 43762 24162
rect 44158 24110 44210 24162
rect 2270 23998 2322 24050
rect 29150 23998 29202 24050
rect 29598 23998 29650 24050
rect 31838 23998 31890 24050
rect 36094 23998 36146 24050
rect 39230 23998 39282 24050
rect 41246 23998 41298 24050
rect 43038 23998 43090 24050
rect 43710 23998 43762 24050
rect 44158 23998 44210 24050
rect 46734 23998 46786 24050
rect 6414 23886 6466 23938
rect 6750 23886 6802 23938
rect 11454 23886 11506 23938
rect 11678 23886 11730 23938
rect 11902 23886 11954 23938
rect 12126 23886 12178 23938
rect 13582 23886 13634 23938
rect 20638 23886 20690 23938
rect 21534 23886 21586 23938
rect 23214 23886 23266 23938
rect 23550 23886 23602 23938
rect 23886 23886 23938 23938
rect 25454 23886 25506 23938
rect 26350 23886 26402 23938
rect 29822 23886 29874 23938
rect 31166 23886 31218 23938
rect 31950 23886 32002 23938
rect 32958 23886 33010 23938
rect 34190 23886 34242 23938
rect 35198 23886 35250 23938
rect 37326 23886 37378 23938
rect 37662 23886 37714 23938
rect 38334 23886 38386 23938
rect 38894 23886 38946 23938
rect 39678 23886 39730 23938
rect 40350 23886 40402 23938
rect 40798 23886 40850 23938
rect 41694 23886 41746 23938
rect 42926 23886 42978 23938
rect 46958 23886 47010 23938
rect 1710 23774 1762 23826
rect 6638 23774 6690 23826
rect 10222 23774 10274 23826
rect 10670 23774 10722 23826
rect 13806 23774 13858 23826
rect 19966 23774 20018 23826
rect 20190 23774 20242 23826
rect 20862 23774 20914 23826
rect 21310 23774 21362 23826
rect 22878 23774 22930 23826
rect 25118 23774 25170 23826
rect 25678 23774 25730 23826
rect 32622 23774 32674 23826
rect 33854 23774 33906 23826
rect 37998 23774 38050 23826
rect 40910 23774 40962 23826
rect 41918 23774 41970 23826
rect 42702 23774 42754 23826
rect 48078 23774 48130 23826
rect 9662 23662 9714 23714
rect 10894 23662 10946 23714
rect 11006 23662 11058 23714
rect 11118 23662 11170 23714
rect 11342 23662 11394 23714
rect 21870 23662 21922 23714
rect 22990 23662 23042 23714
rect 26462 23662 26514 23714
rect 30942 23662 30994 23714
rect 33070 23662 33122 23714
rect 37662 23662 37714 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 1822 23326 1874 23378
rect 6862 23326 6914 23378
rect 14702 23326 14754 23378
rect 23998 23326 24050 23378
rect 29822 23326 29874 23378
rect 38782 23326 38834 23378
rect 40798 23326 40850 23378
rect 41022 23326 41074 23378
rect 41582 23326 41634 23378
rect 45838 23326 45890 23378
rect 5854 23214 5906 23266
rect 9550 23214 9602 23266
rect 13358 23214 13410 23266
rect 13918 23214 13970 23266
rect 14590 23214 14642 23266
rect 15486 23214 15538 23266
rect 15598 23214 15650 23266
rect 16158 23214 16210 23266
rect 19294 23214 19346 23266
rect 21310 23214 21362 23266
rect 22878 23214 22930 23266
rect 23886 23214 23938 23266
rect 26126 23214 26178 23266
rect 29710 23214 29762 23266
rect 35534 23214 35586 23266
rect 38110 23214 38162 23266
rect 41134 23214 41186 23266
rect 4734 23102 4786 23154
rect 11790 23102 11842 23154
rect 12798 23102 12850 23154
rect 14254 23102 14306 23154
rect 15822 23102 15874 23154
rect 21422 23102 21474 23154
rect 22318 23102 22370 23154
rect 24222 23102 24274 23154
rect 25342 23102 25394 23154
rect 26686 23102 26738 23154
rect 27246 23102 27298 23154
rect 27582 23102 27634 23154
rect 28478 23102 28530 23154
rect 29150 23102 29202 23154
rect 30046 23102 30098 23154
rect 33966 23102 34018 23154
rect 37102 23102 37154 23154
rect 39342 23102 39394 23154
rect 39678 23102 39730 23154
rect 40238 23102 40290 23154
rect 45726 23102 45778 23154
rect 4062 22990 4114 23042
rect 6190 22990 6242 23042
rect 12238 22990 12290 23042
rect 13022 22990 13074 23042
rect 20302 22990 20354 23042
rect 25790 22990 25842 23042
rect 26238 22990 26290 23042
rect 28142 22990 28194 23042
rect 34078 22990 34130 23042
rect 35310 22990 35362 23042
rect 10558 22878 10610 22930
rect 12126 22878 12178 22930
rect 14702 22878 14754 22930
rect 34750 22878 34802 22930
rect 39566 22878 39618 22930
rect 45838 22878 45890 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 15710 22542 15762 22594
rect 42590 22542 42642 22594
rect 8542 22430 8594 22482
rect 11790 22430 11842 22482
rect 12910 22430 12962 22482
rect 14702 22430 14754 22482
rect 15038 22430 15090 22482
rect 15486 22430 15538 22482
rect 19406 22430 19458 22482
rect 19742 22430 19794 22482
rect 20302 22430 20354 22482
rect 22094 22430 22146 22482
rect 25902 22430 25954 22482
rect 29262 22430 29314 22482
rect 36990 22430 37042 22482
rect 37438 22430 37490 22482
rect 38446 22430 38498 22482
rect 40014 22430 40066 22482
rect 40574 22430 40626 22482
rect 41022 22430 41074 22482
rect 42254 22430 42306 22482
rect 45502 22430 45554 22482
rect 45950 22430 46002 22482
rect 7086 22318 7138 22370
rect 7422 22318 7474 22370
rect 7758 22318 7810 22370
rect 8430 22318 8482 22370
rect 9326 22318 9378 22370
rect 9774 22318 9826 22370
rect 9998 22318 10050 22370
rect 11566 22318 11618 22370
rect 11678 22318 11730 22370
rect 11902 22318 11954 22370
rect 12014 22318 12066 22370
rect 14590 22318 14642 22370
rect 16718 22318 16770 22370
rect 18174 22318 18226 22370
rect 20078 22318 20130 22370
rect 21758 22318 21810 22370
rect 22206 22318 22258 22370
rect 27246 22318 27298 22370
rect 37662 22318 37714 22370
rect 39454 22318 39506 22370
rect 42030 22318 42082 22370
rect 46174 22318 46226 22370
rect 10670 22206 10722 22258
rect 17614 22206 17666 22258
rect 22878 22206 22930 22258
rect 38334 22206 38386 22258
rect 38558 22206 38610 22258
rect 39790 22206 39842 22258
rect 46846 22206 46898 22258
rect 47070 22206 47122 22258
rect 7534 22094 7586 22146
rect 16046 22094 16098 22146
rect 16830 22094 16882 22146
rect 17054 22094 17106 22146
rect 17278 22094 17330 22146
rect 18510 22094 18562 22146
rect 18846 22094 18898 22146
rect 27582 22094 27634 22146
rect 40462 22094 40514 22146
rect 46958 22094 47010 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 10222 21758 10274 21810
rect 10782 21758 10834 21810
rect 10894 21758 10946 21810
rect 11454 21758 11506 21810
rect 13582 21758 13634 21810
rect 13918 21758 13970 21810
rect 14926 21758 14978 21810
rect 18398 21758 18450 21810
rect 20190 21758 20242 21810
rect 20526 21758 20578 21810
rect 45278 21758 45330 21810
rect 45502 21758 45554 21810
rect 46398 21758 46450 21810
rect 17726 21646 17778 21698
rect 18286 21646 18338 21698
rect 26126 21646 26178 21698
rect 29038 21646 29090 21698
rect 30494 21646 30546 21698
rect 30606 21646 30658 21698
rect 31726 21646 31778 21698
rect 42254 21646 42306 21698
rect 44830 21646 44882 21698
rect 1710 21534 1762 21586
rect 2270 21534 2322 21586
rect 5070 21534 5122 21586
rect 8318 21534 8370 21586
rect 14814 21534 14866 21586
rect 15150 21534 15202 21586
rect 15710 21534 15762 21586
rect 16494 21534 16546 21586
rect 17614 21534 17666 21586
rect 18622 21534 18674 21586
rect 20638 21534 20690 21586
rect 25342 21534 25394 21586
rect 27358 21534 27410 21586
rect 29710 21534 29762 21586
rect 30270 21534 30322 21586
rect 42702 21534 42754 21586
rect 43486 21534 43538 21586
rect 45838 21534 45890 21586
rect 46958 21534 47010 21586
rect 5742 21422 5794 21474
rect 7870 21422 7922 21474
rect 9662 21422 9714 21474
rect 15822 21422 15874 21474
rect 25790 21422 25842 21474
rect 27022 21422 27074 21474
rect 28366 21422 28418 21474
rect 29934 21422 29986 21474
rect 45390 21422 45442 21474
rect 48078 21422 48130 21474
rect 10670 21310 10722 21362
rect 17726 21310 17778 21362
rect 20526 21310 20578 21362
rect 31614 21310 31666 21362
rect 31950 21310 32002 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17390 20974 17442 21026
rect 27022 20974 27074 21026
rect 29598 20974 29650 21026
rect 31278 20974 31330 21026
rect 37774 20974 37826 21026
rect 37998 20974 38050 21026
rect 38558 20974 38610 21026
rect 41470 20974 41522 21026
rect 1822 20862 1874 20914
rect 17166 20862 17218 20914
rect 18958 20862 19010 20914
rect 19630 20862 19682 20914
rect 25230 20862 25282 20914
rect 27358 20862 27410 20914
rect 28590 20862 28642 20914
rect 30046 20862 30098 20914
rect 32622 20862 32674 20914
rect 39118 20862 39170 20914
rect 45614 20862 45666 20914
rect 5966 20750 6018 20802
rect 10110 20750 10162 20802
rect 15486 20750 15538 20802
rect 15710 20750 15762 20802
rect 16046 20750 16098 20802
rect 16942 20750 16994 20802
rect 19294 20750 19346 20802
rect 20302 20750 20354 20802
rect 25902 20750 25954 20802
rect 26126 20750 26178 20802
rect 27246 20750 27298 20802
rect 30158 20750 30210 20802
rect 31614 20750 31666 20802
rect 32958 20750 33010 20802
rect 45390 20750 45442 20802
rect 46734 20750 46786 20802
rect 5742 20638 5794 20690
rect 10558 20638 10610 20690
rect 15598 20638 15650 20690
rect 19966 20638 20018 20690
rect 28030 20638 28082 20690
rect 28142 20638 28194 20690
rect 37662 20638 37714 20690
rect 41694 20638 41746 20690
rect 42142 20638 42194 20690
rect 44830 20638 44882 20690
rect 20190 20526 20242 20578
rect 22542 20526 22594 20578
rect 25678 20526 25730 20578
rect 26014 20526 26066 20578
rect 27806 20526 27858 20578
rect 36094 20526 36146 20578
rect 38222 20526 38274 20578
rect 38670 20526 38722 20578
rect 41134 20526 41186 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 17726 20190 17778 20242
rect 21198 20190 21250 20242
rect 22094 20190 22146 20242
rect 30158 20190 30210 20242
rect 31278 20190 31330 20242
rect 32286 20190 32338 20242
rect 33406 20190 33458 20242
rect 37886 20190 37938 20242
rect 9886 20078 9938 20130
rect 12798 20078 12850 20130
rect 14590 20078 14642 20130
rect 17950 20078 18002 20130
rect 21534 20078 21586 20130
rect 22318 20078 22370 20130
rect 24222 20078 24274 20130
rect 26014 20078 26066 20130
rect 27246 20078 27298 20130
rect 28590 20078 28642 20130
rect 29934 20078 29986 20130
rect 31502 20078 31554 20130
rect 32062 20078 32114 20130
rect 32398 20078 32450 20130
rect 35086 20078 35138 20130
rect 36430 20078 36482 20130
rect 38110 20078 38162 20130
rect 38670 20134 38722 20186
rect 41022 20190 41074 20242
rect 43262 20190 43314 20242
rect 45390 20190 45442 20242
rect 39790 20078 39842 20130
rect 45166 20078 45218 20130
rect 45502 20078 45554 20130
rect 47406 20078 47458 20130
rect 10558 19966 10610 20018
rect 11902 19966 11954 20018
rect 17278 19966 17330 20018
rect 19742 19966 19794 20018
rect 20414 19966 20466 20018
rect 21870 19966 21922 20018
rect 22766 19966 22818 20018
rect 23214 19966 23266 20018
rect 30270 19966 30322 20018
rect 30606 19966 30658 20018
rect 31390 19966 31442 20018
rect 31950 19966 32002 20018
rect 34302 19966 34354 20018
rect 35198 19966 35250 20018
rect 36206 19966 36258 20018
rect 36878 19966 36930 20018
rect 37102 19966 37154 20018
rect 38222 19966 38274 20018
rect 38782 19966 38834 20018
rect 39342 19966 39394 20018
rect 40238 19966 40290 20018
rect 42254 19966 42306 20018
rect 44382 19966 44434 20018
rect 44606 19966 44658 20018
rect 45054 19966 45106 20018
rect 47630 19966 47682 20018
rect 11118 19854 11170 19906
rect 12350 19854 12402 19906
rect 15150 19854 15202 19906
rect 17838 19854 17890 19906
rect 25230 19854 25282 19906
rect 27918 19854 27970 19906
rect 29038 19854 29090 19906
rect 30718 19854 30770 19906
rect 36318 19854 36370 19906
rect 37550 19854 37602 19906
rect 39902 19854 39954 19906
rect 41806 19854 41858 19906
rect 42702 19854 42754 19906
rect 43038 19854 43090 19906
rect 44494 19854 44546 19906
rect 47182 19854 47234 19906
rect 9998 19742 10050 19794
rect 13806 19742 13858 19794
rect 20302 19742 20354 19794
rect 22430 19742 22482 19794
rect 38670 19742 38722 19794
rect 43374 19742 43426 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14030 19406 14082 19458
rect 22766 19406 22818 19458
rect 37550 19406 37602 19458
rect 41582 19406 41634 19458
rect 15038 19294 15090 19346
rect 21534 19294 21586 19346
rect 23998 19294 24050 19346
rect 25566 19294 25618 19346
rect 32622 19294 32674 19346
rect 33742 19294 33794 19346
rect 34190 19294 34242 19346
rect 34750 19294 34802 19346
rect 35310 19294 35362 19346
rect 36206 19294 36258 19346
rect 37214 19294 37266 19346
rect 41022 19294 41074 19346
rect 45838 19294 45890 19346
rect 9774 19182 9826 19234
rect 10334 19182 10386 19234
rect 11230 19182 11282 19234
rect 11790 19182 11842 19234
rect 12014 19182 12066 19234
rect 12462 19182 12514 19234
rect 21982 19182 22034 19234
rect 22318 19182 22370 19234
rect 22542 19182 22594 19234
rect 23550 19182 23602 19234
rect 24894 19182 24946 19234
rect 25454 19182 25506 19234
rect 26126 19182 26178 19234
rect 33406 19182 33458 19234
rect 33630 19182 33682 19234
rect 33966 19182 34018 19234
rect 34526 19182 34578 19234
rect 35982 19182 36034 19234
rect 36990 19182 37042 19234
rect 38334 19182 38386 19234
rect 38670 19182 38722 19234
rect 39006 19182 39058 19234
rect 39678 19182 39730 19234
rect 40238 19182 40290 19234
rect 40910 19182 40962 19234
rect 44942 19182 44994 19234
rect 45390 19182 45442 19234
rect 47182 19182 47234 19234
rect 9886 19070 9938 19122
rect 11342 19070 11394 19122
rect 13470 19070 13522 19122
rect 13918 19070 13970 19122
rect 21758 19070 21810 19122
rect 39790 19070 39842 19122
rect 48078 19070 48130 19122
rect 9214 18958 9266 19010
rect 10446 18958 10498 19010
rect 11006 18958 11058 19010
rect 11454 18958 11506 19010
rect 12238 18958 12290 19010
rect 12574 18958 12626 19010
rect 12910 18958 12962 19010
rect 13694 18958 13746 19010
rect 22206 18958 22258 19010
rect 23102 18958 23154 19010
rect 38110 18958 38162 19010
rect 38222 18958 38274 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 9774 18622 9826 18674
rect 11230 18622 11282 18674
rect 15262 18622 15314 18674
rect 31950 18622 32002 18674
rect 33406 18622 33458 18674
rect 34862 18622 34914 18674
rect 36094 18622 36146 18674
rect 36318 18622 36370 18674
rect 38222 18622 38274 18674
rect 10670 18510 10722 18562
rect 11006 18510 11058 18562
rect 12238 18510 12290 18562
rect 14590 18510 14642 18562
rect 20974 18510 21026 18562
rect 29038 18510 29090 18562
rect 31726 18510 31778 18562
rect 36542 18510 36594 18562
rect 36654 18510 36706 18562
rect 38334 18566 38386 18618
rect 38782 18510 38834 18562
rect 40350 18510 40402 18562
rect 10110 18398 10162 18450
rect 10334 18398 10386 18450
rect 10558 18398 10610 18450
rect 12462 18398 12514 18450
rect 13246 18398 13298 18450
rect 14926 18398 14978 18450
rect 18510 18398 18562 18450
rect 20302 18398 20354 18450
rect 21758 18398 21810 18450
rect 22542 18398 22594 18450
rect 28814 18398 28866 18450
rect 32286 18398 32338 18450
rect 35534 18398 35586 18450
rect 35758 18398 35810 18450
rect 37662 18398 37714 18450
rect 38670 18398 38722 18450
rect 39006 18398 39058 18450
rect 39454 18398 39506 18450
rect 39902 18398 39954 18450
rect 15710 18286 15762 18338
rect 18734 18286 18786 18338
rect 19182 18286 19234 18338
rect 20078 18286 20130 18338
rect 21422 18286 21474 18338
rect 24670 18286 24722 18338
rect 25342 18286 25394 18338
rect 29934 18286 29986 18338
rect 31166 18286 31218 18338
rect 31838 18286 31890 18338
rect 33966 18286 34018 18338
rect 34414 18286 34466 18338
rect 37214 18286 37266 18338
rect 11342 18174 11394 18226
rect 15934 18174 15986 18226
rect 16270 18174 16322 18226
rect 33742 18174 33794 18226
rect 34414 18174 34466 18226
rect 34862 18174 34914 18226
rect 38222 18174 38274 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 18734 17838 18786 17890
rect 36094 17838 36146 17890
rect 11118 17726 11170 17778
rect 14590 17726 14642 17778
rect 26238 17726 26290 17778
rect 28366 17726 28418 17778
rect 29374 17726 29426 17778
rect 31278 17726 31330 17778
rect 31726 17726 31778 17778
rect 32398 17726 32450 17778
rect 34526 17726 34578 17778
rect 35422 17726 35474 17778
rect 37214 17726 37266 17778
rect 39678 17726 39730 17778
rect 40126 17726 40178 17778
rect 42142 17726 42194 17778
rect 13694 17614 13746 17666
rect 14366 17614 14418 17666
rect 15822 17614 15874 17666
rect 16718 17614 16770 17666
rect 18510 17614 18562 17666
rect 20302 17614 20354 17666
rect 20526 17614 20578 17666
rect 25118 17614 25170 17666
rect 25566 17614 25618 17666
rect 30270 17614 30322 17666
rect 34862 17614 34914 17666
rect 39006 17614 39058 17666
rect 39342 17614 39394 17666
rect 42030 17614 42082 17666
rect 14590 17502 14642 17554
rect 15598 17502 15650 17554
rect 17390 17502 17442 17554
rect 19070 17502 19122 17554
rect 19966 17502 20018 17554
rect 36206 17502 36258 17554
rect 37886 17502 37938 17554
rect 39118 17502 39170 17554
rect 42702 17502 42754 17554
rect 43038 17502 43090 17554
rect 43262 17502 43314 17554
rect 20414 17390 20466 17442
rect 29934 17390 29986 17442
rect 30382 17390 30434 17442
rect 30494 17390 30546 17442
rect 30718 17390 30770 17442
rect 31166 17390 31218 17442
rect 36094 17390 36146 17442
rect 38334 17390 38386 17442
rect 43150 17390 43202 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 13918 17054 13970 17106
rect 14814 17054 14866 17106
rect 16382 17054 16434 17106
rect 16606 17054 16658 17106
rect 21646 17054 21698 17106
rect 28590 17054 28642 17106
rect 32286 17054 32338 17106
rect 33630 17054 33682 17106
rect 34190 17054 34242 17106
rect 36542 17054 36594 17106
rect 38782 17054 38834 17106
rect 11118 16942 11170 16994
rect 11230 16942 11282 16994
rect 14254 16942 14306 16994
rect 14702 16942 14754 16994
rect 15038 16942 15090 16994
rect 21422 16942 21474 16994
rect 22206 16942 22258 16994
rect 33294 16942 33346 16994
rect 45726 16942 45778 16994
rect 11454 16830 11506 16882
rect 14142 16830 14194 16882
rect 14478 16830 14530 16882
rect 15262 16830 15314 16882
rect 15486 16830 15538 16882
rect 15822 16830 15874 16882
rect 16158 16830 16210 16882
rect 18734 16830 18786 16882
rect 21086 16830 21138 16882
rect 29934 16830 29986 16882
rect 30606 16830 30658 16882
rect 31838 16830 31890 16882
rect 32062 16830 32114 16882
rect 32398 16830 32450 16882
rect 41582 16830 41634 16882
rect 43262 16830 43314 16882
rect 45054 16830 45106 16882
rect 47070 16830 47122 16882
rect 47742 16830 47794 16882
rect 16270 16718 16322 16770
rect 18846 16718 18898 16770
rect 19182 16718 19234 16770
rect 29822 16718 29874 16770
rect 31278 16718 31330 16770
rect 41694 16718 41746 16770
rect 42142 16718 42194 16770
rect 43038 16718 43090 16770
rect 44942 16718 44994 16770
rect 21310 16606 21362 16658
rect 30270 16606 30322 16658
rect 43598 16606 43650 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 12350 16270 12402 16322
rect 24558 16270 24610 16322
rect 24894 16270 24946 16322
rect 32398 16270 32450 16322
rect 32958 16270 33010 16322
rect 43262 16270 43314 16322
rect 14702 16158 14754 16210
rect 15262 16158 15314 16210
rect 20190 16158 20242 16210
rect 20862 16158 20914 16210
rect 22094 16158 22146 16210
rect 23102 16158 23154 16210
rect 24446 16158 24498 16210
rect 24894 16158 24946 16210
rect 25902 16158 25954 16210
rect 28030 16158 28082 16210
rect 29374 16158 29426 16210
rect 31278 16158 31330 16210
rect 32510 16158 32562 16210
rect 36206 16158 36258 16210
rect 37102 16158 37154 16210
rect 42254 16158 42306 16210
rect 43038 16158 43090 16210
rect 45614 16158 45666 16210
rect 47070 16158 47122 16210
rect 10446 16046 10498 16098
rect 10670 16046 10722 16098
rect 11454 16046 11506 16098
rect 11566 16046 11618 16098
rect 11902 16046 11954 16098
rect 12238 16046 12290 16098
rect 14366 16046 14418 16098
rect 19966 16046 20018 16098
rect 21310 16046 21362 16098
rect 21982 16046 22034 16098
rect 25118 16046 25170 16098
rect 29710 16046 29762 16098
rect 29822 16046 29874 16098
rect 29934 16046 29986 16098
rect 30382 16046 30434 16098
rect 31166 16046 31218 16098
rect 32062 16046 32114 16098
rect 32846 16046 32898 16098
rect 42926 16046 42978 16098
rect 44830 16046 44882 16098
rect 47630 16046 47682 16098
rect 19294 15934 19346 15986
rect 22654 15934 22706 15986
rect 30718 15934 30770 15986
rect 41918 15934 41970 15986
rect 42142 15934 42194 15986
rect 42366 15934 42418 15986
rect 42814 15934 42866 15986
rect 45166 15934 45218 15986
rect 45502 15934 45554 15986
rect 47406 15934 47458 15986
rect 11006 15822 11058 15874
rect 11790 15822 11842 15874
rect 12350 15822 12402 15874
rect 23438 15822 23490 15874
rect 23774 15822 23826 15874
rect 45054 15822 45106 15874
rect 45726 15822 45778 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 12126 15486 12178 15538
rect 12350 15486 12402 15538
rect 12574 15486 12626 15538
rect 13134 15486 13186 15538
rect 21534 15486 21586 15538
rect 24334 15486 24386 15538
rect 25342 15486 25394 15538
rect 25790 15486 25842 15538
rect 30606 15486 30658 15538
rect 37550 15486 37602 15538
rect 11454 15374 11506 15426
rect 11566 15374 11618 15426
rect 11678 15374 11730 15426
rect 13022 15374 13074 15426
rect 16270 15374 16322 15426
rect 18398 15374 18450 15426
rect 22878 15374 22930 15426
rect 24446 15374 24498 15426
rect 35310 15374 35362 15426
rect 35758 15374 35810 15426
rect 35982 15374 36034 15426
rect 36542 15374 36594 15426
rect 36878 15374 36930 15426
rect 38446 15374 38498 15426
rect 40126 15374 40178 15426
rect 40350 15374 40402 15426
rect 13358 15262 13410 15314
rect 17726 15262 17778 15314
rect 21198 15262 21250 15314
rect 22766 15262 22818 15314
rect 24110 15262 24162 15314
rect 31166 15262 31218 15314
rect 31838 15262 31890 15314
rect 36094 15262 36146 15314
rect 37438 15262 37490 15314
rect 37774 15262 37826 15314
rect 12238 15150 12290 15202
rect 17950 15150 18002 15202
rect 26350 15150 26402 15202
rect 35422 15150 35474 15202
rect 38334 15150 38386 15202
rect 11006 15038 11058 15090
rect 22878 15038 22930 15090
rect 31950 15038 32002 15090
rect 35534 15038 35586 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 22430 14702 22482 14754
rect 43710 14702 43762 14754
rect 11566 14590 11618 14642
rect 12350 14590 12402 14642
rect 13470 14590 13522 14642
rect 14702 14590 14754 14642
rect 27470 14590 27522 14642
rect 29710 14590 29762 14642
rect 30158 14590 30210 14642
rect 31166 14590 31218 14642
rect 31614 14590 31666 14642
rect 32062 14590 32114 14642
rect 35870 14590 35922 14642
rect 36542 14590 36594 14642
rect 38334 14590 38386 14642
rect 40014 14590 40066 14642
rect 40462 14590 40514 14642
rect 40910 14590 40962 14642
rect 41806 14590 41858 14642
rect 44830 14590 44882 14642
rect 46734 14590 46786 14642
rect 11118 14478 11170 14530
rect 12574 14478 12626 14530
rect 13022 14478 13074 14530
rect 15710 14478 15762 14530
rect 17614 14478 17666 14530
rect 17838 14478 17890 14530
rect 21534 14478 21586 14530
rect 21758 14478 21810 14530
rect 22878 14478 22930 14530
rect 23326 14478 23378 14530
rect 27918 14478 27970 14530
rect 29150 14478 29202 14530
rect 30494 14478 30546 14530
rect 33294 14478 33346 14530
rect 35422 14478 35474 14530
rect 37214 14478 37266 14530
rect 38222 14478 38274 14530
rect 39118 14478 39170 14530
rect 39790 14478 39842 14530
rect 41134 14478 41186 14530
rect 43822 14478 43874 14530
rect 44046 14478 44098 14530
rect 44270 14478 44322 14530
rect 45054 14478 45106 14530
rect 45390 14478 45442 14530
rect 46958 14478 47010 14530
rect 13582 14366 13634 14418
rect 15374 14366 15426 14418
rect 16046 14366 16098 14418
rect 16494 14366 16546 14418
rect 16606 14366 16658 14418
rect 21422 14366 21474 14418
rect 22318 14366 22370 14418
rect 22654 14366 22706 14418
rect 26574 14366 26626 14418
rect 26910 14366 26962 14418
rect 30606 14366 30658 14418
rect 32734 14366 32786 14418
rect 34414 14366 34466 14418
rect 34974 14366 35026 14418
rect 37102 14366 37154 14418
rect 48078 14366 48130 14418
rect 16270 14254 16322 14306
rect 17390 14254 17442 14306
rect 17726 14254 17778 14306
rect 21198 14254 21250 14306
rect 22094 14254 22146 14306
rect 30830 14254 30882 14306
rect 34302 14254 34354 14306
rect 36878 14254 36930 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 14926 13918 14978 13970
rect 16494 13918 16546 13970
rect 18734 13918 18786 13970
rect 22878 13918 22930 13970
rect 23438 13918 23490 13970
rect 23998 13918 24050 13970
rect 32286 13918 32338 13970
rect 37102 13918 37154 13970
rect 37662 13918 37714 13970
rect 38222 13918 38274 13970
rect 45390 13918 45442 13970
rect 12014 13806 12066 13858
rect 12686 13806 12738 13858
rect 14814 13806 14866 13858
rect 15150 13806 15202 13858
rect 16606 13806 16658 13858
rect 18846 13806 18898 13858
rect 22766 13806 22818 13858
rect 30494 13806 30546 13858
rect 34750 13806 34802 13858
rect 36318 13806 36370 13858
rect 37214 13806 37266 13858
rect 37550 13806 37602 13858
rect 38110 13806 38162 13858
rect 43822 13806 43874 13858
rect 11790 13694 11842 13746
rect 13246 13694 13298 13746
rect 14254 13694 14306 13746
rect 15486 13694 15538 13746
rect 15822 13694 15874 13746
rect 16046 13694 16098 13746
rect 16270 13694 16322 13746
rect 20078 13694 20130 13746
rect 20638 13694 20690 13746
rect 21086 13694 21138 13746
rect 22206 13694 22258 13746
rect 22542 13694 22594 13746
rect 23550 13694 23602 13746
rect 24110 13694 24162 13746
rect 25230 13694 25282 13746
rect 25678 13694 25730 13746
rect 27134 13694 27186 13746
rect 29710 13694 29762 13746
rect 30158 13694 30210 13746
rect 31838 13694 31890 13746
rect 35198 13694 35250 13746
rect 36654 13694 36706 13746
rect 36878 13694 36930 13746
rect 38446 13694 38498 13746
rect 38782 13694 38834 13746
rect 39678 13694 39730 13746
rect 44046 13694 44098 13746
rect 45054 13694 45106 13746
rect 11902 13582 11954 13634
rect 14478 13582 14530 13634
rect 15934 13582 15986 13634
rect 19518 13582 19570 13634
rect 21198 13582 21250 13634
rect 24446 13582 24498 13634
rect 35534 13582 35586 13634
rect 13918 13470 13970 13522
rect 18734 13470 18786 13522
rect 19294 13470 19346 13522
rect 23438 13470 23490 13522
rect 25902 13470 25954 13522
rect 29374 13470 29426 13522
rect 31278 13470 31330 13522
rect 31614 13470 31666 13522
rect 37662 13470 37714 13522
rect 39006 13470 39058 13522
rect 39342 13470 39394 13522
rect 39902 13470 39954 13522
rect 40238 13470 40290 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 18958 13134 19010 13186
rect 14702 13022 14754 13074
rect 15934 13022 15986 13074
rect 17054 13022 17106 13074
rect 20078 13022 20130 13074
rect 24446 13022 24498 13074
rect 25566 13022 25618 13074
rect 26014 13022 26066 13074
rect 29374 13022 29426 13074
rect 30606 13022 30658 13074
rect 32398 13022 32450 13074
rect 37102 13022 37154 13074
rect 41246 13022 41298 13074
rect 43262 13022 43314 13074
rect 12238 12910 12290 12962
rect 13694 12910 13746 12962
rect 14366 12910 14418 12962
rect 14814 12910 14866 12962
rect 16606 12910 16658 12962
rect 19406 12910 19458 12962
rect 24558 12910 24610 12962
rect 29710 12910 29762 12962
rect 30830 12910 30882 12962
rect 32174 12910 32226 12962
rect 34750 12910 34802 12962
rect 34974 12910 35026 12962
rect 35310 12910 35362 12962
rect 36206 12910 36258 12962
rect 39790 12910 39842 12962
rect 40014 12910 40066 12962
rect 40350 12910 40402 12962
rect 42590 12910 42642 12962
rect 13582 12798 13634 12850
rect 15374 12798 15426 12850
rect 16158 12798 16210 12850
rect 19070 12798 19122 12850
rect 30158 12798 30210 12850
rect 31502 12798 31554 12850
rect 32846 12798 32898 12850
rect 36094 12798 36146 12850
rect 39902 12798 39954 12850
rect 41694 12798 41746 12850
rect 12574 12686 12626 12738
rect 13358 12686 13410 12738
rect 18958 12686 19010 12738
rect 19518 12686 19570 12738
rect 19742 12686 19794 12738
rect 34974 12686 35026 12738
rect 35870 12686 35922 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 14030 12350 14082 12402
rect 15934 12350 15986 12402
rect 16046 12350 16098 12402
rect 16606 12350 16658 12402
rect 20414 12350 20466 12402
rect 25454 12350 25506 12402
rect 26350 12350 26402 12402
rect 26910 12350 26962 12402
rect 27582 12350 27634 12402
rect 28142 12350 28194 12402
rect 31278 12350 31330 12402
rect 36542 12350 36594 12402
rect 12350 12238 12402 12290
rect 19070 12238 19122 12290
rect 19406 12238 19458 12290
rect 25342 12238 25394 12290
rect 27806 12238 27858 12290
rect 31838 12238 31890 12290
rect 33182 12238 33234 12290
rect 41022 12238 41074 12290
rect 12686 12126 12738 12178
rect 14702 12126 14754 12178
rect 15150 12126 15202 12178
rect 15486 12126 15538 12178
rect 16158 12126 16210 12178
rect 18174 12126 18226 12178
rect 19630 12126 19682 12178
rect 25678 12126 25730 12178
rect 26238 12126 26290 12178
rect 26574 12126 26626 12178
rect 27470 12126 27522 12178
rect 31614 12126 31666 12178
rect 33294 12126 33346 12178
rect 43374 12126 43426 12178
rect 43822 12126 43874 12178
rect 46734 12126 46786 12178
rect 46958 12126 47010 12178
rect 14254 12014 14306 12066
rect 18734 12014 18786 12066
rect 41134 12014 41186 12066
rect 41470 12014 41522 12066
rect 42366 12014 42418 12066
rect 12686 11902 12738 11954
rect 19966 11902 20018 11954
rect 33182 11902 33234 11954
rect 41694 11902 41746 11954
rect 42030 11902 42082 11954
rect 42590 11902 42642 11954
rect 42926 11902 42978 11954
rect 43374 11902 43426 11954
rect 47742 11902 47794 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 15150 11566 15202 11618
rect 15038 11454 15090 11506
rect 24334 11454 24386 11506
rect 25678 11454 25730 11506
rect 27134 11454 27186 11506
rect 29822 11454 29874 11506
rect 11230 11342 11282 11394
rect 11566 11342 11618 11394
rect 11790 11342 11842 11394
rect 12686 11342 12738 11394
rect 14702 11342 14754 11394
rect 18734 11342 18786 11394
rect 19406 11342 19458 11394
rect 22766 11342 22818 11394
rect 23214 11342 23266 11394
rect 24670 11342 24722 11394
rect 25902 11342 25954 11394
rect 26910 11342 26962 11394
rect 27582 11342 27634 11394
rect 28142 11342 28194 11394
rect 29150 11342 29202 11394
rect 32286 11342 32338 11394
rect 32846 11342 32898 11394
rect 32958 11342 33010 11394
rect 33742 11342 33794 11394
rect 34190 11342 34242 11394
rect 37326 11342 37378 11394
rect 37774 11342 37826 11394
rect 41918 11342 41970 11394
rect 42254 11342 42306 11394
rect 42478 11342 42530 11394
rect 11342 11230 11394 11282
rect 12238 11230 12290 11282
rect 25006 11230 25058 11282
rect 28030 11230 28082 11282
rect 28590 11230 28642 11282
rect 29262 11230 29314 11282
rect 30270 11230 30322 11282
rect 33294 11230 33346 11282
rect 36206 11230 36258 11282
rect 36318 11230 36370 11282
rect 12798 11118 12850 11170
rect 18846 11118 18898 11170
rect 18958 11118 19010 11170
rect 26238 11118 26290 11170
rect 27806 11118 27858 11170
rect 29486 11118 29538 11170
rect 36542 11118 36594 11170
rect 42142 11118 42194 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 23662 10782 23714 10834
rect 24558 10782 24610 10834
rect 24782 10782 24834 10834
rect 26798 10782 26850 10834
rect 26910 10782 26962 10834
rect 30046 10782 30098 10834
rect 34190 10782 34242 10834
rect 12126 10670 12178 10722
rect 21534 10670 21586 10722
rect 23214 10670 23266 10722
rect 23774 10670 23826 10722
rect 24446 10670 24498 10722
rect 28478 10670 28530 10722
rect 32286 10670 32338 10722
rect 32398 10670 32450 10722
rect 32622 10670 32674 10722
rect 33182 10670 33234 10722
rect 33294 10670 33346 10722
rect 35646 10670 35698 10722
rect 44382 10670 44434 10722
rect 12350 10558 12402 10610
rect 13022 10558 13074 10610
rect 17950 10558 18002 10610
rect 18622 10558 18674 10610
rect 19630 10558 19682 10610
rect 20078 10558 20130 10610
rect 20862 10558 20914 10610
rect 22206 10558 22258 10610
rect 22878 10558 22930 10610
rect 25790 10558 25842 10610
rect 27022 10558 27074 10610
rect 27358 10558 27410 10610
rect 29598 10558 29650 10610
rect 34750 10558 34802 10610
rect 35422 10558 35474 10610
rect 37550 10558 37602 10610
rect 39006 10558 39058 10610
rect 43262 10558 43314 10610
rect 43486 10558 43538 10610
rect 44046 10558 44098 10610
rect 13694 10446 13746 10498
rect 17726 10446 17778 10498
rect 19182 10446 19234 10498
rect 20750 10446 20802 10498
rect 22766 10446 22818 10498
rect 26014 10446 26066 10498
rect 26462 10446 26514 10498
rect 28142 10446 28194 10498
rect 36766 10446 36818 10498
rect 37998 10446 38050 10498
rect 23662 10334 23714 10386
rect 33182 10334 33234 10386
rect 39230 10334 39282 10386
rect 43150 10334 43202 10386
rect 43598 10334 43650 10386
rect 44046 10334 44098 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 21870 9998 21922 10050
rect 22206 9998 22258 10050
rect 26126 9998 26178 10050
rect 26462 9998 26514 10050
rect 16270 9886 16322 9938
rect 17166 9886 17218 9938
rect 18174 9886 18226 9938
rect 25006 9886 25058 9938
rect 25902 9886 25954 9938
rect 31278 9886 31330 9938
rect 31838 9886 31890 9938
rect 34190 9886 34242 9938
rect 34862 9886 34914 9938
rect 39230 9886 39282 9938
rect 44270 9886 44322 9938
rect 46734 9886 46786 9938
rect 14366 9774 14418 9826
rect 15598 9774 15650 9826
rect 16606 9774 16658 9826
rect 18398 9774 18450 9826
rect 19854 9774 19906 9826
rect 20190 9774 20242 9826
rect 26910 9774 26962 9826
rect 29822 9774 29874 9826
rect 34974 9774 35026 9826
rect 37998 9774 38050 9826
rect 38670 9774 38722 9826
rect 40798 9774 40850 9826
rect 42142 9774 42194 9826
rect 42814 9774 42866 9826
rect 43486 9774 43538 9826
rect 46958 9774 47010 9826
rect 14590 9662 14642 9714
rect 15822 9662 15874 9714
rect 18734 9662 18786 9714
rect 19630 9662 19682 9714
rect 21646 9662 21698 9714
rect 27022 9662 27074 9714
rect 27582 9662 27634 9714
rect 30718 9662 30770 9714
rect 34526 9662 34578 9714
rect 37438 9662 37490 9714
rect 38110 9662 38162 9714
rect 38334 9662 38386 9714
rect 39342 9662 39394 9714
rect 48078 9662 48130 9714
rect 15486 9550 15538 9602
rect 20078 9550 20130 9602
rect 27246 9550 27298 9602
rect 29486 9550 29538 9602
rect 31726 9550 31778 9602
rect 40910 9550 40962 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 31278 9214 31330 9266
rect 31390 9214 31442 9266
rect 38670 9214 38722 9266
rect 42926 9214 42978 9266
rect 43934 9214 43986 9266
rect 44158 9214 44210 9266
rect 14366 9102 14418 9154
rect 14926 9102 14978 9154
rect 15710 9102 15762 9154
rect 31166 9102 31218 9154
rect 34750 9102 34802 9154
rect 13918 8990 13970 9042
rect 14254 8990 14306 9042
rect 15038 8990 15090 9042
rect 15598 8990 15650 9042
rect 31838 8990 31890 9042
rect 35086 8990 35138 9042
rect 37214 8990 37266 9042
rect 37662 8990 37714 9042
rect 38446 8990 38498 9042
rect 42702 8990 42754 9042
rect 43374 8990 43426 9042
rect 43486 8990 43538 9042
rect 44046 8990 44098 9042
rect 15934 8878 15986 8930
rect 34862 8878 34914 8930
rect 38110 8878 38162 8930
rect 42814 8878 42866 8930
rect 38782 8766 38834 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 35086 8430 35138 8482
rect 15150 8318 15202 8370
rect 16606 8318 16658 8370
rect 18062 8318 18114 8370
rect 18734 8318 18786 8370
rect 20750 8318 20802 8370
rect 21870 8318 21922 8370
rect 23550 8318 23602 8370
rect 31726 8318 31778 8370
rect 41694 8318 41746 8370
rect 14814 8206 14866 8258
rect 15710 8206 15762 8258
rect 16494 8206 16546 8258
rect 17726 8206 17778 8258
rect 18622 8206 18674 8258
rect 21758 8206 21810 8258
rect 22318 8206 22370 8258
rect 23774 8206 23826 8258
rect 27358 8206 27410 8258
rect 31502 8206 31554 8258
rect 34190 8206 34242 8258
rect 34750 8206 34802 8258
rect 35086 8206 35138 8258
rect 40126 8206 40178 8258
rect 17390 8094 17442 8146
rect 17950 8094 18002 8146
rect 19518 8094 19570 8146
rect 20414 8094 20466 8146
rect 32174 8094 32226 8146
rect 34526 8094 34578 8146
rect 35422 8094 35474 8146
rect 41134 8094 41186 8146
rect 20638 7982 20690 8034
rect 24110 7982 24162 8034
rect 27806 7982 27858 8034
rect 27918 7982 27970 8034
rect 28030 7982 28082 8034
rect 34638 7982 34690 8034
rect 39902 7982 39954 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 18398 7646 18450 7698
rect 28702 7646 28754 7698
rect 31838 7646 31890 7698
rect 33406 7646 33458 7698
rect 33518 7646 33570 7698
rect 42030 7646 42082 7698
rect 42142 7646 42194 7698
rect 18622 7534 18674 7586
rect 20974 7534 21026 7586
rect 21310 7534 21362 7586
rect 21870 7534 21922 7586
rect 26350 7534 26402 7586
rect 32062 7534 32114 7586
rect 20302 7422 20354 7474
rect 21646 7422 21698 7474
rect 23774 7422 23826 7474
rect 25230 7422 25282 7474
rect 25790 7422 25842 7474
rect 26910 7422 26962 7474
rect 27358 7422 27410 7474
rect 28142 7422 28194 7474
rect 28366 7422 28418 7474
rect 32174 7422 32226 7474
rect 32958 7422 33010 7474
rect 33630 7422 33682 7474
rect 41470 7422 41522 7474
rect 41918 7422 41970 7474
rect 18398 7310 18450 7362
rect 20526 7310 20578 7362
rect 21758 7310 21810 7362
rect 23886 7310 23938 7362
rect 25678 7310 25730 7362
rect 27806 7310 27858 7362
rect 24558 7198 24610 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 13694 6862 13746 6914
rect 23998 6862 24050 6914
rect 27246 6862 27298 6914
rect 27582 6862 27634 6914
rect 23774 6750 23826 6802
rect 26574 6750 26626 6802
rect 27806 6750 27858 6802
rect 33854 6750 33906 6802
rect 34526 6750 34578 6802
rect 39566 6750 39618 6802
rect 13470 6638 13522 6690
rect 15934 6638 15986 6690
rect 16382 6638 16434 6690
rect 18174 6638 18226 6690
rect 18734 6638 18786 6690
rect 24334 6638 24386 6690
rect 29710 6638 29762 6690
rect 30158 6638 30210 6690
rect 31278 6638 31330 6690
rect 31614 6638 31666 6690
rect 31838 6638 31890 6690
rect 32398 6638 32450 6690
rect 34414 6638 34466 6690
rect 37662 6638 37714 6690
rect 38558 6638 38610 6690
rect 41134 6638 41186 6690
rect 42254 6638 42306 6690
rect 42590 6638 42642 6690
rect 46734 6638 46786 6690
rect 46958 6638 47010 6690
rect 31390 6526 31442 6578
rect 33406 6526 33458 6578
rect 34638 6526 34690 6578
rect 35310 6526 35362 6578
rect 35646 6526 35698 6578
rect 35870 6526 35922 6578
rect 37326 6526 37378 6578
rect 39902 6526 39954 6578
rect 41470 6526 41522 6578
rect 42142 6526 42194 6578
rect 48078 6526 48130 6578
rect 14030 6414 14082 6466
rect 15710 6414 15762 6466
rect 15822 6414 15874 6466
rect 18510 6414 18562 6466
rect 18622 6414 18674 6466
rect 29598 6414 29650 6466
rect 29822 6414 29874 6466
rect 35422 6414 35474 6466
rect 36430 6414 36482 6466
rect 38894 6414 38946 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 16494 6078 16546 6130
rect 20302 6078 20354 6130
rect 30270 6078 30322 6130
rect 33182 6078 33234 6130
rect 35534 6078 35586 6130
rect 38894 6078 38946 6130
rect 39566 6078 39618 6130
rect 41358 6078 41410 6130
rect 13582 5966 13634 6018
rect 16718 5966 16770 6018
rect 16830 5966 16882 6018
rect 18398 5966 18450 6018
rect 20862 5966 20914 6018
rect 26238 5966 26290 6018
rect 28702 5966 28754 6018
rect 32510 5966 32562 6018
rect 33854 5966 33906 6018
rect 39118 5966 39170 6018
rect 41582 5966 41634 6018
rect 43038 5966 43090 6018
rect 13470 5854 13522 5906
rect 14254 5854 14306 5906
rect 15598 5854 15650 5906
rect 16270 5854 16322 5906
rect 17726 5854 17778 5906
rect 18734 5854 18786 5906
rect 18958 5854 19010 5906
rect 19182 5854 19234 5906
rect 20414 5854 20466 5906
rect 20638 5854 20690 5906
rect 20974 5854 21026 5906
rect 22318 5854 22370 5906
rect 22878 5854 22930 5906
rect 25678 5854 25730 5906
rect 29262 5854 29314 5906
rect 29934 5854 29986 5906
rect 31950 5854 32002 5906
rect 35310 5854 35362 5906
rect 36094 5854 36146 5906
rect 36654 5854 36706 5906
rect 37550 5854 37602 5906
rect 37886 5854 37938 5906
rect 39342 5854 39394 5906
rect 39678 5854 39730 5906
rect 41694 5854 41746 5906
rect 42142 5854 42194 5906
rect 42366 5854 42418 5906
rect 15822 5742 15874 5794
rect 17614 5742 17666 5794
rect 22990 5742 23042 5794
rect 25342 5742 25394 5794
rect 32174 5742 32226 5794
rect 33630 5742 33682 5794
rect 36878 5742 36930 5794
rect 37438 5742 37490 5794
rect 14590 5630 14642 5682
rect 19630 5630 19682 5682
rect 20302 5630 20354 5682
rect 38782 5630 38834 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 18958 5294 19010 5346
rect 25006 5294 25058 5346
rect 34974 5294 35026 5346
rect 14590 5182 14642 5234
rect 15038 5182 15090 5234
rect 15934 5182 15986 5234
rect 18734 5182 18786 5234
rect 20526 5182 20578 5234
rect 21534 5182 21586 5234
rect 23102 5182 23154 5234
rect 26014 5182 26066 5234
rect 29486 5182 29538 5234
rect 35534 5182 35586 5234
rect 37214 5182 37266 5234
rect 38894 5182 38946 5234
rect 40910 5182 40962 5234
rect 46622 5182 46674 5234
rect 14366 5070 14418 5122
rect 17278 5070 17330 5122
rect 19294 5070 19346 5122
rect 19854 5070 19906 5122
rect 20750 5070 20802 5122
rect 21758 5070 21810 5122
rect 22430 5070 22482 5122
rect 23326 5070 23378 5122
rect 24334 5070 24386 5122
rect 27582 5070 27634 5122
rect 30606 5070 30658 5122
rect 31502 5070 31554 5122
rect 35646 5070 35698 5122
rect 37774 5070 37826 5122
rect 37998 5070 38050 5122
rect 38334 5070 38386 5122
rect 40462 5070 40514 5122
rect 46958 5070 47010 5122
rect 47742 5070 47794 5122
rect 16158 4958 16210 5010
rect 17950 4958 18002 5010
rect 26126 4958 26178 5010
rect 28030 4958 28082 5010
rect 29374 4958 29426 5010
rect 29598 4958 29650 5010
rect 30382 4958 30434 5010
rect 38110 4958 38162 5010
rect 39006 4958 39058 5010
rect 31950 4846 32002 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19742 4510 19794 4562
rect 23662 4510 23714 4562
rect 23774 4510 23826 4562
rect 30046 4510 30098 4562
rect 35982 4510 36034 4562
rect 38670 4510 38722 4562
rect 38894 4510 38946 4562
rect 39566 4510 39618 4562
rect 14702 4398 14754 4450
rect 22094 4398 22146 4450
rect 25902 4398 25954 4450
rect 29934 4398 29986 4450
rect 30494 4398 30546 4450
rect 35870 4398 35922 4450
rect 46622 4398 46674 4450
rect 14030 4286 14082 4338
rect 14366 4286 14418 4338
rect 22318 4286 22370 4338
rect 23102 4286 23154 4338
rect 23550 4286 23602 4338
rect 27022 4286 27074 4338
rect 27470 4286 27522 4338
rect 30606 4286 30658 4338
rect 38782 4286 38834 4338
rect 39230 4286 39282 4338
rect 39678 4286 39730 4338
rect 46958 4286 47010 4338
rect 13470 4174 13522 4226
rect 18958 4174 19010 4226
rect 19182 4174 19234 4226
rect 22654 4174 22706 4226
rect 25342 4174 25394 4226
rect 48078 4174 48130 4226
rect 13694 4062 13746 4114
rect 19406 4062 19458 4114
rect 30046 4062 30098 4114
rect 36094 4062 36146 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 22990 3614 23042 3666
rect 40238 3614 40290 3666
rect 44046 3614 44098 3666
rect 45278 3614 45330 3666
rect 26910 3502 26962 3554
rect 27358 3502 27410 3554
rect 31390 3502 31442 3554
rect 45614 3502 45666 3554
rect 2718 3390 2770 3442
rect 2942 3390 2994 3442
rect 3278 3390 3330 3442
rect 6750 3390 6802 3442
rect 6974 3390 7026 3442
rect 7310 3390 7362 3442
rect 10782 3390 10834 3442
rect 11006 3390 11058 3442
rect 11342 3390 11394 3442
rect 14814 3390 14866 3442
rect 15038 3390 15090 3442
rect 15374 3390 15426 3442
rect 18846 3390 18898 3442
rect 19070 3390 19122 3442
rect 19406 3390 19458 3442
rect 23438 3390 23490 3442
rect 23886 3390 23938 3442
rect 28478 3390 28530 3442
rect 30942 3390 30994 3442
rect 39342 3390 39394 3442
rect 39790 3390 39842 3442
rect 43150 3390 43202 3442
rect 43598 3390 43650 3442
rect 46398 3390 46450 3442
rect 31166 3278 31218 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 2464 79200 2576 80000
rect 4256 79200 4368 80000
rect 6048 79200 6160 80000
rect 7840 79200 7952 80000
rect 9632 79200 9744 80000
rect 11424 79200 11536 80000
rect 13216 79200 13328 80000
rect 15008 79200 15120 80000
rect 16800 79200 16912 80000
rect 18592 79200 18704 80000
rect 20384 79200 20496 80000
rect 22176 79200 22288 80000
rect 23968 79200 24080 80000
rect 25760 79200 25872 80000
rect 27552 79200 27664 80000
rect 29344 79200 29456 80000
rect 31136 79200 31248 80000
rect 32928 79200 33040 80000
rect 34720 79200 34832 80000
rect 36512 79200 36624 80000
rect 38304 79200 38416 80000
rect 40096 79200 40208 80000
rect 41888 79200 42000 80000
rect 43680 79200 43792 80000
rect 45472 79200 45584 80000
rect 47264 79200 47376 80000
rect 2492 76578 2548 79200
rect 2492 76526 2494 76578
rect 2546 76526 2548 76578
rect 2492 76514 2548 76526
rect 2604 78036 2660 78046
rect 1932 76468 1988 76478
rect 1708 75572 1764 75582
rect 1708 74228 1764 75516
rect 1932 74786 1988 76412
rect 2604 75796 2660 77980
rect 2604 75682 2660 75740
rect 3276 76466 3332 76478
rect 3276 76414 3278 76466
rect 3330 76414 3332 76466
rect 2604 75630 2606 75682
rect 2658 75630 2660 75682
rect 2604 75618 2660 75630
rect 3164 75684 3220 75694
rect 3164 75590 3220 75628
rect 2268 75572 2324 75582
rect 1932 74734 1934 74786
rect 1986 74734 1988 74786
rect 1932 74722 1988 74734
rect 2156 75570 2324 75572
rect 2156 75518 2270 75570
rect 2322 75518 2324 75570
rect 2156 75516 2324 75518
rect 1820 74228 1876 74238
rect 1708 74226 1876 74228
rect 1708 74174 1822 74226
rect 1874 74174 1876 74226
rect 1708 74172 1876 74174
rect 1820 74162 1876 74172
rect 1708 73330 1764 73342
rect 1708 73278 1710 73330
rect 1762 73278 1764 73330
rect 1708 73108 1764 73278
rect 1764 73052 1876 73108
rect 1708 73042 1764 73052
rect 1820 72658 1876 73052
rect 1820 72606 1822 72658
rect 1874 72606 1876 72658
rect 1820 72594 1876 72606
rect 1260 72436 1316 72446
rect 1148 48132 1204 48142
rect 1148 20244 1204 48076
rect 1260 21700 1316 72380
rect 2156 71540 2212 75516
rect 2268 75506 2324 75516
rect 3276 73332 3332 76414
rect 3724 76468 3780 76478
rect 3724 76374 3780 76412
rect 4284 76356 4340 79200
rect 4396 76356 4452 76366
rect 4284 76354 4452 76356
rect 4284 76302 4398 76354
rect 4450 76302 4452 76354
rect 4284 76300 4452 76302
rect 6076 76356 6132 79200
rect 7868 76578 7924 79200
rect 9660 77700 9716 79200
rect 9660 77644 10052 77700
rect 9996 77252 10052 77644
rect 9996 77196 10276 77252
rect 10220 76690 10276 77196
rect 10220 76638 10222 76690
rect 10274 76638 10276 76690
rect 10220 76626 10276 76638
rect 11452 76692 11508 79200
rect 11788 76692 11844 76702
rect 11452 76690 11844 76692
rect 11452 76638 11790 76690
rect 11842 76638 11844 76690
rect 11452 76636 11844 76638
rect 11788 76626 11844 76636
rect 13244 76692 13300 79200
rect 15036 77252 15092 79200
rect 15036 77196 15652 77252
rect 13244 76626 13300 76636
rect 13916 76692 13972 76702
rect 7868 76526 7870 76578
rect 7922 76526 7924 76578
rect 7868 76514 7924 76526
rect 6972 76466 7028 76478
rect 6972 76414 6974 76466
rect 7026 76414 7028 76466
rect 6188 76356 6244 76366
rect 6076 76354 6244 76356
rect 6076 76302 6190 76354
rect 6242 76302 6244 76354
rect 6076 76300 6244 76302
rect 4396 76290 4452 76300
rect 6188 76290 6244 76300
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 3612 75796 3668 75806
rect 3612 75702 3668 75740
rect 5180 75684 5236 75694
rect 4060 75068 4340 75124
rect 4060 75010 4116 75068
rect 4060 74958 4062 75010
rect 4114 74958 4116 75010
rect 4060 74946 4116 74958
rect 4172 74900 4228 74910
rect 3948 74114 4004 74126
rect 4172 74116 4228 74844
rect 3948 74062 3950 74114
rect 4002 74062 4004 74114
rect 3388 74004 3444 74014
rect 3948 74004 4004 74062
rect 3388 74002 3948 74004
rect 3388 73950 3390 74002
rect 3442 73950 3948 74002
rect 3388 73948 3948 73950
rect 3388 73938 3444 73948
rect 3276 73276 3444 73332
rect 2268 73220 2324 73230
rect 2268 73218 3332 73220
rect 2268 73166 2270 73218
rect 2322 73166 3332 73218
rect 2268 73164 3332 73166
rect 2268 73154 2324 73164
rect 2156 71474 2212 71484
rect 2268 70868 2324 70878
rect 2156 70866 2324 70868
rect 2156 70814 2270 70866
rect 2322 70814 2324 70866
rect 2156 70812 2324 70814
rect 1708 70754 1764 70766
rect 1708 70702 1710 70754
rect 1762 70702 1764 70754
rect 1708 70644 1764 70702
rect 1764 70588 1876 70644
rect 1708 70578 1764 70588
rect 1820 70418 1876 70588
rect 1820 70366 1822 70418
rect 1874 70366 1876 70418
rect 1820 70354 1876 70366
rect 1820 68626 1876 68638
rect 1820 68574 1822 68626
rect 1874 68574 1876 68626
rect 1820 68180 1876 68574
rect 1820 67954 1876 68124
rect 1820 67902 1822 67954
rect 1874 67902 1876 67954
rect 1820 67890 1876 67902
rect 1596 66276 1652 66286
rect 1484 62468 1540 62478
rect 1372 56980 1428 56990
rect 1372 36708 1428 56924
rect 1484 46900 1540 62412
rect 1596 60452 1652 66220
rect 1820 66274 1876 66286
rect 1820 66222 1822 66274
rect 1874 66222 1876 66274
rect 1820 65716 1876 66222
rect 1820 65622 1876 65660
rect 2156 65604 2212 70812
rect 2268 70802 2324 70812
rect 2268 68514 2324 68526
rect 2268 68462 2270 68514
rect 2322 68462 2324 68514
rect 2268 67228 2324 68462
rect 2268 67172 2660 67228
rect 2268 66276 2324 66286
rect 2268 66182 2324 66220
rect 2156 65538 2212 65548
rect 1820 63922 1876 63934
rect 1820 63870 1822 63922
rect 1874 63870 1876 63922
rect 1820 63252 1876 63870
rect 2268 63924 2324 63934
rect 2268 63922 2436 63924
rect 2268 63870 2270 63922
rect 2322 63870 2436 63922
rect 2268 63868 2436 63870
rect 2268 63858 2324 63868
rect 1820 63158 1876 63196
rect 2268 62692 2324 62702
rect 2268 62188 2324 62636
rect 2156 62132 2324 62188
rect 2156 61570 2212 62132
rect 2156 61518 2158 61570
rect 2210 61518 2212 61570
rect 1596 60386 1652 60396
rect 1708 60788 1764 60798
rect 1708 60116 1764 60732
rect 1820 60116 1876 60126
rect 1708 60114 1876 60116
rect 1708 60062 1822 60114
rect 1874 60062 1876 60114
rect 1708 60060 1876 60062
rect 1820 60050 1876 60060
rect 1708 58324 1764 58334
rect 1708 58230 1764 58268
rect 2044 58210 2100 58222
rect 2044 58158 2046 58210
rect 2098 58158 2100 58210
rect 2044 57092 2100 58158
rect 2044 57026 2100 57036
rect 1932 56868 1988 56878
rect 2156 56868 2212 61518
rect 1820 56866 2212 56868
rect 1820 56814 1934 56866
rect 1986 56814 2212 56866
rect 1820 56812 2212 56814
rect 2268 60674 2324 60686
rect 2268 60622 2270 60674
rect 2322 60622 2324 60674
rect 1708 56082 1764 56094
rect 1708 56030 1710 56082
rect 1762 56030 1764 56082
rect 1708 55860 1764 56030
rect 1708 55794 1764 55804
rect 1708 54626 1764 54638
rect 1708 54574 1710 54626
rect 1762 54574 1764 54626
rect 1708 52948 1764 54574
rect 1820 53732 1876 56812
rect 1932 56802 1988 56812
rect 2044 56194 2100 56206
rect 2044 56142 2046 56194
rect 2098 56142 2100 56194
rect 1932 54514 1988 54526
rect 1932 54462 1934 54514
rect 1986 54462 1988 54514
rect 1932 54404 1988 54462
rect 1932 54338 1988 54348
rect 1820 53638 1876 53676
rect 2044 53284 2100 56142
rect 1708 52854 1764 52892
rect 1820 53228 2100 53284
rect 1820 49924 1876 53228
rect 2268 52836 2324 60622
rect 2380 56196 2436 63868
rect 2492 58324 2548 58334
rect 2492 58230 2548 58268
rect 2604 56308 2660 67172
rect 2940 61460 2996 61470
rect 2940 61366 2996 61404
rect 3164 57764 3220 57774
rect 2716 57762 3220 57764
rect 2716 57710 3166 57762
rect 3218 57710 3220 57762
rect 2716 57708 3220 57710
rect 2716 56978 2772 57708
rect 3164 57698 3220 57708
rect 2828 57092 2884 57102
rect 2884 57036 3108 57092
rect 2828 57026 2884 57036
rect 2716 56926 2718 56978
rect 2770 56926 2772 56978
rect 2716 56914 2772 56926
rect 2604 56252 2996 56308
rect 2380 56140 2660 56196
rect 2492 55970 2548 55982
rect 2492 55918 2494 55970
rect 2546 55918 2548 55970
rect 2492 55860 2548 55918
rect 2492 55794 2548 55804
rect 2492 54404 2548 54414
rect 2492 54310 2548 54348
rect 2492 53620 2548 53630
rect 2268 52770 2324 52780
rect 2380 53618 2548 53620
rect 2380 53566 2494 53618
rect 2546 53566 2548 53618
rect 2380 53564 2548 53566
rect 2380 52050 2436 53564
rect 2492 53554 2548 53564
rect 2380 51998 2382 52050
rect 2434 51998 2436 52050
rect 2380 51986 2436 51998
rect 2492 52834 2548 52846
rect 2492 52782 2494 52834
rect 2546 52782 2548 52834
rect 2380 51266 2436 51278
rect 2380 51214 2382 51266
rect 2434 51214 2436 51266
rect 2156 50482 2212 50494
rect 2156 50430 2158 50482
rect 2210 50430 2212 50482
rect 2156 50428 2212 50430
rect 1932 50370 1988 50382
rect 1932 50318 1934 50370
rect 1986 50318 1988 50370
rect 1932 50260 1988 50318
rect 1932 50194 1988 50204
rect 2044 50370 2100 50382
rect 2156 50372 2324 50428
rect 2044 50318 2046 50370
rect 2098 50318 2100 50370
rect 2044 50148 2100 50318
rect 2044 50082 2100 50092
rect 1820 49868 2100 49924
rect 1932 49700 1988 49710
rect 1932 49606 1988 49644
rect 2044 49140 2100 49868
rect 1820 49084 2100 49140
rect 2156 49810 2212 49822
rect 2156 49758 2158 49810
rect 2210 49758 2212 49810
rect 1708 49026 1764 49038
rect 1708 48974 1710 49026
rect 1762 48974 1764 49026
rect 1484 46834 1540 46844
rect 1596 48804 1652 48814
rect 1596 38724 1652 48748
rect 1708 48468 1764 48974
rect 1708 48402 1764 48412
rect 1820 43708 1876 49084
rect 2156 48356 2212 49758
rect 2044 48354 2212 48356
rect 2044 48302 2158 48354
rect 2210 48302 2212 48354
rect 2044 48300 2212 48302
rect 1932 45332 1988 45342
rect 2044 45332 2100 48300
rect 2156 48290 2212 48300
rect 2156 47684 2212 47694
rect 2268 47684 2324 50372
rect 2380 50260 2436 51214
rect 2492 50820 2548 52782
rect 2604 51268 2660 56140
rect 2716 52050 2772 52062
rect 2716 51998 2718 52050
rect 2770 51998 2772 52050
rect 2716 51492 2772 51998
rect 2716 51426 2772 51436
rect 2604 51212 2772 51268
rect 2492 50764 2660 50820
rect 2492 50596 2548 50606
rect 2492 50502 2548 50540
rect 2380 50194 2436 50204
rect 2492 50148 2548 50158
rect 2380 49812 2436 49822
rect 2492 49812 2548 50092
rect 2604 50034 2660 50764
rect 2604 49982 2606 50034
rect 2658 49982 2660 50034
rect 2604 49970 2660 49982
rect 2604 49812 2660 49822
rect 2492 49810 2660 49812
rect 2492 49758 2606 49810
rect 2658 49758 2660 49810
rect 2492 49756 2660 49758
rect 2380 49718 2436 49756
rect 2604 49746 2660 49756
rect 2716 49140 2772 51212
rect 2828 50484 2884 50522
rect 2828 50418 2884 50428
rect 2940 50036 2996 56252
rect 2156 47682 2324 47684
rect 2156 47630 2158 47682
rect 2210 47630 2324 47682
rect 2156 47628 2324 47630
rect 2156 47618 2212 47628
rect 2156 45332 2212 45342
rect 2044 45330 2212 45332
rect 2044 45278 2158 45330
rect 2210 45278 2212 45330
rect 2044 45276 2212 45278
rect 1932 45238 1988 45276
rect 2156 44322 2212 45276
rect 2268 45220 2324 47628
rect 2380 49084 2772 49140
rect 2828 49980 2996 50036
rect 2380 45332 2436 49084
rect 2492 48914 2548 48926
rect 2492 48862 2494 48914
rect 2546 48862 2548 48914
rect 2492 48466 2548 48862
rect 2492 48414 2494 48466
rect 2546 48414 2548 48466
rect 2492 48402 2548 48414
rect 2492 48244 2548 48254
rect 2492 48150 2548 48188
rect 2716 48242 2772 48254
rect 2716 48190 2718 48242
rect 2770 48190 2772 48242
rect 2604 48018 2660 48030
rect 2604 47966 2606 48018
rect 2658 47966 2660 48018
rect 2492 47684 2548 47694
rect 2604 47684 2660 47966
rect 2492 47682 2660 47684
rect 2492 47630 2494 47682
rect 2546 47630 2660 47682
rect 2492 47628 2660 47630
rect 2492 47618 2548 47628
rect 2492 47460 2548 47470
rect 2492 47366 2548 47404
rect 2716 47068 2772 48190
rect 2828 47460 2884 49980
rect 2940 49810 2996 49822
rect 2940 49758 2942 49810
rect 2994 49758 2996 49810
rect 2940 49700 2996 49758
rect 2940 49634 2996 49644
rect 2940 47460 2996 47470
rect 2884 47458 2996 47460
rect 2884 47406 2942 47458
rect 2994 47406 2996 47458
rect 2884 47404 2996 47406
rect 2828 47366 2884 47404
rect 2940 47394 2996 47404
rect 2716 47012 2996 47068
rect 2380 45266 2436 45276
rect 2828 45332 2884 45342
rect 2268 45154 2324 45164
rect 2492 45108 2548 45118
rect 2492 45014 2548 45052
rect 2828 45106 2884 45276
rect 2828 45054 2830 45106
rect 2882 45054 2884 45106
rect 2828 45042 2884 45054
rect 2828 44882 2884 44894
rect 2828 44830 2830 44882
rect 2882 44830 2884 44882
rect 2716 44548 2772 44558
rect 2828 44548 2884 44830
rect 2716 44546 2884 44548
rect 2716 44494 2718 44546
rect 2770 44494 2884 44546
rect 2716 44492 2884 44494
rect 2716 44482 2772 44492
rect 2156 44270 2158 44322
rect 2210 44270 2212 44322
rect 1820 43652 2100 43708
rect 1820 40402 1876 40414
rect 1820 40350 1822 40402
rect 1874 40350 1876 40402
rect 1820 39618 1876 40350
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 39284 1876 39566
rect 1820 39218 1876 39228
rect 1596 38658 1652 38668
rect 1708 38834 1764 38846
rect 1708 38782 1710 38834
rect 1762 38782 1764 38834
rect 1708 38612 1764 38782
rect 1764 38556 1876 38612
rect 1708 38546 1764 38556
rect 1820 38162 1876 38556
rect 1820 38110 1822 38162
rect 1874 38110 1876 38162
rect 1820 38098 1876 38110
rect 2044 37716 2100 43652
rect 2156 43650 2212 44270
rect 2940 44322 2996 47012
rect 2940 44270 2942 44322
rect 2994 44270 2996 44322
rect 2380 44210 2436 44222
rect 2380 44158 2382 44210
rect 2434 44158 2436 44210
rect 2380 43708 2436 44158
rect 2156 43598 2158 43650
rect 2210 43598 2212 43650
rect 2156 43586 2212 43598
rect 2268 43652 2436 43708
rect 2492 44098 2548 44110
rect 2492 44046 2494 44098
rect 2546 44046 2548 44098
rect 2268 43586 2324 43596
rect 2380 43540 2436 43550
rect 2380 43446 2436 43484
rect 2268 43426 2324 43438
rect 2268 43374 2270 43426
rect 2322 43374 2324 43426
rect 2156 41076 2212 41086
rect 2156 40982 2212 41020
rect 2268 40516 2324 43374
rect 2492 41188 2548 44046
rect 2604 44100 2660 44110
rect 2604 43538 2660 44044
rect 2604 43486 2606 43538
rect 2658 43486 2660 43538
rect 2604 43474 2660 43486
rect 2940 43538 2996 44270
rect 2940 43486 2942 43538
rect 2994 43486 2996 43538
rect 2940 43316 2996 43486
rect 2940 43250 2996 43260
rect 2716 41412 2772 41422
rect 2492 41132 2660 41188
rect 2492 40964 2548 40974
rect 2492 40870 2548 40908
rect 2492 40516 2548 40526
rect 2268 40514 2548 40516
rect 2268 40462 2494 40514
rect 2546 40462 2548 40514
rect 2268 40460 2548 40462
rect 2492 40450 2548 40460
rect 2492 39732 2548 39742
rect 2604 39732 2660 41132
rect 2492 39730 2660 39732
rect 2492 39678 2494 39730
rect 2546 39678 2660 39730
rect 2492 39676 2660 39678
rect 2492 39666 2548 39676
rect 2604 39284 2660 39294
rect 2604 39058 2660 39228
rect 2604 39006 2606 39058
rect 2658 39006 2660 39058
rect 2604 38994 2660 39006
rect 2156 38724 2212 38734
rect 2716 38668 2772 41356
rect 2828 40962 2884 40974
rect 2828 40910 2830 40962
rect 2882 40910 2884 40962
rect 2828 38836 2884 40910
rect 2940 38836 2996 38846
rect 2828 38834 2996 38836
rect 2828 38782 2942 38834
rect 2994 38782 2996 38834
rect 2828 38780 2996 38782
rect 2156 38630 2212 38668
rect 2604 38612 2772 38668
rect 2044 37660 2212 37716
rect 2044 37492 2100 37502
rect 1932 37436 2044 37492
rect 1372 36642 1428 36652
rect 1820 37154 1876 37166
rect 1820 37102 1822 37154
rect 1874 37102 1876 37154
rect 1596 36484 1652 36494
rect 1596 24052 1652 36428
rect 1708 36260 1764 36270
rect 1820 36260 1876 37102
rect 1708 36258 1876 36260
rect 1708 36206 1710 36258
rect 1762 36206 1876 36258
rect 1708 36204 1876 36206
rect 1708 36148 1764 36204
rect 1708 36082 1764 36092
rect 1820 35700 1876 35710
rect 1932 35700 1988 37436
rect 2044 37426 2100 37436
rect 1820 35698 1988 35700
rect 1820 35646 1822 35698
rect 1874 35646 1988 35698
rect 1820 35644 1988 35646
rect 1708 34130 1764 34142
rect 1708 34078 1710 34130
rect 1762 34078 1764 34130
rect 1708 33684 1764 34078
rect 1708 33618 1764 33628
rect 1820 33124 1876 35644
rect 2156 34132 2212 37660
rect 2268 36596 2324 36606
rect 2268 36502 2324 36540
rect 2268 35588 2324 35598
rect 2268 34914 2324 35532
rect 2268 34862 2270 34914
rect 2322 34862 2324 34914
rect 2268 34850 2324 34862
rect 2492 35586 2548 35598
rect 2492 35534 2494 35586
rect 2546 35534 2548 35586
rect 2492 34802 2548 35534
rect 2492 34750 2494 34802
rect 2546 34750 2548 34802
rect 2492 34738 2548 34750
rect 2604 34244 2660 38612
rect 2940 38164 2996 38780
rect 2940 38098 2996 38108
rect 3052 35364 3108 57036
rect 3164 51266 3220 51278
rect 3164 51214 3166 51266
rect 3218 51214 3220 51266
rect 3164 50596 3220 51214
rect 3164 46340 3220 50540
rect 3276 50260 3332 73164
rect 3388 71428 3444 73276
rect 3388 71362 3444 71372
rect 3388 60452 3444 60462
rect 3388 57428 3444 60396
rect 3948 58828 4004 73948
rect 4060 74060 4228 74116
rect 4060 73330 4116 74060
rect 4284 74004 4340 75068
rect 4844 74900 4900 74910
rect 4844 74806 4900 74844
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4172 73948 4340 74004
rect 4732 74004 4788 74014
rect 4172 73890 4228 73948
rect 4732 73910 4788 73948
rect 5180 73948 5236 75628
rect 5404 75012 5460 75022
rect 5404 74918 5460 74956
rect 6636 75012 6692 75022
rect 6636 74918 6692 74956
rect 5740 74900 5796 74910
rect 5852 74900 5908 74910
rect 5796 74898 5908 74900
rect 5796 74846 5854 74898
rect 5906 74846 5908 74898
rect 5796 74844 5908 74846
rect 5740 74004 5796 74844
rect 5852 74834 5908 74844
rect 5180 73892 5460 73948
rect 5740 73910 5796 73948
rect 4172 73838 4174 73890
rect 4226 73838 4228 73890
rect 4172 73826 4228 73838
rect 4060 73278 4062 73330
rect 4114 73278 4116 73330
rect 4060 73266 4116 73278
rect 4844 73220 4900 73230
rect 4844 73126 4900 73164
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 4956 71540 5012 71550
rect 4284 71428 4340 71438
rect 4284 71092 4340 71372
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 4284 70082 4340 71036
rect 4284 70030 4286 70082
rect 4338 70030 4340 70082
rect 4284 70018 4340 70030
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 4172 65604 4228 65614
rect 4060 61460 4116 61470
rect 4060 61010 4116 61404
rect 4060 60958 4062 61010
rect 4114 60958 4116 61010
rect 4060 60946 4116 60958
rect 3948 58772 4116 58828
rect 3500 57652 3556 57662
rect 3948 57652 4004 57662
rect 3500 57650 4004 57652
rect 3500 57598 3502 57650
rect 3554 57598 3950 57650
rect 4002 57598 4004 57650
rect 3500 57596 4004 57598
rect 3500 57586 3556 57596
rect 3948 57586 4004 57596
rect 3388 57372 3556 57428
rect 3276 50194 3332 50204
rect 3388 54404 3444 54414
rect 3388 49698 3444 54348
rect 3388 49646 3390 49698
rect 3442 49646 3444 49698
rect 3388 48242 3444 49646
rect 3500 48580 3556 57372
rect 4060 52948 4116 58772
rect 4172 53172 4228 65548
rect 4396 65492 4452 65502
rect 4284 65436 4396 65492
rect 4284 63364 4340 65436
rect 4396 65398 4452 65436
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4284 63308 4676 63364
rect 4620 62692 4676 63308
rect 4620 62578 4676 62636
rect 4620 62526 4622 62578
rect 4674 62526 4676 62578
rect 4620 62514 4676 62526
rect 4956 62580 5012 71484
rect 5068 66052 5124 66062
rect 5068 65602 5124 65996
rect 5404 65828 5460 73892
rect 5628 73220 5684 73230
rect 5628 72434 5684 73164
rect 6972 73218 7028 76414
rect 8764 76466 8820 76478
rect 10892 76468 10948 76478
rect 12460 76468 12516 76478
rect 8764 76414 8766 76466
rect 8818 76414 8820 76466
rect 8764 74786 8820 76414
rect 10444 76466 10948 76468
rect 10444 76414 10894 76466
rect 10946 76414 10948 76466
rect 10444 76412 10948 76414
rect 9100 75682 9156 75694
rect 9100 75630 9102 75682
rect 9154 75630 9156 75682
rect 9100 75012 9156 75630
rect 9100 74946 9156 74956
rect 8764 74734 8766 74786
rect 8818 74734 8820 74786
rect 8764 74722 8820 74734
rect 9100 74788 9156 74798
rect 9100 74116 9156 74732
rect 9660 74788 9716 74798
rect 9660 74694 9716 74732
rect 9100 74022 9156 74060
rect 9884 74004 9940 74014
rect 9884 74002 10052 74004
rect 9884 73950 9886 74002
rect 9938 73950 10052 74002
rect 9884 73948 10052 73950
rect 9884 73938 9940 73948
rect 9996 73892 10388 73948
rect 7532 73780 7588 73790
rect 6972 73166 6974 73218
rect 7026 73166 7028 73218
rect 6972 73154 7028 73166
rect 7420 73220 7476 73230
rect 7532 73220 7588 73724
rect 10332 73554 10388 73892
rect 10332 73502 10334 73554
rect 10386 73502 10388 73554
rect 10332 73490 10388 73502
rect 7420 73218 7588 73220
rect 7420 73166 7422 73218
rect 7474 73166 7588 73218
rect 7420 73164 7588 73166
rect 7420 73154 7476 73164
rect 5628 72382 5630 72434
rect 5682 72382 5684 72434
rect 5628 72370 5684 72382
rect 5852 72546 5908 72558
rect 5852 72494 5854 72546
rect 5906 72494 5908 72546
rect 5852 72436 5908 72494
rect 7532 72546 7588 73164
rect 8316 73444 8372 73454
rect 8316 72658 8372 73388
rect 9548 73444 9604 73454
rect 9548 73350 9604 73388
rect 9884 73330 9940 73342
rect 9884 73278 9886 73330
rect 9938 73278 9940 73330
rect 9100 73220 9156 73230
rect 9884 73220 9940 73278
rect 9100 73218 9940 73220
rect 9100 73166 9102 73218
rect 9154 73166 9940 73218
rect 9100 73164 9940 73166
rect 9100 73154 9156 73164
rect 8316 72606 8318 72658
rect 8370 72606 8372 72658
rect 8316 72594 8372 72606
rect 7532 72494 7534 72546
rect 7586 72494 7588 72546
rect 5852 72370 5908 72380
rect 6524 72436 6580 72446
rect 6524 72342 6580 72380
rect 6300 71092 6356 71102
rect 6300 70998 6356 71036
rect 6188 70756 6244 70766
rect 6076 70754 6244 70756
rect 6076 70702 6190 70754
rect 6242 70702 6244 70754
rect 6076 70700 6244 70702
rect 5852 69188 5908 69198
rect 5740 69186 5908 69188
rect 5740 69134 5854 69186
rect 5906 69134 5908 69186
rect 5740 69132 5908 69134
rect 5628 66052 5684 66062
rect 5628 65958 5684 65996
rect 5404 65762 5460 65772
rect 5068 65550 5070 65602
rect 5122 65550 5124 65602
rect 5068 65538 5124 65550
rect 4956 62524 5124 62580
rect 4956 62356 5012 62366
rect 4844 62354 5012 62356
rect 4844 62302 4958 62354
rect 5010 62302 5012 62354
rect 4844 62300 5012 62302
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 4396 60900 4452 60910
rect 4844 60900 4900 62300
rect 4956 62290 5012 62300
rect 5068 62188 5124 62524
rect 5740 62468 5796 69132
rect 5852 69122 5908 69132
rect 5852 68628 5908 68638
rect 5852 68534 5908 68572
rect 6076 68626 6132 70700
rect 6188 70690 6244 70700
rect 6972 70754 7028 70766
rect 6972 70702 6974 70754
rect 7026 70702 7028 70754
rect 6188 70532 6244 70542
rect 6188 69410 6244 70476
rect 6524 70420 6580 70430
rect 6412 70084 6468 70094
rect 6188 69358 6190 69410
rect 6242 69358 6244 69410
rect 6188 69346 6244 69358
rect 6300 70082 6468 70084
rect 6300 70030 6414 70082
rect 6466 70030 6468 70082
rect 6300 70028 6468 70030
rect 6076 68574 6078 68626
rect 6130 68574 6132 68626
rect 6076 68562 6132 68574
rect 5964 68514 6020 68526
rect 5964 68462 5966 68514
rect 6018 68462 6020 68514
rect 5964 68404 6020 68462
rect 6300 68404 6356 70028
rect 6412 70018 6468 70028
rect 6412 69412 6468 69422
rect 6524 69412 6580 70364
rect 6412 69410 6580 69412
rect 6412 69358 6414 69410
rect 6466 69358 6580 69410
rect 6412 69356 6580 69358
rect 6412 69346 6468 69356
rect 6636 69300 6692 69310
rect 6636 69206 6692 69244
rect 6972 69300 7028 70702
rect 7420 70756 7476 70766
rect 7532 70756 7588 72494
rect 8428 71204 8484 71214
rect 8428 70978 8484 71148
rect 9212 71204 9268 71214
rect 9212 71090 9268 71148
rect 9212 71038 9214 71090
rect 9266 71038 9268 71090
rect 9212 71026 9268 71038
rect 8428 70926 8430 70978
rect 8482 70926 8484 70978
rect 7420 70754 7588 70756
rect 7420 70702 7422 70754
rect 7474 70702 7588 70754
rect 7420 70700 7588 70702
rect 8204 70866 8260 70878
rect 8204 70814 8206 70866
rect 8258 70814 8260 70866
rect 8204 70756 8260 70814
rect 7084 70644 7140 70654
rect 7084 69636 7140 70588
rect 7196 70196 7252 70206
rect 7420 70196 7476 70700
rect 8204 70690 8260 70700
rect 7644 70420 7700 70430
rect 8428 70420 8484 70926
rect 7644 70326 7700 70364
rect 8316 70364 8428 70420
rect 8204 70308 8260 70318
rect 8204 70196 8260 70252
rect 7196 70194 7476 70196
rect 7196 70142 7198 70194
rect 7250 70142 7476 70194
rect 7196 70140 7476 70142
rect 7980 70194 8260 70196
rect 7980 70142 8206 70194
rect 8258 70142 8260 70194
rect 7980 70140 8260 70142
rect 7196 70130 7252 70140
rect 7084 69580 7252 69636
rect 6972 69234 7028 69244
rect 7084 69188 7140 69198
rect 7084 69094 7140 69132
rect 6412 68964 6468 68974
rect 6412 68738 6468 68908
rect 6412 68686 6414 68738
rect 6466 68686 6468 68738
rect 6412 68674 6468 68686
rect 5964 68348 6356 68404
rect 6636 68628 6692 68638
rect 6636 67954 6692 68572
rect 6636 67902 6638 67954
rect 6690 67902 6692 67954
rect 6524 67620 6580 67630
rect 6524 66386 6580 67564
rect 6636 67284 6692 67902
rect 7196 67842 7252 69580
rect 7980 69298 8036 70140
rect 8204 70130 8260 70140
rect 8316 69636 8372 70364
rect 8428 70354 8484 70364
rect 8652 70754 8708 70766
rect 8652 70702 8654 70754
rect 8706 70702 8708 70754
rect 8652 70308 8708 70702
rect 8764 70756 8820 70766
rect 8764 70754 9044 70756
rect 8764 70702 8766 70754
rect 8818 70702 9044 70754
rect 8764 70700 9044 70702
rect 8764 70690 8820 70700
rect 8764 70308 8820 70318
rect 8540 70306 8820 70308
rect 8540 70254 8766 70306
rect 8818 70254 8820 70306
rect 8540 70252 8820 70254
rect 7980 69246 7982 69298
rect 8034 69246 8036 69298
rect 7308 68516 7364 68526
rect 7308 68514 7924 68516
rect 7308 68462 7310 68514
rect 7362 68462 7924 68514
rect 7308 68460 7924 68462
rect 7308 68450 7364 68460
rect 7644 67956 7700 67966
rect 7644 67862 7700 67900
rect 7196 67790 7198 67842
rect 7250 67790 7252 67842
rect 7196 67778 7252 67790
rect 7532 67732 7588 67742
rect 7532 67638 7588 67676
rect 7756 67620 7812 67630
rect 7756 67526 7812 67564
rect 6636 67218 6692 67228
rect 7756 67284 7812 67294
rect 6524 66334 6526 66386
rect 6578 66334 6580 66386
rect 6524 66322 6580 66334
rect 6748 67170 6804 67182
rect 6748 67118 6750 67170
rect 6802 67118 6804 67170
rect 6748 66276 6804 67118
rect 6748 66210 6804 66220
rect 7084 67058 7140 67070
rect 7084 67006 7086 67058
rect 7138 67006 7140 67058
rect 5964 66162 6020 66174
rect 5964 66110 5966 66162
rect 6018 66110 6020 66162
rect 5964 64930 6020 66110
rect 5964 64878 5966 64930
rect 6018 64878 6020 64930
rect 5964 64866 6020 64878
rect 6188 65268 6244 65278
rect 6188 64818 6244 65212
rect 6188 64766 6190 64818
rect 6242 64766 6244 64818
rect 6188 64754 6244 64766
rect 6524 64706 6580 64718
rect 6524 64654 6526 64706
rect 6578 64654 6580 64706
rect 6524 64484 6580 64654
rect 6524 64418 6580 64428
rect 6748 64708 6804 64718
rect 6636 63252 6692 63262
rect 6636 63158 6692 63196
rect 6300 62916 6356 62954
rect 6300 62850 6356 62860
rect 5740 62402 5796 62412
rect 6412 62466 6468 62478
rect 6412 62414 6414 62466
rect 6466 62414 6468 62466
rect 5852 62356 5908 62366
rect 6300 62356 6356 62366
rect 5852 62354 6356 62356
rect 5852 62302 5854 62354
rect 5906 62302 6302 62354
rect 6354 62302 6356 62354
rect 5852 62300 6356 62302
rect 5852 62290 5908 62300
rect 6300 62290 6356 62300
rect 6412 62356 6468 62414
rect 6412 62290 6468 62300
rect 6636 62356 6692 62366
rect 6748 62356 6804 64652
rect 6636 62354 6804 62356
rect 6636 62302 6638 62354
rect 6690 62302 6804 62354
rect 6636 62300 6804 62302
rect 6636 62290 6692 62300
rect 4396 60898 4900 60900
rect 4396 60846 4398 60898
rect 4450 60846 4900 60898
rect 4396 60844 4900 60846
rect 4956 62132 5124 62188
rect 5740 62242 5796 62254
rect 5740 62190 5742 62242
rect 5794 62190 5796 62242
rect 5740 62188 5796 62190
rect 5740 62132 6020 62188
rect 4396 60834 4452 60844
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4956 58884 5012 62132
rect 5068 61684 5124 61694
rect 5068 61682 5236 61684
rect 5068 61630 5070 61682
rect 5122 61630 5236 61682
rect 5068 61628 5236 61630
rect 5068 61618 5124 61628
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4956 58818 5012 58828
rect 5180 61572 5236 61628
rect 4476 58762 4740 58772
rect 5180 58436 5236 61516
rect 5852 61572 5908 61582
rect 5516 61460 5572 61470
rect 5516 60788 5572 61404
rect 5740 61458 5796 61470
rect 5740 61406 5742 61458
rect 5794 61406 5796 61458
rect 5740 61348 5796 61406
rect 5852 61458 5908 61516
rect 5852 61406 5854 61458
rect 5906 61406 5908 61458
rect 5852 61394 5908 61406
rect 5740 61282 5796 61292
rect 5180 58370 5236 58380
rect 5292 60676 5348 60686
rect 5516 60676 5572 60732
rect 5292 60674 5572 60676
rect 5292 60622 5294 60674
rect 5346 60622 5572 60674
rect 5292 60620 5572 60622
rect 5852 61236 5908 61246
rect 5852 60676 5908 61180
rect 5964 60900 6020 62132
rect 6300 61572 6356 61582
rect 6300 61478 6356 61516
rect 6076 61348 6132 61358
rect 6076 61346 6580 61348
rect 6076 61294 6078 61346
rect 6130 61294 6580 61346
rect 6076 61292 6580 61294
rect 6076 61282 6132 61292
rect 5964 60844 6468 60900
rect 6412 60786 6468 60844
rect 6412 60734 6414 60786
rect 6466 60734 6468 60786
rect 5964 60676 6020 60686
rect 5852 60674 6020 60676
rect 5852 60622 5966 60674
rect 6018 60622 6020 60674
rect 5852 60620 6020 60622
rect 5292 58996 5348 60620
rect 5964 59780 6020 60620
rect 6300 60562 6356 60574
rect 6300 60510 6302 60562
rect 6354 60510 6356 60562
rect 5852 59724 6020 59780
rect 6188 59778 6244 59790
rect 6188 59726 6190 59778
rect 6242 59726 6244 59778
rect 5628 58996 5684 59006
rect 5292 58994 5684 58996
rect 5292 58942 5630 58994
rect 5682 58942 5684 58994
rect 5292 58940 5684 58942
rect 4620 58212 4676 58222
rect 4620 57650 4676 58156
rect 4620 57598 4622 57650
rect 4674 57598 4676 57650
rect 4620 57586 4676 57598
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4844 56978 4900 56990
rect 4844 56926 4846 56978
rect 4898 56926 4900 56978
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4844 54628 4900 56926
rect 4844 54562 4900 54572
rect 5068 55970 5124 55982
rect 5068 55918 5070 55970
rect 5122 55918 5124 55970
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4620 53844 4676 53854
rect 4172 53106 4228 53116
rect 4284 53842 4676 53844
rect 4284 53790 4622 53842
rect 4674 53790 4676 53842
rect 4284 53788 4676 53790
rect 3948 52892 4116 52948
rect 3612 52052 3668 52062
rect 3612 51958 3668 51996
rect 3836 51940 3892 51950
rect 3724 50708 3780 50718
rect 3724 50614 3780 50652
rect 3836 50484 3892 51884
rect 3836 50034 3892 50428
rect 3836 49982 3838 50034
rect 3890 49982 3892 50034
rect 3836 49970 3892 49982
rect 3500 48524 3780 48580
rect 3612 48356 3668 48366
rect 3612 48262 3668 48300
rect 3388 48190 3390 48242
rect 3442 48190 3444 48242
rect 3388 47572 3444 48190
rect 3388 47506 3444 47516
rect 3500 48244 3556 48254
rect 3500 46786 3556 48188
rect 3500 46734 3502 46786
rect 3554 46734 3556 46786
rect 3500 46722 3556 46734
rect 3612 47684 3668 47694
rect 3612 46564 3668 47628
rect 3500 46508 3668 46564
rect 3164 46284 3332 46340
rect 3164 45220 3220 45230
rect 3164 45126 3220 45164
rect 3276 44660 3332 46284
rect 3164 44604 3332 44660
rect 3388 45220 3444 45230
rect 3164 43708 3220 44604
rect 3276 44212 3332 44222
rect 3388 44212 3444 45164
rect 3276 44210 3388 44212
rect 3276 44158 3278 44210
rect 3330 44158 3388 44210
rect 3276 44156 3388 44158
rect 3276 44146 3332 44156
rect 3388 44118 3444 44156
rect 3500 43988 3556 46508
rect 3388 43932 3556 43988
rect 3612 44996 3668 45006
rect 3612 44098 3668 44940
rect 3612 44046 3614 44098
rect 3666 44046 3668 44098
rect 3612 43988 3668 44046
rect 3164 43652 3332 43708
rect 3164 42642 3220 42654
rect 3164 42590 3166 42642
rect 3218 42590 3220 42642
rect 3164 41972 3220 42590
rect 3164 41906 3220 41916
rect 3164 41074 3220 41086
rect 3164 41022 3166 41074
rect 3218 41022 3220 41074
rect 3164 40964 3220 41022
rect 3164 39732 3220 40908
rect 3164 39666 3220 39676
rect 2716 35308 3108 35364
rect 2716 34356 2772 35308
rect 2716 34354 2884 34356
rect 2716 34302 2718 34354
rect 2770 34302 2884 34354
rect 2716 34300 2884 34302
rect 2716 34290 2772 34300
rect 2380 34188 2660 34244
rect 2044 34076 2212 34132
rect 2268 34132 2324 34142
rect 2044 33684 2100 34076
rect 2268 34038 2324 34076
rect 2044 33618 2100 33628
rect 2156 33908 2212 33918
rect 2380 33908 2436 34188
rect 2716 34020 2772 34030
rect 2716 33926 2772 33964
rect 2156 33570 2212 33852
rect 2156 33518 2158 33570
rect 2210 33518 2212 33570
rect 2156 33460 2212 33518
rect 1932 33404 2212 33460
rect 1932 33346 1988 33404
rect 1932 33294 1934 33346
rect 1986 33294 1988 33346
rect 1932 33282 1988 33294
rect 1708 33068 1876 33124
rect 1932 33124 1988 33134
rect 1708 30996 1764 33068
rect 1820 32788 1876 32798
rect 1932 32788 1988 33068
rect 1820 32786 1988 32788
rect 1820 32734 1822 32786
rect 1874 32734 1988 32786
rect 1820 32732 1988 32734
rect 1820 32722 1876 32732
rect 2044 32340 2100 32350
rect 1932 31668 1988 31678
rect 1932 31574 1988 31612
rect 1932 31220 1988 31230
rect 1708 30994 1876 30996
rect 1708 30942 1710 30994
rect 1762 30942 1876 30994
rect 1708 30940 1876 30942
rect 1708 30930 1764 30940
rect 1708 29988 1764 29998
rect 1708 29426 1764 29932
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 29092 1764 29374
rect 1820 29316 1876 30940
rect 1932 30324 1988 31164
rect 1932 30210 1988 30268
rect 1932 30158 1934 30210
rect 1986 30158 1988 30210
rect 1932 30146 1988 30158
rect 1820 29250 1876 29260
rect 1708 29036 1876 29092
rect 1820 28756 1876 29036
rect 1820 28690 1876 28700
rect 1708 28644 1764 28654
rect 1708 28550 1764 28588
rect 1820 27746 1876 27758
rect 1820 27694 1822 27746
rect 1874 27694 1876 27746
rect 1820 27074 1876 27694
rect 2044 27188 2100 32284
rect 2156 31778 2212 33404
rect 2156 31726 2158 31778
rect 2210 31726 2212 31778
rect 2156 31714 2212 31726
rect 2268 33852 2436 33908
rect 2268 31556 2324 33852
rect 2380 33572 2436 33582
rect 2380 33234 2436 33516
rect 2380 33182 2382 33234
rect 2434 33182 2436 33234
rect 2380 33170 2436 33182
rect 2492 33458 2548 33470
rect 2492 33406 2494 33458
rect 2546 33406 2548 33458
rect 2492 33236 2548 33406
rect 2828 33460 2884 34300
rect 2940 33908 2996 33918
rect 2996 33852 3220 33908
rect 2940 33814 2996 33852
rect 2940 33460 2996 33470
rect 2828 33458 2996 33460
rect 2828 33406 2942 33458
rect 2994 33406 2996 33458
rect 2828 33404 2996 33406
rect 2940 33394 2996 33404
rect 2492 33180 2884 33236
rect 2828 33012 2884 33180
rect 2716 32956 2884 33012
rect 2492 32788 2548 32798
rect 2492 32562 2548 32732
rect 2492 32510 2494 32562
rect 2546 32510 2548 32562
rect 2492 32498 2548 32510
rect 2716 32562 2772 32956
rect 2716 32510 2718 32562
rect 2770 32510 2772 32562
rect 2716 32498 2772 32510
rect 2828 32788 2884 32798
rect 2716 32116 2772 32126
rect 2716 32002 2772 32060
rect 2716 31950 2718 32002
rect 2770 31950 2772 32002
rect 2716 31938 2772 31950
rect 2492 31778 2548 31790
rect 2492 31726 2494 31778
rect 2546 31726 2548 31778
rect 2492 31668 2548 31726
rect 2828 31778 2884 32732
rect 3164 32674 3220 33852
rect 3164 32622 3166 32674
rect 3218 32622 3220 32674
rect 3164 32610 3220 32622
rect 2940 32564 2996 32574
rect 2940 32470 2996 32508
rect 2828 31726 2830 31778
rect 2882 31726 2884 31778
rect 2828 31714 2884 31726
rect 3052 32450 3108 32462
rect 3052 32398 3054 32450
rect 3106 32398 3108 32450
rect 2492 31602 2548 31612
rect 2156 31500 2324 31556
rect 2604 31556 2660 31566
rect 2604 31554 2772 31556
rect 2604 31502 2606 31554
rect 2658 31502 2772 31554
rect 2604 31500 2772 31502
rect 2156 29428 2212 31500
rect 2604 31490 2660 31500
rect 2492 30884 2548 30894
rect 2492 30882 2660 30884
rect 2492 30830 2494 30882
rect 2546 30830 2660 30882
rect 2492 30828 2660 30830
rect 2492 30818 2548 30828
rect 2604 30098 2660 30828
rect 2604 30046 2606 30098
rect 2658 30046 2660 30098
rect 2604 30034 2660 30046
rect 2268 29988 2324 29998
rect 2268 29894 2324 29932
rect 2716 29876 2772 31500
rect 2940 30884 2996 30894
rect 2940 30210 2996 30828
rect 2940 30158 2942 30210
rect 2994 30158 2996 30210
rect 2940 30146 2996 30158
rect 2492 29820 2772 29876
rect 2268 29428 2324 29438
rect 2156 29426 2324 29428
rect 2156 29374 2270 29426
rect 2322 29374 2324 29426
rect 2156 29372 2324 29374
rect 2268 29362 2324 29372
rect 2492 28754 2548 29820
rect 2492 28702 2494 28754
rect 2546 28702 2548 28754
rect 2492 28690 2548 28702
rect 2604 28644 2660 28654
rect 2492 28084 2548 28094
rect 2604 28084 2660 28588
rect 3052 28196 3108 32398
rect 3276 31780 3332 43652
rect 3388 39508 3444 43932
rect 3612 43922 3668 43932
rect 3724 44324 3780 48524
rect 3836 47572 3892 47582
rect 3836 47478 3892 47516
rect 3836 46676 3892 46686
rect 3836 45332 3892 46620
rect 3836 45266 3892 45276
rect 3948 44436 4004 52892
rect 4172 52164 4228 52174
rect 4172 52070 4228 52108
rect 4060 51938 4116 51950
rect 4060 51886 4062 51938
rect 4114 51886 4116 51938
rect 4060 50484 4116 51886
rect 4172 51492 4228 51502
rect 4172 51398 4228 51436
rect 4060 49812 4116 50428
rect 4284 50482 4340 53788
rect 4620 53778 4676 53788
rect 5068 53508 5124 55918
rect 5068 53414 5124 53452
rect 5180 54516 5236 54526
rect 4956 52946 5012 52958
rect 4956 52894 4958 52946
rect 5010 52894 5012 52946
rect 4620 52836 4676 52846
rect 4620 52834 4900 52836
rect 4620 52782 4622 52834
rect 4674 52782 4900 52834
rect 4620 52780 4900 52782
rect 4620 52770 4676 52780
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4732 52388 4788 52398
rect 4732 51378 4788 52332
rect 4844 52276 4900 52780
rect 4956 52386 5012 52894
rect 5180 52388 5236 54460
rect 4956 52334 4958 52386
rect 5010 52334 5012 52386
rect 4956 52322 5012 52334
rect 5068 52332 5236 52388
rect 4844 52210 4900 52220
rect 4732 51326 4734 51378
rect 4786 51326 4788 51378
rect 4732 51314 4788 51326
rect 4844 52050 4900 52062
rect 4844 51998 4846 52050
rect 4898 51998 4900 52050
rect 4844 51380 4900 51998
rect 4956 52052 5012 52062
rect 4956 51958 5012 51996
rect 5068 51716 5124 52332
rect 4844 51314 4900 51324
rect 4956 51660 5124 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4284 50430 4286 50482
rect 4338 50430 4340 50482
rect 4284 50418 4340 50430
rect 4508 50596 4564 50606
rect 4060 49746 4116 49756
rect 4508 49698 4564 50540
rect 4508 49646 4510 49698
rect 4562 49646 4564 49698
rect 4508 49588 4564 49646
rect 4284 49532 4564 49588
rect 4956 50482 5012 51660
rect 4956 50430 4958 50482
rect 5010 50430 5012 50482
rect 4956 49698 5012 50430
rect 4956 49646 4958 49698
rect 5010 49646 5012 49698
rect 4284 49476 4340 49532
rect 4060 49420 4340 49476
rect 4476 49420 4740 49430
rect 4060 45780 4116 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4732 48804 4788 48814
rect 4732 48802 4900 48804
rect 4732 48750 4734 48802
rect 4786 48750 4900 48802
rect 4732 48748 4900 48750
rect 4732 48738 4788 48748
rect 4396 48468 4452 48478
rect 4396 48354 4452 48412
rect 4844 48468 4900 48748
rect 4844 48374 4900 48412
rect 4396 48302 4398 48354
rect 4450 48302 4452 48354
rect 4396 48290 4452 48302
rect 4284 48244 4340 48254
rect 4172 47460 4228 47470
rect 4284 47460 4340 48188
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4732 47684 4788 47694
rect 4956 47684 5012 49646
rect 4788 47628 5012 47684
rect 4732 47618 4788 47628
rect 4844 47460 4900 47470
rect 4284 47404 4452 47460
rect 4172 47346 4228 47404
rect 4172 47294 4174 47346
rect 4226 47294 4228 47346
rect 4172 46676 4228 47294
rect 4396 47348 4452 47404
rect 4844 47366 4900 47404
rect 4396 47254 4452 47292
rect 4956 47348 5012 47358
rect 4956 47254 5012 47292
rect 4172 46610 4228 46620
rect 4284 47234 4340 47246
rect 5180 47236 5236 47246
rect 4284 47182 4286 47234
rect 4338 47182 4340 47234
rect 4284 45892 4340 47182
rect 5068 47234 5236 47236
rect 5068 47182 5182 47234
rect 5234 47182 5236 47234
rect 5068 47180 5236 47182
rect 4844 47124 4900 47134
rect 4844 46674 4900 47068
rect 5068 47012 5124 47180
rect 5180 47170 5236 47180
rect 4844 46622 4846 46674
rect 4898 46622 4900 46674
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4396 45892 4452 45902
rect 4284 45890 4452 45892
rect 4284 45838 4398 45890
rect 4450 45838 4452 45890
rect 4284 45836 4452 45838
rect 4396 45826 4452 45836
rect 4732 45892 4788 45902
rect 4844 45892 4900 46622
rect 4732 45890 4900 45892
rect 4732 45838 4734 45890
rect 4786 45838 4900 45890
rect 4732 45836 4900 45838
rect 4956 46956 5124 47012
rect 4956 45890 5012 46956
rect 4956 45838 4958 45890
rect 5010 45838 5012 45890
rect 4732 45826 4788 45836
rect 4956 45826 5012 45838
rect 4060 45724 4340 45780
rect 3948 44370 4004 44380
rect 3724 43762 3780 44268
rect 4172 44324 4228 44334
rect 3948 44212 4004 44222
rect 3948 44118 4004 44156
rect 4172 44210 4228 44268
rect 4172 44158 4174 44210
rect 4226 44158 4228 44210
rect 4172 44146 4228 44158
rect 4060 44100 4116 44110
rect 4060 44006 4116 44044
rect 4284 43988 4340 45724
rect 4844 45666 4900 45678
rect 4844 45614 4846 45666
rect 4898 45614 4900 45666
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4732 44100 4788 44110
rect 4732 44006 4788 44044
rect 3724 43710 3726 43762
rect 3778 43710 3780 43762
rect 3724 43698 3780 43710
rect 4172 43932 4340 43988
rect 3612 43652 3668 43662
rect 3388 39442 3444 39452
rect 3500 41076 3556 41086
rect 3388 38948 3444 38958
rect 3388 38834 3444 38892
rect 3388 38782 3390 38834
rect 3442 38782 3444 38834
rect 3388 38770 3444 38782
rect 3388 34020 3444 34030
rect 3388 33926 3444 33964
rect 3388 33572 3444 33582
rect 3388 33458 3444 33516
rect 3388 33406 3390 33458
rect 3442 33406 3444 33458
rect 3388 33394 3444 33406
rect 2492 28082 2660 28084
rect 2492 28030 2494 28082
rect 2546 28030 2660 28082
rect 2492 28028 2660 28030
rect 2828 28140 3108 28196
rect 3164 31724 3332 31780
rect 3388 32788 3444 32798
rect 2268 27860 2324 27870
rect 2268 27766 2324 27804
rect 2156 27188 2212 27198
rect 2044 27186 2212 27188
rect 2044 27134 2158 27186
rect 2210 27134 2212 27186
rect 2044 27132 2212 27134
rect 2156 27122 2212 27132
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 26908 1876 27022
rect 2492 26908 2548 28028
rect 1708 26852 1876 26908
rect 2044 26852 2548 26908
rect 2604 27076 2660 27086
rect 2604 26962 2660 27020
rect 2604 26910 2606 26962
rect 2658 26910 2660 26962
rect 2604 26898 2660 26910
rect 1708 26292 1764 26852
rect 1708 26226 1764 26236
rect 2044 26290 2100 26852
rect 2716 26404 2772 26414
rect 2828 26404 2884 28140
rect 3164 28084 3220 31724
rect 3276 31554 3332 31566
rect 3276 31502 3278 31554
rect 3330 31502 3332 31554
rect 3276 30324 3332 31502
rect 3276 30258 3332 30268
rect 3388 29988 3444 32732
rect 3500 30212 3556 41020
rect 3612 38668 3668 43596
rect 3724 42756 3780 42766
rect 3724 42662 3780 42700
rect 3724 41076 3780 41086
rect 3724 40982 3780 41020
rect 3948 39060 4004 39070
rect 3836 39004 3948 39060
rect 3612 38612 3780 38668
rect 3612 38500 3668 38510
rect 3612 34356 3668 38444
rect 3724 37826 3780 38612
rect 3836 38050 3892 39004
rect 3948 38966 4004 39004
rect 3836 37998 3838 38050
rect 3890 37998 3892 38050
rect 3836 37986 3892 37998
rect 3724 37774 3726 37826
rect 3778 37774 3780 37826
rect 3724 35028 3780 37774
rect 3948 37828 4004 37838
rect 3724 34962 3780 34972
rect 3836 36372 3892 36382
rect 3836 34802 3892 36316
rect 3836 34750 3838 34802
rect 3890 34750 3892 34802
rect 3836 34738 3892 34750
rect 3612 34290 3668 34300
rect 3836 34020 3892 34030
rect 3836 33458 3892 33964
rect 3836 33406 3838 33458
rect 3890 33406 3892 33458
rect 3836 33394 3892 33406
rect 3836 32564 3892 32574
rect 3836 32450 3892 32508
rect 3836 32398 3838 32450
rect 3890 32398 3892 32450
rect 3836 32004 3892 32398
rect 3836 31938 3892 31948
rect 3836 31778 3892 31790
rect 3836 31726 3838 31778
rect 3890 31726 3892 31778
rect 3836 31668 3892 31726
rect 3836 31602 3892 31612
rect 3500 30156 3668 30212
rect 3500 29988 3556 29998
rect 3388 29986 3556 29988
rect 3388 29934 3502 29986
rect 3554 29934 3556 29986
rect 3388 29932 3556 29934
rect 3500 29922 3556 29932
rect 3388 28084 3444 28094
rect 3164 28082 3444 28084
rect 3164 28030 3390 28082
rect 3442 28030 3444 28082
rect 3164 28028 3444 28030
rect 2940 27860 2996 27870
rect 2940 27766 2996 27804
rect 3276 27076 3332 28028
rect 3388 28018 3444 28028
rect 2716 26402 2884 26404
rect 2716 26350 2718 26402
rect 2770 26350 2884 26402
rect 2716 26348 2884 26350
rect 2940 26964 2996 27002
rect 3276 26982 3332 27020
rect 3612 27860 3668 30156
rect 2716 26338 2772 26348
rect 2044 26238 2046 26290
rect 2098 26238 2100 26290
rect 2044 26226 2100 26238
rect 1596 23986 1652 23996
rect 2268 24052 2324 24062
rect 2268 23958 2324 23996
rect 1708 23828 1764 23838
rect 1764 23772 1876 23828
rect 1708 23734 1764 23772
rect 1820 23378 1876 23772
rect 1820 23326 1822 23378
rect 1874 23326 1876 23378
rect 1820 23314 1876 23326
rect 1260 21634 1316 21644
rect 2268 21812 2324 21822
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21364 1764 21534
rect 2268 21586 2324 21756
rect 2268 21534 2270 21586
rect 2322 21534 2324 21586
rect 2268 21522 2324 21534
rect 1708 20916 1764 21308
rect 1820 20916 1876 20926
rect 1708 20914 1876 20916
rect 1708 20862 1822 20914
rect 1874 20862 1876 20914
rect 1708 20860 1876 20862
rect 1820 20850 1876 20860
rect 1148 20178 1204 20188
rect 2940 20188 2996 26908
rect 3612 26962 3668 27804
rect 3612 26910 3614 26962
rect 3666 26910 3668 26962
rect 3612 23604 3668 26910
rect 3612 23538 3668 23548
rect 2940 20132 3332 20188
rect 2716 3444 2772 3454
rect 2940 3444 2996 3454
rect 2716 3442 2996 3444
rect 2716 3390 2718 3442
rect 2770 3390 2942 3442
rect 2994 3390 2996 3442
rect 2716 3388 2996 3390
rect 2716 800 2772 3388
rect 2940 3378 2996 3388
rect 3276 3442 3332 20132
rect 3948 20020 4004 37772
rect 4060 35028 4116 35038
rect 4060 34934 4116 34972
rect 4172 34356 4228 43932
rect 4844 43876 4900 45614
rect 5180 45220 5236 45230
rect 4508 43820 4900 43876
rect 4956 44100 5012 44110
rect 4508 43540 4564 43820
rect 4956 43708 5012 44044
rect 4732 43652 4788 43662
rect 4956 43652 5124 43708
rect 4284 43538 4564 43540
rect 4284 43486 4510 43538
rect 4562 43486 4564 43538
rect 4284 43484 4564 43486
rect 4284 42756 4340 43484
rect 4508 43474 4564 43484
rect 4620 43540 4676 43550
rect 4620 43446 4676 43484
rect 4732 43428 4788 43596
rect 4956 43538 5012 43550
rect 4956 43486 4958 43538
rect 5010 43486 5012 43538
rect 4732 43362 4788 43372
rect 4844 43426 4900 43438
rect 4844 43374 4846 43426
rect 4898 43374 4900 43426
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4844 42868 4900 43374
rect 4620 42812 4900 42868
rect 4396 42756 4452 42766
rect 4284 42754 4452 42756
rect 4284 42702 4398 42754
rect 4450 42702 4452 42754
rect 4284 42700 4452 42702
rect 4396 42690 4452 42700
rect 4620 42084 4676 42812
rect 4956 42756 5012 43486
rect 5068 43204 5124 43652
rect 5068 43138 5124 43148
rect 4956 42690 5012 42700
rect 4956 42530 5012 42542
rect 4956 42478 4958 42530
rect 5010 42478 5012 42530
rect 4732 42084 4788 42094
rect 4620 42082 4788 42084
rect 4620 42030 4734 42082
rect 4786 42030 4788 42082
rect 4620 42028 4788 42030
rect 4732 42018 4788 42028
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4956 41076 5012 42478
rect 5180 42532 5236 45164
rect 5292 45108 5348 58940
rect 5628 58930 5684 58940
rect 5740 58212 5796 58222
rect 5740 58118 5796 58156
rect 5852 57988 5908 59724
rect 5964 59106 6020 59118
rect 5964 59054 5966 59106
rect 6018 59054 6020 59106
rect 5964 58994 6020 59054
rect 6188 59108 6244 59726
rect 6188 59042 6244 59052
rect 5964 58942 5966 58994
rect 6018 58942 6020 58994
rect 5964 58930 6020 58942
rect 6300 58884 6356 60510
rect 6412 60002 6468 60734
rect 6524 60340 6580 61292
rect 6636 60898 6692 60910
rect 6636 60846 6638 60898
rect 6690 60846 6692 60898
rect 6636 60788 6692 60846
rect 6748 60788 6804 62300
rect 6972 63252 7028 63262
rect 6972 62354 7028 63196
rect 6972 62302 6974 62354
rect 7026 62302 7028 62354
rect 6860 61348 6916 61358
rect 6860 61254 6916 61292
rect 6972 61236 7028 62302
rect 6972 61170 7028 61180
rect 6972 60788 7028 60798
rect 6748 60786 7028 60788
rect 6748 60734 6974 60786
rect 7026 60734 7028 60786
rect 6748 60732 7028 60734
rect 6636 60722 6692 60732
rect 6524 60284 6804 60340
rect 6748 60114 6804 60284
rect 6748 60062 6750 60114
rect 6802 60062 6804 60114
rect 6748 60050 6804 60062
rect 6412 59950 6414 60002
rect 6466 59950 6468 60002
rect 6412 59938 6468 59950
rect 6860 60002 6916 60014
rect 6860 59950 6862 60002
rect 6914 59950 6916 60002
rect 6076 58828 6356 58884
rect 6412 59108 6468 59118
rect 5964 58548 6020 58558
rect 5964 58322 6020 58492
rect 5964 58270 5966 58322
rect 6018 58270 6020 58322
rect 5964 58258 6020 58270
rect 6076 58324 6132 58828
rect 6300 58548 6356 58558
rect 6300 58454 6356 58492
rect 6076 58322 6356 58324
rect 6076 58270 6078 58322
rect 6130 58270 6356 58322
rect 6076 58268 6356 58270
rect 6076 58258 6132 58268
rect 5740 57932 5908 57988
rect 5740 56980 5796 57932
rect 5852 57764 5908 57774
rect 5964 57764 6020 57774
rect 5852 57762 5964 57764
rect 5852 57710 5854 57762
rect 5906 57710 5964 57762
rect 5852 57708 5964 57710
rect 5852 57698 5908 57708
rect 5740 56914 5796 56924
rect 5964 56754 6020 57708
rect 6300 57652 6356 58268
rect 6412 58322 6468 59052
rect 6412 58270 6414 58322
rect 6466 58270 6468 58322
rect 6412 58258 6468 58270
rect 6524 59106 6580 59118
rect 6524 59054 6526 59106
rect 6578 59054 6580 59106
rect 6524 58996 6580 59054
rect 6860 59108 6916 59950
rect 6860 59014 6916 59052
rect 6524 57764 6580 58940
rect 6748 58994 6804 59006
rect 6748 58942 6750 58994
rect 6802 58942 6804 58994
rect 6748 58884 6804 58942
rect 6748 58828 6916 58884
rect 6748 58548 6804 58558
rect 6636 58436 6692 58446
rect 6636 58342 6692 58380
rect 6524 57698 6580 57708
rect 6412 57652 6468 57662
rect 6300 57650 6468 57652
rect 6300 57598 6414 57650
rect 6466 57598 6468 57650
rect 6300 57596 6468 57598
rect 6412 57586 6468 57596
rect 6748 57650 6804 58492
rect 6860 58434 6916 58828
rect 6860 58382 6862 58434
rect 6914 58382 6916 58434
rect 6860 58370 6916 58382
rect 6748 57598 6750 57650
rect 6802 57598 6804 57650
rect 6748 57586 6804 57598
rect 6076 57538 6132 57550
rect 6076 57486 6078 57538
rect 6130 57486 6132 57538
rect 6076 57428 6132 57486
rect 6076 56868 6132 57372
rect 6636 57538 6692 57550
rect 6636 57486 6638 57538
rect 6690 57486 6692 57538
rect 6188 56868 6244 56878
rect 6076 56866 6356 56868
rect 6076 56814 6190 56866
rect 6242 56814 6356 56866
rect 6076 56812 6356 56814
rect 6188 56802 6244 56812
rect 5964 56702 5966 56754
rect 6018 56702 6020 56754
rect 5964 56420 6020 56702
rect 5964 56364 6244 56420
rect 5740 56196 5796 56206
rect 5516 53508 5572 53518
rect 5404 52722 5460 52734
rect 5404 52670 5406 52722
rect 5458 52670 5460 52722
rect 5404 47124 5460 52670
rect 5516 50428 5572 53452
rect 5628 52164 5684 52174
rect 5628 52070 5684 52108
rect 5628 51380 5684 51390
rect 5628 51286 5684 51324
rect 5628 50708 5684 50718
rect 5628 50594 5684 50652
rect 5628 50542 5630 50594
rect 5682 50542 5684 50594
rect 5628 50530 5684 50542
rect 5740 50428 5796 56140
rect 6188 55970 6244 56364
rect 6188 55918 6190 55970
rect 6242 55918 6244 55970
rect 6188 55860 6244 55918
rect 5964 55804 6244 55860
rect 5852 54516 5908 54526
rect 5852 54422 5908 54460
rect 5964 54292 6020 55804
rect 5852 54236 6020 54292
rect 6076 55410 6132 55422
rect 6076 55358 6078 55410
rect 6130 55358 6132 55410
rect 6076 54740 6132 55358
rect 6076 54514 6132 54684
rect 6188 54628 6244 54638
rect 6188 54534 6244 54572
rect 6076 54462 6078 54514
rect 6130 54462 6132 54514
rect 5852 52500 5908 54236
rect 6076 53956 6132 54462
rect 6076 53890 6132 53900
rect 5852 52434 5908 52444
rect 5964 53620 6020 53630
rect 5964 52946 6020 53564
rect 5964 52894 5966 52946
rect 6018 52894 6020 52946
rect 5964 52388 6020 52894
rect 5964 52322 6020 52332
rect 6076 53620 6132 53630
rect 6300 53620 6356 56812
rect 6636 56866 6692 57486
rect 6636 56814 6638 56866
rect 6690 56814 6692 56866
rect 6636 56802 6692 56814
rect 6972 56868 7028 60732
rect 7084 60452 7140 67006
rect 7308 65828 7364 65838
rect 7196 65604 7252 65614
rect 7196 65378 7252 65548
rect 7196 65326 7198 65378
rect 7250 65326 7252 65378
rect 7196 64708 7252 65326
rect 7196 64642 7252 64652
rect 7196 64484 7252 64494
rect 7196 63140 7252 64428
rect 7196 63074 7252 63084
rect 7084 60386 7140 60396
rect 7196 62916 7252 62926
rect 7196 62244 7252 62860
rect 7308 62468 7364 65772
rect 7644 65604 7700 65614
rect 7644 65510 7700 65548
rect 7756 65602 7812 67228
rect 7756 65550 7758 65602
rect 7810 65550 7812 65602
rect 7756 65380 7812 65550
rect 7644 65268 7700 65278
rect 7644 65174 7700 65212
rect 7756 63252 7812 65324
rect 7756 63186 7812 63196
rect 7644 63140 7700 63150
rect 7308 62412 7476 62468
rect 7308 62244 7364 62254
rect 7196 62242 7364 62244
rect 7196 62190 7310 62242
rect 7362 62190 7364 62242
rect 7196 62188 7364 62190
rect 7196 61348 7252 62188
rect 7308 62178 7364 62188
rect 7308 61796 7364 61806
rect 7308 61682 7364 61740
rect 7308 61630 7310 61682
rect 7362 61630 7364 61682
rect 7308 61618 7364 61630
rect 7196 58828 7252 61292
rect 7308 59444 7364 59454
rect 7420 59444 7476 62412
rect 7308 59442 7420 59444
rect 7308 59390 7310 59442
rect 7362 59390 7420 59442
rect 7308 59388 7420 59390
rect 7308 59378 7364 59388
rect 7420 59350 7476 59388
rect 7196 58772 7364 58828
rect 7196 57876 7252 57886
rect 7084 57650 7140 57662
rect 7084 57598 7086 57650
rect 7138 57598 7140 57650
rect 7084 57540 7140 57598
rect 7084 57474 7140 57484
rect 7084 56868 7140 56878
rect 6972 56812 7084 56868
rect 7084 56802 7140 56812
rect 6636 56642 6692 56654
rect 6636 56590 6638 56642
rect 6690 56590 6692 56642
rect 6524 55970 6580 55982
rect 6524 55918 6526 55970
rect 6578 55918 6580 55970
rect 6524 54516 6580 55918
rect 6524 54450 6580 54460
rect 6076 53618 6356 53620
rect 6076 53566 6078 53618
rect 6130 53566 6356 53618
rect 6076 53564 6356 53566
rect 6636 53620 6692 56590
rect 7084 56308 7140 56318
rect 7196 56308 7252 57820
rect 7084 56306 7252 56308
rect 7084 56254 7086 56306
rect 7138 56254 7252 56306
rect 7084 56252 7252 56254
rect 7084 56242 7140 56252
rect 7308 56084 7364 58772
rect 7420 58436 7476 58446
rect 7420 58342 7476 58380
rect 7532 58210 7588 58222
rect 7532 58158 7534 58210
rect 7586 58158 7588 58210
rect 7420 58100 7476 58110
rect 7420 56866 7476 58044
rect 7420 56814 7422 56866
rect 7474 56814 7476 56866
rect 7420 56802 7476 56814
rect 6076 51044 6132 53564
rect 6636 53554 6692 53564
rect 6748 56028 7364 56084
rect 6748 53284 6804 56028
rect 7084 54292 7140 54302
rect 6972 54290 7140 54292
rect 6972 54238 7086 54290
rect 7138 54238 7140 54290
rect 6972 54236 7140 54238
rect 6860 53618 6916 53630
rect 6860 53566 6862 53618
rect 6914 53566 6916 53618
rect 6860 53396 6916 53566
rect 6972 53396 7028 54236
rect 7084 54226 7140 54236
rect 7532 53396 7588 58158
rect 7644 57876 7700 63084
rect 7756 62356 7812 62394
rect 7756 62290 7812 62300
rect 7868 62188 7924 68460
rect 7980 68514 8036 69246
rect 8204 69580 8372 69636
rect 8428 69972 8484 69982
rect 7980 68462 7982 68514
rect 8034 68462 8036 68514
rect 7980 68450 8036 68462
rect 8092 68726 8148 68738
rect 8092 68674 8094 68726
rect 8146 68674 8148 68726
rect 8092 68628 8148 68674
rect 7980 67620 8036 67630
rect 8092 67620 8148 68572
rect 8204 67954 8260 69580
rect 8428 69412 8484 69916
rect 8316 69410 8484 69412
rect 8316 69358 8430 69410
rect 8482 69358 8484 69410
rect 8316 69356 8484 69358
rect 8316 68626 8372 69356
rect 8428 69346 8484 69356
rect 8540 69188 8596 70252
rect 8764 70242 8820 70252
rect 8988 70306 9044 70700
rect 9884 70644 9940 73164
rect 10444 72658 10500 76412
rect 10892 76402 10948 76412
rect 12012 76466 12516 76468
rect 12012 76414 12462 76466
rect 12514 76414 12516 76466
rect 12012 76412 12516 76414
rect 10668 74898 10724 74910
rect 10668 74846 10670 74898
rect 10722 74846 10724 74898
rect 10668 74788 10724 74846
rect 10668 74004 10724 74732
rect 11340 74788 11396 74798
rect 11340 74786 11844 74788
rect 11340 74734 11342 74786
rect 11394 74734 11844 74786
rect 11340 74732 11844 74734
rect 11340 74722 11396 74732
rect 10892 74004 10948 74014
rect 10668 73948 10892 74004
rect 10668 73330 10724 73342
rect 10668 73278 10670 73330
rect 10722 73278 10724 73330
rect 10668 72770 10724 73278
rect 10668 72718 10670 72770
rect 10722 72718 10724 72770
rect 10668 72706 10724 72718
rect 10444 72606 10446 72658
rect 10498 72606 10500 72658
rect 10444 72594 10500 72606
rect 10892 72658 10948 73948
rect 11788 73444 11844 74732
rect 12012 74226 12068 76412
rect 12460 76402 12516 76412
rect 13468 76466 13524 76478
rect 13468 76414 13470 76466
rect 13522 76414 13524 76466
rect 13468 74786 13524 76414
rect 13468 74734 13470 74786
rect 13522 74734 13524 74786
rect 13468 74722 13524 74734
rect 13580 76468 13636 76478
rect 12012 74174 12014 74226
rect 12066 74174 12068 74226
rect 12012 74162 12068 74174
rect 13468 74228 13524 74238
rect 13580 74228 13636 76412
rect 13916 76354 13972 76636
rect 15148 76468 15204 76478
rect 15148 76374 15204 76412
rect 13916 76302 13918 76354
rect 13970 76302 13972 76354
rect 13916 76290 13972 76302
rect 15596 76354 15652 77196
rect 16828 77026 16884 79200
rect 16828 76974 16830 77026
rect 16882 76974 16884 77026
rect 16828 76962 16884 76974
rect 17948 77026 18004 77038
rect 17948 76974 17950 77026
rect 18002 76974 18004 77026
rect 17948 76578 18004 76974
rect 18620 77026 18676 79200
rect 18620 76974 18622 77026
rect 18674 76974 18676 77026
rect 18620 76962 18676 76974
rect 19180 77026 19236 77038
rect 19180 76974 19182 77026
rect 19234 76974 19236 77026
rect 17948 76526 17950 76578
rect 18002 76526 18004 76578
rect 17948 76514 18004 76526
rect 19180 76578 19236 76974
rect 20412 77026 20468 79200
rect 20412 76974 20414 77026
rect 20466 76974 20468 77026
rect 20412 76962 20468 76974
rect 21532 77026 21588 77038
rect 21532 76974 21534 77026
rect 21586 76974 21588 77026
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 21532 76690 21588 76974
rect 22204 77026 22260 79200
rect 23996 77476 24052 79200
rect 23996 77420 24500 77476
rect 22204 76974 22206 77026
rect 22258 76974 22260 77026
rect 22204 76962 22260 76974
rect 23100 77026 23156 77038
rect 23100 76974 23102 77026
rect 23154 76974 23156 77026
rect 21532 76638 21534 76690
rect 21586 76638 21588 76690
rect 21532 76626 21588 76638
rect 19180 76526 19182 76578
rect 19234 76526 19236 76578
rect 19180 76514 19236 76526
rect 17052 76468 17108 76478
rect 15596 76302 15598 76354
rect 15650 76302 15652 76354
rect 15596 76290 15652 76302
rect 16828 76466 17108 76468
rect 16828 76414 17054 76466
rect 17106 76414 17108 76466
rect 16828 76412 17108 76414
rect 14700 75684 14756 75694
rect 13692 75458 13748 75470
rect 13692 75406 13694 75458
rect 13746 75406 13748 75458
rect 13692 74900 13748 75406
rect 14700 75010 14756 75628
rect 15932 75684 15988 75694
rect 15932 75570 15988 75628
rect 15932 75518 15934 75570
rect 15986 75518 15988 75570
rect 15932 75506 15988 75518
rect 16268 75570 16324 75582
rect 16268 75518 16270 75570
rect 16322 75518 16324 75570
rect 14700 74958 14702 75010
rect 14754 74958 14756 75010
rect 14700 74946 14756 74958
rect 14028 74900 14084 74910
rect 13692 74898 14084 74900
rect 13692 74846 14030 74898
rect 14082 74846 14084 74898
rect 13692 74844 14084 74846
rect 13468 74226 13636 74228
rect 13468 74174 13470 74226
rect 13522 74174 13636 74226
rect 13468 74172 13636 74174
rect 13468 74162 13524 74172
rect 12460 74004 12516 74014
rect 12460 73910 12516 73948
rect 14028 74004 14084 74844
rect 15596 74340 15652 74350
rect 15596 74226 15652 74284
rect 15596 74174 15598 74226
rect 15650 74174 15652 74226
rect 15596 74162 15652 74174
rect 14028 73938 14084 73948
rect 11788 73378 11844 73388
rect 13804 73332 13860 73342
rect 13804 73330 14196 73332
rect 13804 73278 13806 73330
rect 13858 73278 14196 73330
rect 13804 73276 14196 73278
rect 13804 73266 13860 73276
rect 11116 73218 11172 73230
rect 11116 73166 11118 73218
rect 11170 73166 11172 73218
rect 11004 72772 11060 72782
rect 11116 72772 11172 73166
rect 11004 72770 11172 72772
rect 11004 72718 11006 72770
rect 11058 72718 11172 72770
rect 11004 72716 11172 72718
rect 11004 72706 11060 72716
rect 10892 72606 10894 72658
rect 10946 72606 10948 72658
rect 10892 72594 10948 72606
rect 11116 71316 11172 72716
rect 11116 71250 11172 71260
rect 12796 72436 12852 72446
rect 12796 71090 12852 72380
rect 12796 71038 12798 71090
rect 12850 71038 12852 71090
rect 9884 70578 9940 70588
rect 9996 70978 10052 70990
rect 9996 70926 9998 70978
rect 10050 70926 10052 70978
rect 8988 70254 8990 70306
rect 9042 70254 9044 70306
rect 8988 70242 9044 70254
rect 9996 70420 10052 70926
rect 10668 70868 10724 70878
rect 11788 70868 11844 70878
rect 10668 70866 11396 70868
rect 10668 70814 10670 70866
rect 10722 70814 11396 70866
rect 10668 70812 11396 70814
rect 10668 70802 10724 70812
rect 8316 68574 8318 68626
rect 8370 68574 8372 68626
rect 8316 68562 8372 68574
rect 8428 69132 8596 69188
rect 8652 70082 8708 70094
rect 8652 70030 8654 70082
rect 8706 70030 8708 70082
rect 8204 67902 8206 67954
rect 8258 67902 8260 67954
rect 8204 67732 8260 67902
rect 8204 67666 8260 67676
rect 8036 67564 8148 67620
rect 7980 67554 8036 67564
rect 8316 65492 8372 65502
rect 8316 65398 8372 65436
rect 8428 65266 8484 69132
rect 8540 68964 8596 68974
rect 8652 68964 8708 70030
rect 9772 70082 9828 70094
rect 9772 70030 9774 70082
rect 9826 70030 9828 70082
rect 8596 68908 8708 68964
rect 8764 69410 8820 69422
rect 8764 69358 8766 69410
rect 8818 69358 8820 69410
rect 8764 69300 8820 69358
rect 8764 68964 8820 69244
rect 9772 68964 9828 70030
rect 9996 69410 10052 70364
rect 10444 70420 10500 70430
rect 10444 70326 10500 70364
rect 9996 69358 9998 69410
rect 10050 69358 10052 69410
rect 9996 69346 10052 69358
rect 10220 70196 10276 70206
rect 9996 68964 10052 68974
rect 9772 68908 9996 68964
rect 8540 68898 8596 68908
rect 8764 67396 8820 68908
rect 9548 68628 9604 68638
rect 9548 68534 9604 68572
rect 9996 68514 10052 68908
rect 9996 68462 9998 68514
rect 10050 68462 10052 68514
rect 9996 68450 10052 68462
rect 10220 68068 10276 70140
rect 8428 65214 8430 65266
rect 8482 65214 8484 65266
rect 8428 64930 8484 65214
rect 8428 64878 8430 64930
rect 8482 64878 8484 64930
rect 8428 64866 8484 64878
rect 8540 67340 8820 67396
rect 9884 68012 10276 68068
rect 7980 64596 8036 64606
rect 8316 64596 8372 64606
rect 7980 64594 8372 64596
rect 7980 64542 7982 64594
rect 8034 64542 8318 64594
rect 8370 64542 8372 64594
rect 7980 64540 8372 64542
rect 7980 64530 8036 64540
rect 8316 64372 8372 64540
rect 8540 64372 8596 67340
rect 9884 67058 9940 68012
rect 9884 67006 9886 67058
rect 9938 67006 9940 67058
rect 9884 66994 9940 67006
rect 10108 67842 10164 67854
rect 10108 67790 10110 67842
rect 10162 67790 10164 67842
rect 9436 66276 9492 66286
rect 9436 66182 9492 66220
rect 10108 66276 10164 67790
rect 10220 67732 10276 68012
rect 10668 69298 10724 69310
rect 10668 69246 10670 69298
rect 10722 69246 10724 69298
rect 10332 67732 10388 67742
rect 10220 67730 10388 67732
rect 10220 67678 10334 67730
rect 10386 67678 10388 67730
rect 10220 67676 10388 67678
rect 10332 67666 10388 67676
rect 10668 67396 10724 69246
rect 10668 67330 10724 67340
rect 10556 66948 10612 66958
rect 10556 66946 11284 66948
rect 10556 66894 10558 66946
rect 10610 66894 11284 66946
rect 10556 66892 11284 66894
rect 10556 66882 10612 66892
rect 10108 66210 10164 66220
rect 8652 66164 8708 66174
rect 8652 66162 8820 66164
rect 8652 66110 8654 66162
rect 8706 66110 8820 66162
rect 8652 66108 8820 66110
rect 8652 66098 8708 66108
rect 8652 65380 8708 65390
rect 8652 65286 8708 65324
rect 8764 64820 8820 66108
rect 11116 65492 11172 65502
rect 11004 65490 11172 65492
rect 11004 65438 11118 65490
rect 11170 65438 11172 65490
rect 11004 65436 11172 65438
rect 10108 65378 10164 65390
rect 10108 65326 10110 65378
rect 10162 65326 10164 65378
rect 8988 65266 9044 65278
rect 8988 65214 8990 65266
rect 9042 65214 9044 65266
rect 8876 64820 8932 64830
rect 8764 64818 8932 64820
rect 8764 64766 8878 64818
rect 8930 64766 8932 64818
rect 8764 64764 8932 64766
rect 8876 64754 8932 64764
rect 8988 64706 9044 65214
rect 9324 64932 9380 64942
rect 9884 64932 9940 64942
rect 9324 64930 9940 64932
rect 9324 64878 9326 64930
rect 9378 64878 9886 64930
rect 9938 64878 9940 64930
rect 9324 64876 9940 64878
rect 9324 64866 9380 64876
rect 9884 64866 9940 64876
rect 8988 64654 8990 64706
rect 9042 64654 9044 64706
rect 8988 64642 9044 64654
rect 9548 64708 9604 64718
rect 9548 64614 9604 64652
rect 9884 64706 9940 64718
rect 9884 64654 9886 64706
rect 9938 64654 9940 64706
rect 8764 64596 8820 64606
rect 8764 64502 8820 64540
rect 8316 64316 8820 64372
rect 7644 57782 7700 57820
rect 7756 62132 7924 62188
rect 8204 62356 8260 62366
rect 7644 56868 7700 56878
rect 7644 56774 7700 56812
rect 7756 56194 7812 62132
rect 7868 61796 7924 61806
rect 7868 60786 7924 61740
rect 7868 60734 7870 60786
rect 7922 60734 7924 60786
rect 7868 60722 7924 60734
rect 8092 60452 8148 60462
rect 7868 60116 7924 60126
rect 7868 60114 8036 60116
rect 7868 60062 7870 60114
rect 7922 60062 8036 60114
rect 7868 60060 8036 60062
rect 7868 60050 7924 60060
rect 7980 59220 8036 60060
rect 8092 59442 8148 60396
rect 8092 59390 8094 59442
rect 8146 59390 8148 59442
rect 8092 59378 8148 59390
rect 7868 59106 7924 59118
rect 7868 59054 7870 59106
rect 7922 59054 7924 59106
rect 7868 58996 7924 59054
rect 7868 58930 7924 58940
rect 7868 58100 7924 58110
rect 7980 58100 8036 59164
rect 8204 58324 8260 62300
rect 8428 62354 8484 62366
rect 8428 62302 8430 62354
rect 8482 62302 8484 62354
rect 8428 61796 8484 62302
rect 8428 61730 8484 61740
rect 8652 62356 8708 62366
rect 8652 61012 8708 62300
rect 8316 61010 8708 61012
rect 8316 60958 8654 61010
rect 8706 60958 8708 61010
rect 8316 60956 8708 60958
rect 8316 59218 8372 60956
rect 8652 60946 8708 60956
rect 8428 60788 8484 60798
rect 8428 60786 8596 60788
rect 8428 60734 8430 60786
rect 8482 60734 8596 60786
rect 8428 60732 8596 60734
rect 8428 60722 8484 60732
rect 8316 59166 8318 59218
rect 8370 59166 8372 59218
rect 8316 59154 8372 59166
rect 8316 58324 8372 58334
rect 8204 58268 8316 58324
rect 8316 58230 8372 58268
rect 8428 58322 8484 58334
rect 8428 58270 8430 58322
rect 8482 58270 8484 58322
rect 7924 58044 8036 58100
rect 8092 58210 8148 58222
rect 8092 58158 8094 58210
rect 8146 58158 8148 58210
rect 7868 58034 7924 58044
rect 8092 57876 8148 58158
rect 8428 57988 8484 58270
rect 8428 57922 8484 57932
rect 8092 57810 8148 57820
rect 8540 57764 8596 60732
rect 8652 59444 8708 59454
rect 8652 58884 8708 59388
rect 8652 58268 8708 58828
rect 8764 58660 8820 64316
rect 8988 64148 9044 64158
rect 8988 64054 9044 64092
rect 9884 64148 9940 64654
rect 10108 64708 10164 65326
rect 10556 65378 10612 65390
rect 10556 65326 10558 65378
rect 10610 65326 10612 65378
rect 10556 64708 10612 65326
rect 10892 65380 10948 65390
rect 10892 65044 10948 65324
rect 10892 64978 10948 64988
rect 10780 64820 10836 64830
rect 10108 64642 10164 64652
rect 10332 64652 10612 64708
rect 10668 64708 10724 64718
rect 9884 64082 9940 64092
rect 10220 64596 10276 64606
rect 10332 64596 10388 64652
rect 10276 64540 10388 64596
rect 9772 63924 9828 63934
rect 10220 63924 10276 64540
rect 10556 64482 10612 64494
rect 10556 64430 10558 64482
rect 10610 64430 10612 64482
rect 10332 64372 10388 64382
rect 10332 64146 10388 64316
rect 10556 64260 10612 64430
rect 10556 64194 10612 64204
rect 10332 64094 10334 64146
rect 10386 64094 10388 64146
rect 10332 64082 10388 64094
rect 9772 63922 10276 63924
rect 9772 63870 9774 63922
rect 9826 63870 10276 63922
rect 9772 63868 10276 63870
rect 9772 63858 9828 63868
rect 8988 62244 9044 62254
rect 8988 62150 9044 62188
rect 10108 62244 10164 63868
rect 10444 62580 10500 62590
rect 10444 62354 10500 62524
rect 10668 62468 10724 64652
rect 10780 64594 10836 64764
rect 10780 64542 10782 64594
rect 10834 64542 10836 64594
rect 10780 64530 10836 64542
rect 10892 64594 10948 64606
rect 10892 64542 10894 64594
rect 10946 64542 10948 64594
rect 10780 64036 10836 64074
rect 10780 63970 10836 63980
rect 10892 63924 10948 64542
rect 11004 64146 11060 65436
rect 11116 65426 11172 65436
rect 11228 65268 11284 66892
rect 11340 65490 11396 70812
rect 11340 65438 11342 65490
rect 11394 65438 11396 65490
rect 11340 65426 11396 65438
rect 11452 70644 11508 70654
rect 11228 65212 11396 65268
rect 11340 64818 11396 65212
rect 11340 64766 11342 64818
rect 11394 64766 11396 64818
rect 11340 64754 11396 64766
rect 11116 64706 11172 64718
rect 11116 64654 11118 64706
rect 11170 64654 11172 64706
rect 11116 64260 11172 64654
rect 11116 64194 11172 64204
rect 11228 64372 11284 64382
rect 11004 64094 11006 64146
rect 11058 64094 11060 64146
rect 11004 64082 11060 64094
rect 11228 64146 11284 64316
rect 11452 64260 11508 70588
rect 11788 70308 11844 70812
rect 12796 70588 12852 71038
rect 12572 70532 12852 70588
rect 12908 72324 12964 72334
rect 11788 70242 11844 70252
rect 12460 70420 12516 70430
rect 12460 70194 12516 70364
rect 12460 70142 12462 70194
rect 12514 70142 12516 70194
rect 12460 70130 12516 70142
rect 12012 69524 12068 69534
rect 11900 69468 12012 69524
rect 11676 67396 11732 67406
rect 11732 67340 11844 67396
rect 11676 67330 11732 67340
rect 11788 65940 11844 67340
rect 11900 66162 11956 69468
rect 12012 69458 12068 69468
rect 12572 66724 12628 70532
rect 12796 69524 12852 69534
rect 12796 69430 12852 69468
rect 12908 67060 12964 72268
rect 13692 70978 13748 70990
rect 13692 70926 13694 70978
rect 13746 70926 13748 70978
rect 13692 70420 13748 70926
rect 13692 70354 13748 70364
rect 14140 70196 14196 73276
rect 14476 73218 14532 73230
rect 14476 73166 14478 73218
rect 14530 73166 14532 73218
rect 14476 71092 14532 73166
rect 14476 71036 14756 71092
rect 14476 70868 14532 70878
rect 14476 70866 14644 70868
rect 14476 70814 14478 70866
rect 14530 70814 14644 70866
rect 14476 70812 14644 70814
rect 14476 70802 14532 70812
rect 13132 70082 13188 70094
rect 13132 70030 13134 70082
rect 13186 70030 13188 70082
rect 13132 67956 13188 70030
rect 14140 69410 14196 70140
rect 14140 69358 14142 69410
rect 14194 69358 14196 69410
rect 14140 69346 14196 69358
rect 13132 67900 13524 67956
rect 12684 67004 13188 67060
rect 12684 66946 12740 67004
rect 12684 66894 12686 66946
rect 12738 66894 12740 66946
rect 12684 66882 12740 66894
rect 12572 66668 12740 66724
rect 12236 66500 12292 66510
rect 12236 66498 12516 66500
rect 12236 66446 12238 66498
rect 12290 66446 12516 66498
rect 12236 66444 12516 66446
rect 12236 66434 12292 66444
rect 11900 66110 11902 66162
rect 11954 66110 11956 66162
rect 11900 66052 11956 66110
rect 12236 66164 12292 66174
rect 12236 66052 12292 66108
rect 11900 65996 12292 66052
rect 12348 66162 12404 66174
rect 12348 66110 12350 66162
rect 12402 66110 12404 66162
rect 11788 65884 12292 65940
rect 11564 65490 11620 65502
rect 11564 65438 11566 65490
rect 11618 65438 11620 65490
rect 11564 64932 11620 65438
rect 11564 64866 11620 64876
rect 11788 65492 11844 65502
rect 11564 64596 11620 64606
rect 11564 64502 11620 64540
rect 11788 64594 11844 65436
rect 12012 65490 12068 65502
rect 12012 65438 12014 65490
rect 12066 65438 12068 65490
rect 12012 65156 12068 65438
rect 12236 65490 12292 65884
rect 12236 65438 12238 65490
rect 12290 65438 12292 65490
rect 12236 65426 12292 65438
rect 12348 65268 12404 66110
rect 12460 65602 12516 66444
rect 12460 65550 12462 65602
rect 12514 65550 12516 65602
rect 12460 65538 12516 65550
rect 12572 65492 12628 65502
rect 12572 65398 12628 65436
rect 12348 65202 12404 65212
rect 12012 65100 12180 65156
rect 12012 64932 12068 64942
rect 12012 64706 12068 64876
rect 12012 64654 12014 64706
rect 12066 64654 12068 64706
rect 12012 64642 12068 64654
rect 11788 64542 11790 64594
rect 11842 64542 11844 64594
rect 11788 64372 11844 64542
rect 11788 64316 11956 64372
rect 11452 64194 11508 64204
rect 11228 64094 11230 64146
rect 11282 64094 11284 64146
rect 11228 64082 11284 64094
rect 11788 64036 11844 64046
rect 11788 63942 11844 63980
rect 11340 63924 11396 63934
rect 11676 63924 11732 63934
rect 10892 63922 11732 63924
rect 10892 63870 11342 63922
rect 11394 63870 11678 63922
rect 11730 63870 11732 63922
rect 10892 63868 11732 63870
rect 10780 63812 10836 63822
rect 10836 63756 10948 63812
rect 10780 63746 10836 63756
rect 10668 62466 10836 62468
rect 10668 62414 10670 62466
rect 10722 62414 10836 62466
rect 10668 62412 10836 62414
rect 10668 62402 10724 62412
rect 10444 62302 10446 62354
rect 10498 62302 10500 62354
rect 10444 62290 10500 62302
rect 10108 62178 10164 62188
rect 10108 61570 10164 61582
rect 10108 61518 10110 61570
rect 10162 61518 10164 61570
rect 9436 61458 9492 61470
rect 9436 61406 9438 61458
rect 9490 61406 9492 61458
rect 9100 59106 9156 59118
rect 9100 59054 9102 59106
rect 9154 59054 9156 59106
rect 9100 58828 9156 59054
rect 9436 58996 9492 61406
rect 9660 60788 9716 60798
rect 9660 60694 9716 60732
rect 10108 60452 10164 61518
rect 10108 60386 10164 60396
rect 10668 60452 10724 60462
rect 10668 60002 10724 60396
rect 10668 59950 10670 60002
rect 10722 59950 10724 60002
rect 10668 59938 10724 59950
rect 9996 59892 10052 59902
rect 9884 59890 10052 59892
rect 9884 59838 9998 59890
rect 10050 59838 10052 59890
rect 9884 59836 10052 59838
rect 9548 59220 9604 59230
rect 9548 59126 9604 59164
rect 9436 58940 9716 58996
rect 8764 58594 8820 58604
rect 8876 58772 9604 58828
rect 8764 58436 8820 58446
rect 8876 58436 8932 58772
rect 9436 58660 9492 58670
rect 8764 58434 8932 58436
rect 8764 58382 8766 58434
rect 8818 58382 8932 58434
rect 8764 58380 8932 58382
rect 9100 58436 9156 58446
rect 9100 58434 9380 58436
rect 9100 58382 9102 58434
rect 9154 58382 9380 58434
rect 9100 58380 9380 58382
rect 8764 58370 8820 58380
rect 9100 58370 9156 58380
rect 8652 58212 8932 58268
rect 8876 58210 8932 58212
rect 8876 58158 8878 58210
rect 8930 58158 8932 58210
rect 8428 57708 8596 57764
rect 8764 57764 8820 57802
rect 8092 57538 8148 57550
rect 8092 57486 8094 57538
rect 8146 57486 8148 57538
rect 7980 56868 8036 56878
rect 8092 56868 8148 57486
rect 7980 56866 8092 56868
rect 7980 56814 7982 56866
rect 8034 56814 8092 56866
rect 7980 56812 8092 56814
rect 8428 56868 8484 57708
rect 8764 57698 8820 57708
rect 8764 57540 8820 57578
rect 8764 57474 8820 57484
rect 8540 57428 8596 57438
rect 8540 57334 8596 57372
rect 8876 57204 8932 58158
rect 9212 58210 9268 58222
rect 9212 58158 9214 58210
rect 9266 58158 9268 58210
rect 8988 57204 9044 57214
rect 8876 57148 8988 57204
rect 8988 57138 9044 57148
rect 8988 56868 9044 56878
rect 8428 56812 8708 56868
rect 7756 56142 7758 56194
rect 7810 56142 7812 56194
rect 7756 55298 7812 56142
rect 7868 56754 7924 56766
rect 7868 56702 7870 56754
rect 7922 56702 7924 56754
rect 7868 55860 7924 56702
rect 7868 55794 7924 55804
rect 7756 55246 7758 55298
rect 7810 55246 7812 55298
rect 7756 55234 7812 55246
rect 6860 53340 7252 53396
rect 6748 53228 6916 53284
rect 6188 52948 6244 52958
rect 6188 52946 6692 52948
rect 6188 52894 6190 52946
rect 6242 52894 6692 52946
rect 6188 52892 6692 52894
rect 6188 52882 6244 52892
rect 6300 52724 6356 52734
rect 6188 52388 6244 52398
rect 6188 52274 6244 52332
rect 6188 52222 6190 52274
rect 6242 52222 6244 52274
rect 6188 52210 6244 52222
rect 6300 52052 6356 52668
rect 6636 52274 6692 52892
rect 6748 52834 6804 52846
rect 6748 52782 6750 52834
rect 6802 52782 6804 52834
rect 6748 52724 6804 52782
rect 6748 52658 6804 52668
rect 6636 52222 6638 52274
rect 6690 52222 6692 52274
rect 6636 52210 6692 52222
rect 6300 51378 6356 51996
rect 6300 51326 6302 51378
rect 6354 51326 6356 51378
rect 6300 51314 6356 51326
rect 6524 52050 6580 52062
rect 6524 51998 6526 52050
rect 6578 51998 6580 52050
rect 6524 51380 6580 51998
rect 6748 52052 6804 52062
rect 6860 52052 6916 53228
rect 7196 52162 7252 53340
rect 7196 52110 7198 52162
rect 7250 52110 7252 52162
rect 7196 52098 7252 52110
rect 7308 53340 7588 53396
rect 6860 51996 7028 52052
rect 6748 51958 6804 51996
rect 6188 51044 6244 51054
rect 6076 50988 6188 51044
rect 6188 50978 6244 50988
rect 6524 50706 6580 51324
rect 6524 50654 6526 50706
rect 6578 50654 6580 50706
rect 6524 50428 6580 50654
rect 5516 50372 5684 50428
rect 5740 50372 6020 50428
rect 5516 49698 5572 49710
rect 5516 49646 5518 49698
rect 5570 49646 5572 49698
rect 5516 49476 5572 49646
rect 5516 49410 5572 49420
rect 5404 47058 5460 47068
rect 5404 46788 5460 46798
rect 5404 46694 5460 46732
rect 5628 45892 5684 50372
rect 5852 49588 5908 49598
rect 5740 46788 5796 46798
rect 5740 46694 5796 46732
rect 5852 46340 5908 49532
rect 5740 45892 5796 45902
rect 5628 45836 5740 45892
rect 5740 45798 5796 45836
rect 5292 45052 5796 45108
rect 5292 43650 5348 45052
rect 5740 44434 5796 45052
rect 5740 44382 5742 44434
rect 5794 44382 5796 44434
rect 5740 44370 5796 44382
rect 5852 44212 5908 46284
rect 5740 44156 5908 44212
rect 5516 44100 5572 44110
rect 5292 43598 5294 43650
rect 5346 43598 5348 43650
rect 5292 43586 5348 43598
rect 5404 43650 5460 43662
rect 5404 43598 5406 43650
rect 5458 43598 5460 43650
rect 5404 42868 5460 43598
rect 5404 42802 5460 42812
rect 5404 42532 5460 42542
rect 5180 42466 5236 42476
rect 5292 42476 5404 42532
rect 5516 42532 5572 44044
rect 5628 43538 5684 43550
rect 5628 43486 5630 43538
rect 5682 43486 5684 43538
rect 5628 42756 5684 43486
rect 5740 43092 5796 44156
rect 5740 43026 5796 43036
rect 5852 43650 5908 43662
rect 5852 43598 5854 43650
rect 5906 43598 5908 43650
rect 5852 43540 5908 43598
rect 5628 42662 5684 42700
rect 5740 42532 5796 42570
rect 5516 42476 5684 42532
rect 5292 42084 5348 42476
rect 5404 42466 5460 42476
rect 5068 42028 5348 42084
rect 5068 41970 5124 42028
rect 5068 41918 5070 41970
rect 5122 41918 5124 41970
rect 5068 41906 5124 41918
rect 5516 41858 5572 41870
rect 5516 41806 5518 41858
rect 5570 41806 5572 41858
rect 5068 41748 5124 41758
rect 5068 41746 5236 41748
rect 5068 41694 5070 41746
rect 5122 41694 5236 41746
rect 5068 41692 5236 41694
rect 5068 41682 5124 41692
rect 5068 41076 5124 41086
rect 4956 41020 5068 41076
rect 5068 41010 5124 41020
rect 4732 40628 4788 40638
rect 4732 40534 4788 40572
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4620 39730 4676 39742
rect 4620 39678 4622 39730
rect 4674 39678 4676 39730
rect 4284 39508 4340 39518
rect 4284 38612 4340 39452
rect 4620 39060 4676 39678
rect 4620 38994 4676 39004
rect 4844 38948 4900 38958
rect 4844 38668 4900 38892
rect 4844 38612 5012 38668
rect 4284 38546 4340 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4396 37268 4452 37278
rect 4396 37174 4452 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4396 36708 4452 36718
rect 4396 36596 4452 36652
rect 4396 36594 4564 36596
rect 4396 36542 4398 36594
rect 4450 36542 4564 36594
rect 4396 36540 4564 36542
rect 4396 36530 4452 36540
rect 4508 36482 4564 36540
rect 4508 36430 4510 36482
rect 4562 36430 4564 36482
rect 4508 36418 4564 36430
rect 4956 36372 5012 38612
rect 5068 38610 5124 38622
rect 5068 38558 5070 38610
rect 5122 38558 5124 38610
rect 5068 37378 5124 38558
rect 5068 37326 5070 37378
rect 5122 37326 5124 37378
rect 5068 37314 5124 37326
rect 5180 36820 5236 41692
rect 5516 41636 5572 41806
rect 5516 40628 5572 41580
rect 5516 40534 5572 40572
rect 5628 40404 5684 42476
rect 5740 42466 5796 42476
rect 5852 42530 5908 43484
rect 5852 42478 5854 42530
rect 5906 42478 5908 42530
rect 5852 42466 5908 42478
rect 5740 40404 5796 40414
rect 5628 40402 5796 40404
rect 5628 40350 5742 40402
rect 5794 40350 5796 40402
rect 5628 40348 5796 40350
rect 5740 40338 5796 40348
rect 5964 40180 6020 50372
rect 6412 50372 6580 50428
rect 6860 50708 6916 50718
rect 6076 48468 6132 48478
rect 6076 48374 6132 48412
rect 6412 48354 6468 50372
rect 6860 49922 6916 50652
rect 6860 49870 6862 49922
rect 6914 49870 6916 49922
rect 6860 49858 6916 49870
rect 6412 48302 6414 48354
rect 6466 48302 6468 48354
rect 6412 48290 6468 48302
rect 6636 49810 6692 49822
rect 6636 49758 6638 49810
rect 6690 49758 6692 49810
rect 6636 49476 6692 49758
rect 6636 48468 6692 49420
rect 6636 48242 6692 48412
rect 6636 48190 6638 48242
rect 6690 48190 6692 48242
rect 6636 48178 6692 48190
rect 6748 46900 6804 46910
rect 6076 46788 6132 46798
rect 6076 46786 6468 46788
rect 6076 46734 6078 46786
rect 6130 46734 6468 46786
rect 6076 46732 6468 46734
rect 6076 46722 6132 46732
rect 6412 46002 6468 46732
rect 6412 45950 6414 46002
rect 6466 45950 6468 46002
rect 6412 45938 6468 45950
rect 6748 45332 6804 46844
rect 6300 45276 6804 45332
rect 6860 45332 6916 45342
rect 6300 44436 6356 45276
rect 6300 44342 6356 44380
rect 6524 44210 6580 44222
rect 6524 44158 6526 44210
rect 6578 44158 6580 44210
rect 6524 44100 6580 44158
rect 6524 44034 6580 44044
rect 6636 44098 6692 44110
rect 6636 44046 6638 44098
rect 6690 44046 6692 44098
rect 6636 43876 6692 44046
rect 6636 43810 6692 43820
rect 6860 44098 6916 45276
rect 6860 44046 6862 44098
rect 6914 44046 6916 44098
rect 6636 43650 6692 43662
rect 6636 43598 6638 43650
rect 6690 43598 6692 43650
rect 6188 43540 6244 43550
rect 6636 43540 6692 43598
rect 6860 43650 6916 44046
rect 6860 43598 6862 43650
rect 6914 43598 6916 43650
rect 6860 43586 6916 43598
rect 6188 43538 6580 43540
rect 6188 43486 6190 43538
rect 6242 43486 6580 43538
rect 6188 43484 6580 43486
rect 6188 43474 6244 43484
rect 6188 43092 6244 43102
rect 6188 42308 6244 43036
rect 6524 42980 6580 43484
rect 6636 43474 6692 43484
rect 6748 43426 6804 43438
rect 6748 43374 6750 43426
rect 6802 43374 6804 43426
rect 6636 42980 6692 42990
rect 6524 42978 6692 42980
rect 6524 42926 6638 42978
rect 6690 42926 6692 42978
rect 6524 42924 6692 42926
rect 6636 42756 6692 42924
rect 6636 42690 6692 42700
rect 6524 42644 6580 42654
rect 6076 42252 6244 42308
rect 6412 42642 6580 42644
rect 6412 42590 6526 42642
rect 6578 42590 6580 42642
rect 6412 42588 6580 42590
rect 6076 41412 6132 42252
rect 6188 41860 6244 41870
rect 6412 41860 6468 42588
rect 6524 42578 6580 42588
rect 6748 42420 6804 43374
rect 6972 43092 7028 51996
rect 7308 51490 7364 53340
rect 7532 53172 7588 53182
rect 7532 53078 7588 53116
rect 7308 51438 7310 51490
rect 7362 51438 7364 51490
rect 7308 50708 7364 51438
rect 7644 51380 7700 51390
rect 7308 50652 7588 50708
rect 7532 50594 7588 50652
rect 7532 50542 7534 50594
rect 7586 50542 7588 50594
rect 7532 50530 7588 50542
rect 7644 50484 7700 51324
rect 7644 50418 7700 50428
rect 7756 51044 7812 51054
rect 7756 49810 7812 50988
rect 7756 49758 7758 49810
rect 7810 49758 7812 49810
rect 7756 49746 7812 49758
rect 7868 50034 7924 50046
rect 7868 49982 7870 50034
rect 7922 49982 7924 50034
rect 7196 49026 7252 49038
rect 7196 48974 7198 49026
rect 7250 48974 7252 49026
rect 7196 48244 7252 48974
rect 7644 49028 7700 49038
rect 7868 49028 7924 49982
rect 7644 49026 7924 49028
rect 7644 48974 7646 49026
rect 7698 48974 7924 49026
rect 7644 48972 7924 48974
rect 7532 48916 7588 48926
rect 7196 48178 7252 48188
rect 7420 48914 7588 48916
rect 7420 48862 7534 48914
rect 7586 48862 7588 48914
rect 7420 48860 7588 48862
rect 7084 45332 7140 45342
rect 7084 44100 7140 45276
rect 7420 44996 7476 48860
rect 7532 48850 7588 48860
rect 7644 47458 7700 48972
rect 7980 48916 8036 56812
rect 8092 56774 8148 56812
rect 8428 56642 8484 56654
rect 8428 56590 8430 56642
rect 8482 56590 8484 56642
rect 8204 55860 8260 55870
rect 8316 55860 8372 55870
rect 8260 55858 8372 55860
rect 8260 55806 8318 55858
rect 8370 55806 8372 55858
rect 8260 55804 8372 55806
rect 8092 54516 8148 54526
rect 8092 54422 8148 54460
rect 8092 52834 8148 52846
rect 8092 52782 8094 52834
rect 8146 52782 8148 52834
rect 8092 52500 8148 52782
rect 8092 52434 8148 52444
rect 8204 50428 8260 55804
rect 8316 55794 8372 55804
rect 8428 54404 8484 56590
rect 8540 54740 8596 54750
rect 8540 54646 8596 54684
rect 8428 54338 8484 54348
rect 8316 53506 8372 53518
rect 8316 53454 8318 53506
rect 8370 53454 8372 53506
rect 8316 52162 8372 53454
rect 8428 52834 8484 52846
rect 8428 52782 8430 52834
rect 8482 52782 8484 52834
rect 8428 52724 8484 52782
rect 8428 52658 8484 52668
rect 8316 52110 8318 52162
rect 8370 52110 8372 52162
rect 8316 52052 8372 52110
rect 8372 51996 8596 52052
rect 8316 51986 8372 51996
rect 8540 51604 8596 51996
rect 8652 51940 8708 56812
rect 8988 56774 9044 56812
rect 9212 56866 9268 58158
rect 9324 57652 9380 58380
rect 9436 58322 9492 58604
rect 9436 58270 9438 58322
rect 9490 58270 9492 58322
rect 9436 58258 9492 58270
rect 9548 58322 9604 58772
rect 9548 58270 9550 58322
rect 9602 58270 9604 58322
rect 9548 58100 9604 58270
rect 9548 58034 9604 58044
rect 9660 57874 9716 58940
rect 9660 57822 9662 57874
rect 9714 57822 9716 57874
rect 9660 57810 9716 57822
rect 9772 58210 9828 58222
rect 9772 58158 9774 58210
rect 9826 58158 9828 58210
rect 9436 57652 9492 57662
rect 9324 57650 9492 57652
rect 9324 57598 9438 57650
rect 9490 57598 9492 57650
rect 9324 57596 9492 57598
rect 9436 57586 9492 57596
rect 9212 56814 9214 56866
rect 9266 56814 9268 56866
rect 9212 56802 9268 56814
rect 9660 56868 9716 56878
rect 9772 56868 9828 58158
rect 9884 57988 9940 59836
rect 9996 59826 10052 59836
rect 9996 59108 10052 59118
rect 9996 58828 10052 59052
rect 10556 59108 10612 59118
rect 10556 59106 10724 59108
rect 10556 59054 10558 59106
rect 10610 59054 10724 59106
rect 10556 59052 10724 59054
rect 10556 59042 10612 59052
rect 10668 58996 10724 59052
rect 9996 58772 10612 58828
rect 10108 58266 10164 58278
rect 9996 58212 10052 58222
rect 9996 58118 10052 58156
rect 10108 58214 10110 58266
rect 10162 58214 10164 58266
rect 10108 57988 10164 58214
rect 10556 58212 10612 58772
rect 10668 58772 10724 58940
rect 10668 58706 10724 58716
rect 10612 58156 10724 58212
rect 10556 58118 10612 58156
rect 9884 57932 10052 57988
rect 9884 57764 9940 57774
rect 9884 57670 9940 57708
rect 9660 56866 9828 56868
rect 9660 56814 9662 56866
rect 9714 56814 9828 56866
rect 9660 56812 9828 56814
rect 9884 56868 9940 56878
rect 9660 56802 9716 56812
rect 9884 56774 9940 56812
rect 9548 56644 9604 56654
rect 9996 56644 10052 57932
rect 10108 57922 10164 57932
rect 10668 57876 10724 58156
rect 10668 57810 10724 57820
rect 10556 57762 10612 57774
rect 10556 57710 10558 57762
rect 10610 57710 10612 57762
rect 9548 56642 10052 56644
rect 9548 56590 9550 56642
rect 9602 56590 10052 56642
rect 9548 56588 10052 56590
rect 10108 57650 10164 57662
rect 10556 57652 10612 57710
rect 10108 57598 10110 57650
rect 10162 57598 10164 57650
rect 10108 57540 10164 57598
rect 9548 56578 9604 56588
rect 10108 56308 10164 57484
rect 10444 57596 10612 57652
rect 10780 57652 10836 62412
rect 10892 61348 10948 63756
rect 11116 62580 11172 62590
rect 11116 62486 11172 62524
rect 11340 62188 11396 63868
rect 11676 63858 11732 63868
rect 11900 63700 11956 64316
rect 12012 64148 12068 64158
rect 12124 64148 12180 65100
rect 12684 64932 12740 66668
rect 13020 66050 13076 66062
rect 13020 65998 13022 66050
rect 13074 65998 13076 66050
rect 13020 65828 13076 65998
rect 12236 64876 12740 64932
rect 12796 65268 12852 65278
rect 12236 64484 12292 64876
rect 12348 64764 12740 64820
rect 12348 64706 12404 64764
rect 12348 64654 12350 64706
rect 12402 64654 12404 64706
rect 12348 64642 12404 64654
rect 12684 64708 12740 64764
rect 12796 64708 12852 65212
rect 12908 64708 12964 64718
rect 12684 64706 12964 64708
rect 12684 64654 12910 64706
rect 12962 64654 12964 64706
rect 12684 64652 12964 64654
rect 12572 64596 12628 64606
rect 12572 64502 12628 64540
rect 12236 64482 12404 64484
rect 12236 64430 12238 64482
rect 12290 64430 12404 64482
rect 12236 64428 12404 64430
rect 12236 64418 12292 64428
rect 12012 64146 12180 64148
rect 12012 64094 12014 64146
rect 12066 64094 12180 64146
rect 12012 64092 12180 64094
rect 12236 64148 12292 64158
rect 12012 64082 12068 64092
rect 11900 63634 11956 63644
rect 11228 62132 11396 62188
rect 11452 62580 11508 62590
rect 11228 61572 11284 62132
rect 11228 61478 11284 61516
rect 11340 61348 11396 61358
rect 10892 61346 11396 61348
rect 10892 61294 10894 61346
rect 10946 61294 11342 61346
rect 11394 61294 11396 61346
rect 10892 61292 11396 61294
rect 10892 61282 10948 61292
rect 11228 60786 11284 60798
rect 11228 60734 11230 60786
rect 11282 60734 11284 60786
rect 11228 60452 11284 60734
rect 11228 60386 11284 60396
rect 11340 58884 11396 61292
rect 11228 58828 11396 58884
rect 11004 58210 11060 58222
rect 11004 58158 11006 58210
rect 11058 58158 11060 58210
rect 11004 58100 11060 58158
rect 10444 57540 10500 57596
rect 10780 57586 10836 57596
rect 10892 57650 10948 57662
rect 10892 57598 10894 57650
rect 10946 57598 10948 57650
rect 10444 57474 10500 57484
rect 10332 56868 10388 56878
rect 10892 56868 10948 57598
rect 10332 56642 10388 56812
rect 10332 56590 10334 56642
rect 10386 56590 10388 56642
rect 10332 56308 10388 56590
rect 9996 56252 10388 56308
rect 10444 56812 10948 56868
rect 10444 56306 10500 56812
rect 11004 56756 11060 58044
rect 10444 56254 10446 56306
rect 10498 56254 10500 56306
rect 9660 55970 9716 55982
rect 9660 55918 9662 55970
rect 9714 55918 9716 55970
rect 9660 55860 9716 55918
rect 9660 55794 9716 55804
rect 9660 55636 9716 55646
rect 8876 53172 8932 53182
rect 8764 52946 8820 52958
rect 8764 52894 8766 52946
rect 8818 52894 8820 52946
rect 8764 52500 8820 52894
rect 8876 52612 8932 53116
rect 9100 53060 9156 53070
rect 9548 53060 9604 53070
rect 9100 53058 9604 53060
rect 9100 53006 9102 53058
rect 9154 53006 9550 53058
rect 9602 53006 9604 53058
rect 9100 53004 9604 53006
rect 9100 52994 9156 53004
rect 9548 52994 9604 53004
rect 8876 52546 8932 52556
rect 9548 52836 9604 52846
rect 8764 52434 8820 52444
rect 9212 52274 9268 52286
rect 9212 52222 9214 52274
rect 9266 52222 9268 52274
rect 9100 52164 9156 52174
rect 8652 51874 8708 51884
rect 8876 52162 9156 52164
rect 8876 52110 9102 52162
rect 9154 52110 9156 52162
rect 8876 52108 9156 52110
rect 8316 51378 8372 51390
rect 8316 51326 8318 51378
rect 8370 51326 8372 51378
rect 8316 50596 8372 51326
rect 8316 50530 8372 50540
rect 8428 51266 8484 51278
rect 8428 51214 8430 51266
rect 8482 51214 8484 51266
rect 8428 50484 8484 51214
rect 8204 50372 8372 50428
rect 8428 50418 8484 50428
rect 7644 47406 7646 47458
rect 7698 47406 7700 47458
rect 7644 47394 7700 47406
rect 7756 48860 8036 48916
rect 8204 49028 8260 49038
rect 7644 47236 7700 47246
rect 7644 47142 7700 47180
rect 7532 46900 7588 46910
rect 7532 46806 7588 46844
rect 7420 44930 7476 44940
rect 7532 44994 7588 45006
rect 7532 44942 7534 44994
rect 7586 44942 7588 44994
rect 7532 44772 7588 44942
rect 7308 44716 7588 44772
rect 7084 44006 7140 44044
rect 7196 44212 7252 44222
rect 7308 44212 7364 44716
rect 7196 44210 7364 44212
rect 7196 44158 7198 44210
rect 7250 44158 7364 44210
rect 7196 44156 7364 44158
rect 7644 44436 7700 44446
rect 7084 43538 7140 43550
rect 7084 43486 7086 43538
rect 7138 43486 7140 43538
rect 7084 43428 7140 43486
rect 7084 43362 7140 43372
rect 6972 43026 7028 43036
rect 7084 42980 7140 42990
rect 7084 42886 7140 42924
rect 6972 42644 7028 42654
rect 6972 42550 7028 42588
rect 6748 42354 6804 42364
rect 6188 41858 6468 41860
rect 6188 41806 6190 41858
rect 6242 41806 6468 41858
rect 6188 41804 6468 41806
rect 6188 41636 6244 41804
rect 6188 41570 6244 41580
rect 7084 41636 7140 41646
rect 6076 41356 6356 41412
rect 5740 40124 6020 40180
rect 6076 41076 6132 41086
rect 5628 39394 5684 39406
rect 5628 39342 5630 39394
rect 5682 39342 5684 39394
rect 5404 38948 5460 38958
rect 5404 38854 5460 38892
rect 5628 38668 5684 39342
rect 5516 38612 5684 38668
rect 5740 38668 5796 40124
rect 5964 39508 6020 39518
rect 6076 39508 6132 41020
rect 5964 39506 6132 39508
rect 5964 39454 5966 39506
rect 6018 39454 6132 39506
rect 5964 39452 6132 39454
rect 5964 39442 6020 39452
rect 5740 38612 6020 38668
rect 5516 38610 5572 38612
rect 5516 38558 5518 38610
rect 5570 38558 5572 38610
rect 5516 38546 5572 38558
rect 5180 36764 5348 36820
rect 5292 36484 5348 36764
rect 5852 36484 5908 36494
rect 5292 36482 5908 36484
rect 5292 36430 5854 36482
rect 5906 36430 5908 36482
rect 5292 36428 5908 36430
rect 5068 36372 5124 36382
rect 4956 36316 5068 36372
rect 5068 36278 5124 36316
rect 4844 36258 4900 36270
rect 4844 36206 4846 36258
rect 4898 36206 4900 36258
rect 4620 35588 4676 35598
rect 4844 35588 4900 36206
rect 5180 36260 5236 36270
rect 5180 36166 5236 36204
rect 5292 35810 5348 36428
rect 5852 36418 5908 36428
rect 5292 35758 5294 35810
rect 5346 35758 5348 35810
rect 5292 35746 5348 35758
rect 5628 36258 5684 36270
rect 5628 36206 5630 36258
rect 5682 36206 5684 36258
rect 4284 35586 4900 35588
rect 4284 35534 4622 35586
rect 4674 35534 4900 35586
rect 4284 35532 4900 35534
rect 4956 35588 5012 35598
rect 4284 35140 4340 35532
rect 4620 35522 4676 35532
rect 4956 35494 5012 35532
rect 4956 35364 5012 35374
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35308 4956 35364
rect 4620 35140 4676 35150
rect 4844 35140 4900 35308
rect 4956 35298 5012 35308
rect 5628 35364 5684 36206
rect 5628 35298 5684 35308
rect 5740 36258 5796 36270
rect 5740 36206 5742 36258
rect 5794 36206 5796 36258
rect 4284 35084 4452 35140
rect 4284 34916 4340 34926
rect 4284 34822 4340 34860
rect 4396 34804 4452 35084
rect 4620 35138 4900 35140
rect 4620 35086 4622 35138
rect 4674 35086 4900 35138
rect 4620 35084 4900 35086
rect 4620 35074 4676 35084
rect 5068 35028 5124 35038
rect 5068 34934 5124 34972
rect 5740 34916 5796 36206
rect 5964 35140 6020 38612
rect 6076 36260 6132 36270
rect 6076 36166 6132 36204
rect 5964 35084 6132 35140
rect 4396 34738 4452 34748
rect 5516 34860 5796 34916
rect 5964 34916 6020 34926
rect 4284 34356 4340 34366
rect 4172 34354 4340 34356
rect 4172 34302 4286 34354
rect 4338 34302 4340 34354
rect 4172 34300 4340 34302
rect 4284 34244 4340 34300
rect 4620 34356 4676 34366
rect 4620 34262 4676 34300
rect 5068 34356 5124 34366
rect 4284 34178 4340 34188
rect 5068 34130 5124 34300
rect 5180 34244 5236 34254
rect 5180 34150 5236 34188
rect 5068 34078 5070 34130
rect 5122 34078 5124 34130
rect 5068 34066 5124 34078
rect 4732 34020 4788 34030
rect 4788 33964 4900 34020
rect 4732 33954 4788 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33460 4340 33470
rect 4844 33460 4900 33964
rect 4284 32788 4340 33404
rect 4284 32694 4340 32732
rect 4732 33404 4900 33460
rect 4732 32786 4788 33404
rect 4732 32734 4734 32786
rect 4786 32734 4788 32786
rect 4732 32722 4788 32734
rect 4844 33236 4900 33246
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 32004 4900 33180
rect 4732 31948 4900 32004
rect 5068 32450 5124 32462
rect 5068 32398 5070 32450
rect 5122 32398 5124 32450
rect 4620 31554 4676 31566
rect 4620 31502 4622 31554
rect 4674 31502 4676 31554
rect 4620 31444 4676 31502
rect 4284 31388 4620 31444
rect 4284 30436 4340 31388
rect 4620 31350 4676 31388
rect 4620 30884 4676 30894
rect 4732 30884 4788 31948
rect 5068 31780 5124 32398
rect 4620 30882 4788 30884
rect 4620 30830 4622 30882
rect 4674 30830 4788 30882
rect 4620 30828 4788 30830
rect 4844 31724 5124 31780
rect 4844 31666 4900 31724
rect 4844 31614 4846 31666
rect 4898 31614 4900 31666
rect 4844 30996 4900 31614
rect 4956 31554 5012 31566
rect 4956 31502 4958 31554
rect 5010 31502 5012 31554
rect 4956 31444 5012 31502
rect 5180 31556 5236 31566
rect 5180 31554 5460 31556
rect 5180 31502 5182 31554
rect 5234 31502 5460 31554
rect 5180 31500 5460 31502
rect 5180 31490 5236 31500
rect 4956 31378 5012 31388
rect 4620 30818 4676 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30380 4452 30436
rect 4396 30210 4452 30380
rect 4508 30324 4564 30334
rect 4844 30324 4900 30940
rect 4956 30884 5012 30894
rect 4956 30790 5012 30828
rect 4508 30322 4900 30324
rect 4508 30270 4510 30322
rect 4562 30270 4900 30322
rect 4508 30268 4900 30270
rect 4508 30258 4564 30268
rect 4396 30158 4398 30210
rect 4450 30158 4452 30210
rect 4284 30098 4340 30110
rect 4284 30046 4286 30098
rect 4338 30046 4340 30098
rect 4060 26964 4116 27002
rect 4060 26898 4116 26908
rect 4284 25618 4340 30046
rect 4396 29652 4452 30158
rect 5180 30212 5236 30222
rect 5180 30118 5236 30156
rect 5404 30100 5460 31500
rect 5516 30994 5572 34860
rect 5964 34822 6020 34860
rect 5740 34692 5796 34702
rect 5740 34598 5796 34636
rect 5740 34242 5796 34254
rect 5740 34190 5742 34242
rect 5794 34190 5796 34242
rect 5740 33236 5796 34190
rect 5964 33348 6020 33358
rect 5740 33142 5796 33180
rect 5852 33346 6020 33348
rect 5852 33294 5966 33346
rect 6018 33294 6020 33346
rect 5852 33292 6020 33294
rect 5628 32562 5684 32574
rect 5628 32510 5630 32562
rect 5682 32510 5684 32562
rect 5628 31668 5684 32510
rect 5628 31612 5796 31668
rect 5740 31444 5796 31612
rect 5740 31378 5796 31388
rect 5516 30942 5518 30994
rect 5570 30942 5572 30994
rect 5516 30660 5572 30942
rect 5516 30594 5572 30604
rect 5404 30044 5684 30100
rect 4396 29586 4452 29596
rect 5404 29652 5460 29662
rect 5404 29558 5460 29596
rect 5628 29538 5684 30044
rect 5740 29986 5796 29998
rect 5740 29934 5742 29986
rect 5794 29934 5796 29986
rect 5740 29876 5796 29934
rect 5740 29810 5796 29820
rect 5628 29486 5630 29538
rect 5682 29486 5684 29538
rect 5628 29474 5684 29486
rect 5740 29540 5796 29550
rect 5740 29446 5796 29484
rect 4844 29316 4900 29326
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4620 28756 4676 28766
rect 4620 28662 4676 28700
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 26404 4900 29260
rect 5740 29092 5796 29102
rect 5628 29036 5740 29092
rect 5068 28644 5124 28654
rect 4956 26964 5012 26974
rect 4956 26516 5012 26908
rect 5068 26908 5124 28588
rect 5628 28420 5684 29036
rect 5740 29026 5796 29036
rect 5852 28756 5908 33292
rect 5964 33282 6020 33292
rect 6076 32564 6132 35084
rect 6188 34914 6244 34926
rect 6188 34862 6190 34914
rect 6242 34862 6244 34914
rect 6188 34580 6244 34862
rect 6188 34356 6244 34524
rect 6188 34290 6244 34300
rect 6076 32498 6132 32508
rect 6188 34018 6244 34030
rect 6188 33966 6190 34018
rect 6242 33966 6244 34018
rect 5964 32340 6020 32350
rect 5964 32246 6020 32284
rect 5964 31556 6020 31566
rect 6076 31556 6132 31566
rect 5964 31554 6076 31556
rect 5964 31502 5966 31554
rect 6018 31502 6076 31554
rect 5964 31500 6076 31502
rect 5964 31490 6020 31500
rect 5964 30212 6020 30222
rect 5964 29650 6020 30156
rect 5964 29598 5966 29650
rect 6018 29598 6020 29650
rect 5964 29586 6020 29598
rect 6076 29876 6132 31500
rect 6188 31444 6244 33966
rect 6300 33460 6356 41356
rect 6748 41298 6804 41310
rect 6748 41246 6750 41298
rect 6802 41246 6804 41298
rect 6748 41076 6804 41246
rect 6748 41010 6804 41020
rect 7084 40516 7140 41580
rect 7196 40962 7252 44156
rect 7644 43538 7700 44380
rect 7644 43486 7646 43538
rect 7698 43486 7700 43538
rect 7644 43474 7700 43486
rect 7532 43426 7588 43438
rect 7532 43374 7534 43426
rect 7586 43374 7588 43426
rect 7308 42756 7364 42766
rect 7308 42662 7364 42700
rect 7308 42420 7364 42430
rect 7364 42364 7476 42420
rect 7308 42354 7364 42364
rect 7196 40910 7198 40962
rect 7250 40910 7252 40962
rect 7196 40852 7252 40910
rect 7196 40786 7252 40796
rect 7196 40516 7252 40526
rect 7084 40514 7252 40516
rect 7084 40462 7198 40514
rect 7250 40462 7252 40514
rect 7084 40460 7252 40462
rect 7196 40450 7252 40460
rect 6748 40178 6804 40190
rect 6748 40126 6750 40178
rect 6802 40126 6804 40178
rect 6748 39620 6804 40126
rect 6860 39844 6916 39854
rect 7420 39844 7476 42364
rect 7532 40068 7588 43374
rect 7756 42868 7812 48860
rect 8204 48692 8260 48972
rect 7980 48636 8260 48692
rect 7980 47346 8036 48636
rect 8204 48244 8260 48254
rect 8204 47460 8260 48188
rect 8204 47394 8260 47404
rect 7980 47294 7982 47346
rect 8034 47294 8036 47346
rect 7980 47282 8036 47294
rect 8316 47124 8372 50372
rect 8540 49922 8596 51548
rect 8540 49870 8542 49922
rect 8594 49870 8596 49922
rect 8540 49858 8596 49870
rect 8652 51716 8708 51726
rect 8540 48468 8596 48478
rect 8204 47068 8372 47124
rect 8428 48412 8540 48468
rect 7980 46562 8036 46574
rect 7980 46510 7982 46562
rect 8034 46510 8036 46562
rect 7980 45892 8036 46510
rect 7868 45108 7924 45118
rect 7868 45014 7924 45052
rect 7644 42812 7812 42868
rect 7868 44212 7924 44222
rect 7980 44212 8036 45836
rect 7868 44210 8036 44212
rect 7868 44158 7870 44210
rect 7922 44158 8036 44210
rect 7868 44156 8036 44158
rect 7644 41972 7700 42812
rect 7644 41906 7700 41916
rect 7756 42642 7812 42654
rect 7756 42590 7758 42642
rect 7810 42590 7812 42642
rect 7532 40002 7588 40012
rect 7756 39844 7812 42590
rect 7420 39788 7700 39844
rect 6860 39750 6916 39788
rect 7084 39620 7140 39630
rect 7420 39620 7476 39630
rect 6748 39618 7420 39620
rect 6748 39566 7086 39618
rect 7138 39566 7420 39618
rect 6748 39564 7420 39566
rect 7084 39554 7140 39564
rect 7420 39526 7476 39564
rect 6524 39394 6580 39406
rect 6524 39342 6526 39394
rect 6578 39342 6580 39394
rect 6524 37156 6580 39342
rect 6524 37090 6580 37100
rect 7084 39396 7140 39406
rect 6860 36708 6916 36718
rect 6860 36372 6916 36652
rect 6860 35810 6916 36316
rect 6860 35758 6862 35810
rect 6914 35758 6916 35810
rect 6860 35746 6916 35758
rect 6972 35586 7028 35598
rect 6972 35534 6974 35586
rect 7026 35534 7028 35586
rect 6860 35252 6916 35262
rect 6860 35028 6916 35196
rect 6412 34972 6916 35028
rect 6412 34244 6468 34972
rect 6636 34804 6692 34814
rect 6748 34804 6804 34814
rect 6636 34802 6748 34804
rect 6636 34750 6638 34802
rect 6690 34750 6748 34802
rect 6636 34748 6748 34750
rect 6636 34738 6692 34748
rect 6412 34178 6468 34188
rect 6300 33394 6356 33404
rect 6524 34130 6580 34142
rect 6524 34078 6526 34130
rect 6578 34078 6580 34130
rect 6524 33908 6580 34078
rect 6524 33236 6580 33852
rect 6748 33346 6804 34748
rect 6860 34802 6916 34972
rect 6860 34750 6862 34802
rect 6914 34750 6916 34802
rect 6860 34738 6916 34750
rect 6972 34916 7028 35534
rect 6972 34580 7028 34860
rect 6860 34524 7028 34580
rect 6860 34130 6916 34524
rect 6860 34078 6862 34130
rect 6914 34078 6916 34130
rect 6860 34066 6916 34078
rect 6748 33294 6750 33346
rect 6802 33294 6804 33346
rect 6748 33282 6804 33294
rect 6972 33572 7028 33582
rect 6412 33180 6580 33236
rect 6636 33234 6692 33246
rect 6636 33182 6638 33234
rect 6690 33182 6692 33234
rect 6300 32676 6356 32686
rect 6300 32562 6356 32620
rect 6300 32510 6302 32562
rect 6354 32510 6356 32562
rect 6300 32498 6356 32510
rect 6412 31890 6468 33180
rect 6524 32452 6580 32462
rect 6524 32358 6580 32396
rect 6412 31838 6414 31890
rect 6466 31838 6468 31890
rect 6412 31826 6468 31838
rect 6636 31778 6692 33182
rect 6636 31726 6638 31778
rect 6690 31726 6692 31778
rect 6636 31714 6692 31726
rect 6748 32004 6804 32014
rect 6188 31378 6244 31388
rect 6524 31444 6580 31454
rect 6412 30996 6468 31006
rect 6412 30902 6468 30940
rect 6524 30210 6580 31388
rect 6524 30158 6526 30210
rect 6578 30158 6580 30210
rect 6524 30146 6580 30158
rect 6636 30322 6692 30334
rect 6636 30270 6638 30322
rect 6690 30270 6692 30322
rect 6076 29092 6132 29820
rect 6636 29876 6692 30270
rect 6636 29810 6692 29820
rect 6076 29026 6132 29036
rect 5740 28644 5796 28654
rect 5852 28644 5908 28700
rect 5740 28642 6020 28644
rect 5740 28590 5742 28642
rect 5794 28590 6020 28642
rect 5740 28588 6020 28590
rect 5740 28578 5796 28588
rect 5740 28420 5796 28430
rect 5628 28418 5796 28420
rect 5628 28366 5742 28418
rect 5794 28366 5796 28418
rect 5628 28364 5796 28366
rect 5740 28354 5796 28364
rect 5852 26964 5908 27002
rect 5068 26852 5348 26908
rect 5852 26898 5908 26908
rect 4956 26460 5236 26516
rect 4844 26348 5012 26404
rect 4956 26292 5012 26348
rect 5068 26292 5124 26302
rect 4956 26236 5068 26292
rect 5068 26226 5124 26236
rect 4844 26178 4900 26190
rect 4844 26126 4846 26178
rect 4898 26126 4900 26178
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25566 4286 25618
rect 4338 25566 4340 25618
rect 4284 25172 4340 25566
rect 4620 25508 4676 25518
rect 4620 25414 4676 25452
rect 4284 25106 4340 25116
rect 4844 25060 4900 26126
rect 5068 25620 5124 25630
rect 5180 25620 5236 26460
rect 5292 26180 5348 26852
rect 5628 26292 5684 26302
rect 5516 26236 5628 26292
rect 5292 26178 5460 26180
rect 5292 26126 5294 26178
rect 5346 26126 5460 26178
rect 5292 26124 5460 26126
rect 5292 26114 5348 26124
rect 5068 25618 5236 25620
rect 5068 25566 5070 25618
rect 5122 25566 5236 25618
rect 5068 25564 5236 25566
rect 5068 25554 5124 25564
rect 5292 25508 5348 25518
rect 4844 24994 4900 25004
rect 5180 25172 5236 25182
rect 4732 24836 4788 24846
rect 4732 24742 4788 24780
rect 5180 24834 5236 25116
rect 5292 24946 5348 25452
rect 5292 24894 5294 24946
rect 5346 24894 5348 24946
rect 5292 24882 5348 24894
rect 5180 24782 5182 24834
rect 5234 24782 5236 24834
rect 5180 24770 5236 24782
rect 4844 24724 4900 24734
rect 4844 24722 5012 24724
rect 4844 24670 4846 24722
rect 4898 24670 5012 24722
rect 4844 24668 5012 24670
rect 4844 24658 4900 24668
rect 4732 24500 4788 24510
rect 4956 24500 5012 24668
rect 5292 24500 5348 24510
rect 4732 24498 4900 24500
rect 4732 24446 4734 24498
rect 4786 24446 4900 24498
rect 4732 24444 4900 24446
rect 4956 24498 5348 24500
rect 4956 24446 5294 24498
rect 5346 24446 5348 24498
rect 4956 24444 5348 24446
rect 4732 24434 4788 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4732 23156 4788 23166
rect 4844 23156 4900 24444
rect 5292 24434 5348 24444
rect 4732 23154 4900 23156
rect 4732 23102 4734 23154
rect 4786 23102 4900 23154
rect 4732 23100 4900 23102
rect 4732 23090 4788 23100
rect 4060 23042 4116 23054
rect 4060 22990 4062 23042
rect 4114 22990 4116 23042
rect 4060 20804 4116 22990
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5068 21588 5124 21598
rect 5068 21494 5124 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4060 20738 4116 20748
rect 3948 19954 4004 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5404 17444 5460 26124
rect 5516 21588 5572 26236
rect 5628 26198 5684 26236
rect 5852 25620 5908 25630
rect 5628 25508 5684 25518
rect 5628 25414 5684 25452
rect 5852 25506 5908 25564
rect 5852 25454 5854 25506
rect 5906 25454 5908 25506
rect 5852 25442 5908 25454
rect 5964 25508 6020 28588
rect 6748 27300 6804 31948
rect 6860 31892 6916 31902
rect 6860 31106 6916 31836
rect 6860 31054 6862 31106
rect 6914 31054 6916 31106
rect 6860 31042 6916 31054
rect 6748 27186 6804 27244
rect 6748 27134 6750 27186
rect 6802 27134 6804 27186
rect 6748 27122 6804 27134
rect 6188 26852 6244 26862
rect 6188 26850 6468 26852
rect 6188 26798 6190 26850
rect 6242 26798 6468 26850
rect 6188 26796 6468 26798
rect 6188 26786 6244 26796
rect 6412 26402 6468 26796
rect 6412 26350 6414 26402
rect 6466 26350 6468 26402
rect 6412 26338 6468 26350
rect 6748 25620 6804 25630
rect 6300 25508 6356 25518
rect 5964 25506 6692 25508
rect 5964 25454 6302 25506
rect 6354 25454 6692 25506
rect 5964 25452 6692 25454
rect 6300 25442 6356 25452
rect 5852 25284 5908 25294
rect 5852 24834 5908 25228
rect 5852 24782 5854 24834
rect 5906 24782 5908 24834
rect 5852 23380 5908 24782
rect 6076 25060 6132 25070
rect 6076 24722 6132 25004
rect 6076 24670 6078 24722
rect 6130 24670 6132 24722
rect 6076 24658 6132 24670
rect 6412 24836 6468 24846
rect 6412 23938 6468 24780
rect 6412 23886 6414 23938
rect 6466 23886 6468 23938
rect 6412 23874 6468 23886
rect 6636 23826 6692 25452
rect 6748 24834 6804 25564
rect 6860 25060 6916 25070
rect 6860 24946 6916 25004
rect 6860 24894 6862 24946
rect 6914 24894 6916 24946
rect 6860 24882 6916 24894
rect 6748 24782 6750 24834
rect 6802 24782 6804 24834
rect 6748 23938 6804 24782
rect 6748 23886 6750 23938
rect 6802 23886 6804 23938
rect 6748 23874 6804 23886
rect 6636 23774 6638 23826
rect 6690 23774 6692 23826
rect 6636 23762 6692 23774
rect 5852 23266 5908 23324
rect 5852 23214 5854 23266
rect 5906 23214 5908 23266
rect 5852 23202 5908 23214
rect 6412 23604 6468 23614
rect 6188 23044 6244 23054
rect 6188 22950 6244 22988
rect 5628 21588 5684 21598
rect 5516 21532 5628 21588
rect 5628 21522 5684 21532
rect 5740 21474 5796 21486
rect 5740 21422 5742 21474
rect 5794 21422 5796 21474
rect 5740 20690 5796 21422
rect 5964 20804 6020 20814
rect 5964 20710 6020 20748
rect 5740 20638 5742 20690
rect 5794 20638 5796 20690
rect 5740 20626 5796 20638
rect 6412 18116 6468 23548
rect 6860 23380 6916 23390
rect 6860 23286 6916 23324
rect 6972 21812 7028 33516
rect 7084 33346 7140 39340
rect 7644 39284 7700 39788
rect 7756 39508 7812 39788
rect 7756 39442 7812 39452
rect 7644 39228 7812 39284
rect 7196 38948 7252 38958
rect 7196 38854 7252 38892
rect 7308 38836 7364 38846
rect 7196 37156 7252 37166
rect 7308 37156 7364 38780
rect 7644 38500 7700 38510
rect 7644 37716 7700 38444
rect 7644 37650 7700 37660
rect 7644 37268 7700 37278
rect 7196 37154 7364 37156
rect 7196 37102 7198 37154
rect 7250 37102 7364 37154
rect 7196 37100 7364 37102
rect 7532 37156 7588 37166
rect 7196 37090 7252 37100
rect 7420 36258 7476 36270
rect 7420 36206 7422 36258
rect 7474 36206 7476 36258
rect 7420 35252 7476 36206
rect 7420 35186 7476 35196
rect 7532 35028 7588 37100
rect 7084 33294 7086 33346
rect 7138 33294 7140 33346
rect 7084 33282 7140 33294
rect 7196 34972 7588 35028
rect 7644 37154 7700 37212
rect 7644 37102 7646 37154
rect 7698 37102 7700 37154
rect 7644 35028 7700 37102
rect 7756 36482 7812 39228
rect 7868 38724 7924 44156
rect 8204 41188 8260 47068
rect 8316 46900 8372 46910
rect 8316 46806 8372 46844
rect 8316 45220 8372 45230
rect 8316 45106 8372 45164
rect 8316 45054 8318 45106
rect 8370 45054 8372 45106
rect 8316 44660 8372 45054
rect 8428 44996 8484 48412
rect 8540 48402 8596 48412
rect 8540 46002 8596 46014
rect 8540 45950 8542 46002
rect 8594 45950 8596 46002
rect 8540 45332 8596 45950
rect 8540 45266 8596 45276
rect 8652 44996 8708 51660
rect 8764 51380 8820 51390
rect 8764 51286 8820 51324
rect 8876 51154 8932 52108
rect 9100 52098 9156 52108
rect 8876 51102 8878 51154
rect 8930 51102 8932 51154
rect 8876 51090 8932 51102
rect 8876 50484 8932 50494
rect 9212 50428 9268 52222
rect 8764 50260 8820 50270
rect 8764 47012 8820 50204
rect 8764 46946 8820 46956
rect 8876 46786 8932 50428
rect 8988 50372 9268 50428
rect 8988 49028 9044 50372
rect 8988 48934 9044 48972
rect 9548 48692 9604 52780
rect 9660 51716 9716 55580
rect 9996 54628 10052 56252
rect 10108 55300 10164 55310
rect 10444 55300 10500 56254
rect 10892 56700 11060 56756
rect 10108 55298 10500 55300
rect 10108 55246 10110 55298
rect 10162 55246 10500 55298
rect 10108 55244 10500 55246
rect 10668 56082 10724 56094
rect 10668 56030 10670 56082
rect 10722 56030 10724 56082
rect 10108 55234 10164 55244
rect 10332 54628 10388 54638
rect 9996 54626 10388 54628
rect 9996 54574 10334 54626
rect 10386 54574 10388 54626
rect 9996 54572 10388 54574
rect 9772 53620 9828 53630
rect 9772 53170 9828 53564
rect 9772 53118 9774 53170
rect 9826 53118 9828 53170
rect 9772 53106 9828 53118
rect 10108 53058 10164 54572
rect 10332 54562 10388 54572
rect 10108 53006 10110 53058
rect 10162 53006 10164 53058
rect 10108 52994 10164 53006
rect 10220 54404 10276 54414
rect 9884 52948 9940 52958
rect 9884 52854 9940 52892
rect 10220 52162 10276 54348
rect 10668 53956 10724 56030
rect 10780 55188 10836 55198
rect 10780 55094 10836 55132
rect 10668 53900 10836 53956
rect 10556 53620 10612 53630
rect 10556 53526 10612 53564
rect 10556 53058 10612 53070
rect 10556 53006 10558 53058
rect 10610 53006 10612 53058
rect 10332 52948 10388 52958
rect 10332 52854 10388 52892
rect 10220 52110 10222 52162
rect 10274 52110 10276 52162
rect 10220 52098 10276 52110
rect 10556 52724 10612 53006
rect 10780 53060 10836 53900
rect 10780 52994 10836 53004
rect 9660 51650 9716 51660
rect 9772 51604 9828 51614
rect 9772 51510 9828 51548
rect 10332 51268 10388 51278
rect 10332 51174 10388 51212
rect 10556 51268 10612 52668
rect 10556 51202 10612 51212
rect 10668 52948 10724 52958
rect 9772 50596 9828 50606
rect 9772 50428 9828 50540
rect 10220 50484 10276 50522
rect 9772 50372 10052 50428
rect 10220 50418 10276 50428
rect 9436 48636 9604 48692
rect 9884 49026 9940 49038
rect 9884 48974 9886 49026
rect 9938 48974 9940 49026
rect 8988 48468 9044 48478
rect 8988 48374 9044 48412
rect 8876 46734 8878 46786
rect 8930 46734 8932 46786
rect 8876 45332 8932 46734
rect 8988 48244 9044 48254
rect 8988 46788 9044 48188
rect 9436 47572 9492 48636
rect 9548 48468 9604 48478
rect 9548 48374 9604 48412
rect 9884 48468 9940 48974
rect 9884 48402 9940 48412
rect 9996 48132 10052 50372
rect 8988 46722 9044 46732
rect 9100 47516 9492 47572
rect 9772 48130 10052 48132
rect 9772 48078 9998 48130
rect 10050 48078 10052 48130
rect 9772 48076 10052 48078
rect 8876 45266 8932 45276
rect 8876 45108 8932 45118
rect 8428 44940 8596 44996
rect 8316 44594 8372 44604
rect 8428 44772 8484 44782
rect 8428 41412 8484 44716
rect 8540 43428 8596 44940
rect 8652 44930 8708 44940
rect 8764 45052 8876 45108
rect 8540 43334 8596 43372
rect 8652 44660 8708 44670
rect 8652 42978 8708 44604
rect 8652 42926 8654 42978
rect 8706 42926 8708 42978
rect 8652 42914 8708 42926
rect 8764 42866 8820 45052
rect 8876 45042 8932 45052
rect 8988 44994 9044 45006
rect 8988 44942 8990 44994
rect 9042 44942 9044 44994
rect 8876 43650 8932 43662
rect 8876 43598 8878 43650
rect 8930 43598 8932 43650
rect 8876 42980 8932 43598
rect 8988 43652 9044 44942
rect 9100 44996 9156 47516
rect 9100 44930 9156 44940
rect 9212 47236 9268 47246
rect 8988 43586 9044 43596
rect 8876 42914 8932 42924
rect 9100 43540 9156 43550
rect 8764 42814 8766 42866
rect 8818 42814 8820 42866
rect 8764 42802 8820 42814
rect 9100 42642 9156 43484
rect 9100 42590 9102 42642
rect 9154 42590 9156 42642
rect 9100 42578 9156 42590
rect 8428 41346 8484 41356
rect 8540 41972 8596 41982
rect 8204 41132 8372 41188
rect 8092 41076 8148 41086
rect 7980 41074 8148 41076
rect 7980 41022 8094 41074
rect 8146 41022 8148 41074
rect 7980 41020 8148 41022
rect 7980 40292 8036 41020
rect 8092 41010 8148 41020
rect 8204 40962 8260 40974
rect 8204 40910 8206 40962
rect 8258 40910 8260 40962
rect 7980 40236 8148 40292
rect 8092 39620 8148 40236
rect 8092 39554 8148 39564
rect 7980 39508 8036 39518
rect 7980 39414 8036 39452
rect 8204 39508 8260 40910
rect 8092 39396 8148 39406
rect 8092 38948 8148 39340
rect 8092 38854 8148 38892
rect 7868 38658 7924 38668
rect 7980 38836 8036 38846
rect 7756 36430 7758 36482
rect 7810 36430 7812 36482
rect 7756 36418 7812 36430
rect 7868 37826 7924 37838
rect 7868 37774 7870 37826
rect 7922 37774 7924 37826
rect 7196 32788 7252 34972
rect 7532 34802 7588 34814
rect 7532 34750 7534 34802
rect 7586 34750 7588 34802
rect 7532 34692 7588 34750
rect 7084 32732 7252 32788
rect 7420 32900 7476 32910
rect 7084 31780 7140 32732
rect 7084 31714 7140 31724
rect 7196 32562 7252 32574
rect 7196 32510 7198 32562
rect 7250 32510 7252 32562
rect 7196 32452 7252 32510
rect 7196 31108 7252 32396
rect 7420 32450 7476 32844
rect 7420 32398 7422 32450
rect 7474 32398 7476 32450
rect 7420 32386 7476 32398
rect 7532 32228 7588 34636
rect 7644 32452 7700 34972
rect 7868 35700 7924 37774
rect 7980 36596 8036 38780
rect 8204 38668 8260 39452
rect 8316 40402 8372 41132
rect 8428 40964 8484 40974
rect 8428 40870 8484 40908
rect 8540 40628 8596 41916
rect 8988 41860 9044 41870
rect 8988 41766 9044 41804
rect 8428 40516 8484 40526
rect 8540 40516 8596 40572
rect 8428 40514 8596 40516
rect 8428 40462 8430 40514
rect 8482 40462 8596 40514
rect 8428 40460 8596 40462
rect 8428 40450 8484 40460
rect 8316 40350 8318 40402
rect 8370 40350 8372 40402
rect 8316 40292 8372 40350
rect 8316 38836 8372 40236
rect 8540 39396 8596 40460
rect 9212 39730 9268 47180
rect 9548 46788 9604 46798
rect 9436 46786 9604 46788
rect 9436 46734 9550 46786
rect 9602 46734 9604 46786
rect 9436 46732 9604 46734
rect 9212 39678 9214 39730
rect 9266 39678 9268 39730
rect 9212 39666 9268 39678
rect 9324 45780 9380 45790
rect 9324 45666 9380 45724
rect 9324 45614 9326 45666
rect 9378 45614 9380 45666
rect 9324 43652 9380 45614
rect 8988 39508 9044 39518
rect 9212 39508 9268 39518
rect 9044 39506 9268 39508
rect 9044 39454 9214 39506
rect 9266 39454 9268 39506
rect 9044 39452 9268 39454
rect 8988 39442 9044 39452
rect 9212 39442 9268 39452
rect 8540 39330 8596 39340
rect 8316 38770 8372 38780
rect 8988 38836 9044 38846
rect 8428 38722 8484 38734
rect 8428 38670 8430 38722
rect 8482 38670 8484 38722
rect 8428 38668 8484 38670
rect 8204 38612 8484 38668
rect 7980 36482 8036 36540
rect 7980 36430 7982 36482
rect 8034 36430 8036 36482
rect 7980 36418 8036 36430
rect 8092 38388 8148 38398
rect 8092 35924 8148 38332
rect 8204 38276 8260 38286
rect 8204 37268 8260 38220
rect 8428 38162 8484 38612
rect 8428 38110 8430 38162
rect 8482 38110 8484 38162
rect 8428 38098 8484 38110
rect 8876 38164 8932 38174
rect 8876 38050 8932 38108
rect 8876 37998 8878 38050
rect 8930 37998 8932 38050
rect 8876 37986 8932 37998
rect 8988 37492 9044 38780
rect 8988 37490 9156 37492
rect 8988 37438 8990 37490
rect 9042 37438 9156 37490
rect 8988 37436 9156 37438
rect 8988 37426 9044 37436
rect 8204 37202 8260 37212
rect 8316 37156 8372 37166
rect 8316 36482 8372 37100
rect 8316 36430 8318 36482
rect 8370 36430 8372 36482
rect 8316 36418 8372 36430
rect 8764 36596 8820 36606
rect 8204 36260 8260 36270
rect 8204 36258 8484 36260
rect 8204 36206 8206 36258
rect 8258 36206 8484 36258
rect 8204 36204 8484 36206
rect 8204 36194 8260 36204
rect 8092 35868 8372 35924
rect 8092 35700 8148 35710
rect 7868 35698 8148 35700
rect 7868 35646 8094 35698
rect 8146 35646 8148 35698
rect 7868 35644 8148 35646
rect 7756 34804 7812 34814
rect 7756 34710 7812 34748
rect 7756 32788 7812 32798
rect 7756 32562 7812 32732
rect 7756 32510 7758 32562
rect 7810 32510 7812 32562
rect 7756 32498 7812 32510
rect 7644 32386 7700 32396
rect 7532 32172 7700 32228
rect 7196 31042 7252 31052
rect 7308 31890 7364 31902
rect 7308 31838 7310 31890
rect 7362 31838 7364 31890
rect 7308 30996 7364 31838
rect 7532 31892 7588 31902
rect 7420 31778 7476 31790
rect 7420 31726 7422 31778
rect 7474 31726 7476 31778
rect 7420 31556 7476 31726
rect 7420 31490 7476 31500
rect 7308 30930 7364 30940
rect 7532 29652 7588 31836
rect 7532 29558 7588 29596
rect 7420 27300 7476 27310
rect 7420 25506 7476 27244
rect 7644 26908 7700 32172
rect 7756 31666 7812 31678
rect 7756 31614 7758 31666
rect 7810 31614 7812 31666
rect 7756 31108 7812 31614
rect 7756 31042 7812 31052
rect 7868 31106 7924 35644
rect 8092 35634 8148 35644
rect 7980 34690 8036 34702
rect 7980 34638 7982 34690
rect 8034 34638 8036 34690
rect 7980 34356 8036 34638
rect 7980 34290 8036 34300
rect 8092 34690 8148 34702
rect 8092 34638 8094 34690
rect 8146 34638 8148 34690
rect 7980 34018 8036 34030
rect 7980 33966 7982 34018
rect 8034 33966 8036 34018
rect 7980 32564 8036 33966
rect 8092 33348 8148 34638
rect 8092 33282 8148 33292
rect 8204 33236 8260 33246
rect 7980 32498 8036 32508
rect 8092 32788 8148 32798
rect 8092 32004 8148 32732
rect 8204 32674 8260 33180
rect 8204 32622 8206 32674
rect 8258 32622 8260 32674
rect 8204 32610 8260 32622
rect 7868 31054 7870 31106
rect 7922 31054 7924 31106
rect 7868 31042 7924 31054
rect 7980 31948 8148 32004
rect 7868 30884 7924 30894
rect 7756 30324 7812 30334
rect 7756 30098 7812 30268
rect 7756 30046 7758 30098
rect 7810 30046 7812 30098
rect 7756 30034 7812 30046
rect 7868 29652 7924 30828
rect 7980 30100 8036 31948
rect 8092 31780 8148 31790
rect 8092 31220 8148 31724
rect 8316 31220 8372 35868
rect 8428 35586 8484 36204
rect 8428 35534 8430 35586
rect 8482 35534 8484 35586
rect 8428 35522 8484 35534
rect 8652 35474 8708 35486
rect 8652 35422 8654 35474
rect 8706 35422 8708 35474
rect 8428 34914 8484 34926
rect 8428 34862 8430 34914
rect 8482 34862 8484 34914
rect 8428 33908 8484 34862
rect 8540 34356 8596 34366
rect 8540 34242 8596 34300
rect 8540 34190 8542 34242
rect 8594 34190 8596 34242
rect 8540 34178 8596 34190
rect 8428 33814 8484 33852
rect 8652 33460 8708 35422
rect 8652 33394 8708 33404
rect 8764 33236 8820 36540
rect 9100 36036 9156 37436
rect 9100 35980 9268 36036
rect 8876 35308 8932 35318
rect 9212 35308 9268 35980
rect 8876 35026 8932 35252
rect 8988 35196 9268 35308
rect 9212 35028 9268 35196
rect 8876 34974 8878 35026
rect 8930 34974 8932 35026
rect 8876 33906 8932 34974
rect 8876 33854 8878 33906
rect 8930 33854 8932 33906
rect 8876 33842 8932 33854
rect 8988 34972 9268 35028
rect 8764 33180 8932 33236
rect 8652 32900 8708 32910
rect 8652 32788 8708 32844
rect 8652 32786 8820 32788
rect 8652 32734 8654 32786
rect 8706 32734 8820 32786
rect 8652 32732 8820 32734
rect 8652 32722 8708 32732
rect 8092 31106 8148 31164
rect 8092 31054 8094 31106
rect 8146 31054 8148 31106
rect 8092 31042 8148 31054
rect 8204 31164 8372 31220
rect 8428 32676 8484 32686
rect 8092 30100 8148 30110
rect 7980 30098 8148 30100
rect 7980 30046 8094 30098
rect 8146 30046 8148 30098
rect 7980 30044 8148 30046
rect 8092 30034 8148 30044
rect 7980 29652 8036 29662
rect 7868 29650 8036 29652
rect 7868 29598 7982 29650
rect 8034 29598 8036 29650
rect 7868 29596 8036 29598
rect 7980 29586 8036 29596
rect 8204 27188 8260 31164
rect 8316 30996 8372 31006
rect 8316 30902 8372 30940
rect 8428 30994 8484 32620
rect 8428 30942 8430 30994
rect 8482 30942 8484 30994
rect 8428 30324 8484 30942
rect 8428 30258 8484 30268
rect 8540 32340 8596 32350
rect 8540 30210 8596 32284
rect 8652 31556 8708 31566
rect 8652 30884 8708 31500
rect 8652 30818 8708 30828
rect 8540 30158 8542 30210
rect 8594 30158 8596 30210
rect 8540 30146 8596 30158
rect 8764 29988 8820 32732
rect 8876 31556 8932 33180
rect 8876 31490 8932 31500
rect 8876 30770 8932 30782
rect 8876 30718 8878 30770
rect 8930 30718 8932 30770
rect 8876 30100 8932 30718
rect 8876 30034 8932 30044
rect 8652 29932 8820 29988
rect 8652 29652 8708 29932
rect 8988 29876 9044 34972
rect 9324 34916 9380 43596
rect 9436 43316 9492 46732
rect 9548 46722 9604 46732
rect 9548 45780 9604 45790
rect 9548 45686 9604 45724
rect 9772 45108 9828 48076
rect 9996 48066 10052 48076
rect 10332 50372 10388 50382
rect 9884 46900 9940 46910
rect 9884 46806 9940 46844
rect 10220 46676 10276 46686
rect 9996 46674 10276 46676
rect 9996 46622 10222 46674
rect 10274 46622 10276 46674
rect 9996 46620 10276 46622
rect 9996 45892 10052 46620
rect 10220 46610 10276 46620
rect 9884 45780 9940 45790
rect 9996 45780 10052 45836
rect 9884 45778 10052 45780
rect 9884 45726 9886 45778
rect 9938 45726 10052 45778
rect 9884 45724 10052 45726
rect 10220 45780 10276 45790
rect 9884 45714 9940 45724
rect 10220 45686 10276 45724
rect 9772 45042 9828 45052
rect 9660 44996 9716 45006
rect 9660 44884 9716 44940
rect 10108 44994 10164 45006
rect 10108 44942 10110 44994
rect 10162 44942 10164 44994
rect 9660 44828 9828 44884
rect 9436 42756 9492 43260
rect 9548 43540 9604 43550
rect 9772 43540 9828 44828
rect 10108 43764 10164 44942
rect 10108 43698 10164 43708
rect 10220 43652 10276 43662
rect 10332 43652 10388 50316
rect 10668 50372 10724 52892
rect 10892 52836 10948 56700
rect 11116 56644 11172 56654
rect 11004 56588 11116 56644
rect 11004 55636 11060 56588
rect 11116 56550 11172 56588
rect 11228 56420 11284 58828
rect 11452 58436 11508 62524
rect 11788 61572 11844 61582
rect 11788 61458 11844 61516
rect 11788 61406 11790 61458
rect 11842 61406 11844 61458
rect 11788 61394 11844 61406
rect 11564 61346 11620 61358
rect 11564 61294 11566 61346
rect 11618 61294 11620 61346
rect 11564 61236 11620 61294
rect 11564 61170 11620 61180
rect 12012 61348 12068 61358
rect 12012 60898 12068 61292
rect 12012 60846 12014 60898
rect 12066 60846 12068 60898
rect 12012 60834 12068 60846
rect 12124 61346 12180 61358
rect 12124 61294 12126 61346
rect 12178 61294 12180 61346
rect 12124 60564 12180 61294
rect 12124 60498 12180 60508
rect 11564 58996 11620 59006
rect 11620 58940 11732 58996
rect 11564 58930 11620 58940
rect 11004 55570 11060 55580
rect 11116 56364 11284 56420
rect 11340 58380 11508 58436
rect 10780 52780 10948 52836
rect 11004 53620 11060 53630
rect 10780 52500 10836 52780
rect 11004 52500 11060 53564
rect 11116 52724 11172 56364
rect 11228 53730 11284 53742
rect 11228 53678 11230 53730
rect 11282 53678 11284 53730
rect 11228 53060 11284 53678
rect 11228 52966 11284 53004
rect 11116 52668 11284 52724
rect 10780 52434 10836 52444
rect 10892 52444 11060 52500
rect 10892 51380 10948 52444
rect 11004 52276 11060 52286
rect 11004 52274 11172 52276
rect 11004 52222 11006 52274
rect 11058 52222 11172 52274
rect 11004 52220 11172 52222
rect 11004 52210 11060 52220
rect 11004 51380 11060 51390
rect 10892 51378 11060 51380
rect 10892 51326 11006 51378
rect 11058 51326 11060 51378
rect 10892 51324 11060 51326
rect 11004 51314 11060 51324
rect 10668 50306 10724 50316
rect 11116 50370 11172 52220
rect 11116 50318 11118 50370
rect 11170 50318 11172 50370
rect 11116 50306 11172 50318
rect 10444 50260 10500 50270
rect 10444 44436 10500 50204
rect 11004 49924 11060 49934
rect 10892 49868 11004 49924
rect 10556 49700 10612 49710
rect 10892 49700 10948 49868
rect 11004 49830 11060 49868
rect 11116 49812 11172 49850
rect 11116 49746 11172 49756
rect 10612 49644 10948 49700
rect 10556 49606 10612 49644
rect 11004 49588 11060 49598
rect 10892 49586 11060 49588
rect 10892 49534 11006 49586
rect 11058 49534 11060 49586
rect 10892 49532 11060 49534
rect 10556 49026 10612 49038
rect 10556 48974 10558 49026
rect 10610 48974 10612 49026
rect 10556 48916 10612 48974
rect 10556 48860 10836 48916
rect 10780 48466 10836 48860
rect 10780 48414 10782 48466
rect 10834 48414 10836 48466
rect 10780 48402 10836 48414
rect 10668 48244 10724 48254
rect 10892 48244 10948 49532
rect 11004 49522 11060 49532
rect 11116 49588 11172 49598
rect 11004 48356 11060 48366
rect 11116 48356 11172 49532
rect 11228 48804 11284 52668
rect 11340 50260 11396 58380
rect 11564 58324 11620 58334
rect 11452 58212 11508 58222
rect 11564 58212 11620 58268
rect 11452 58210 11620 58212
rect 11452 58158 11454 58210
rect 11506 58158 11620 58210
rect 11452 58156 11620 58158
rect 11452 58146 11508 58156
rect 11676 57764 11732 58940
rect 12236 58436 12292 64092
rect 12348 63812 12404 64428
rect 12572 63812 12628 63822
rect 12348 63810 12628 63812
rect 12348 63758 12574 63810
rect 12626 63758 12628 63810
rect 12348 63756 12628 63758
rect 12572 62132 12628 63756
rect 12572 62066 12628 62076
rect 12684 61572 12740 64652
rect 12908 64642 12964 64652
rect 12796 64482 12852 64494
rect 12796 64430 12798 64482
rect 12850 64430 12852 64482
rect 12796 64148 12852 64430
rect 13020 64372 13076 65772
rect 13020 64306 13076 64316
rect 13132 64260 13188 67004
rect 13468 65716 13524 67900
rect 14476 67620 14532 67630
rect 13916 67060 13972 67070
rect 14476 67060 14532 67564
rect 14588 67282 14644 70812
rect 14588 67230 14590 67282
rect 14642 67230 14644 67282
rect 14588 67218 14644 67230
rect 13916 67058 14644 67060
rect 13916 67006 13918 67058
rect 13970 67006 14478 67058
rect 14530 67006 14644 67058
rect 13916 67004 14644 67006
rect 13916 66994 13972 67004
rect 14476 66994 14532 67004
rect 14476 66836 14532 66846
rect 14140 66834 14532 66836
rect 14140 66782 14478 66834
rect 14530 66782 14532 66834
rect 14140 66780 14532 66782
rect 14140 66498 14196 66780
rect 14476 66770 14532 66780
rect 14588 66612 14644 67004
rect 14700 66836 14756 71036
rect 15372 70644 15428 70654
rect 15260 70084 15316 70094
rect 15372 70084 15428 70588
rect 16268 70196 16324 75518
rect 16828 74786 16884 76412
rect 17052 76402 17108 76412
rect 20076 76466 20132 76478
rect 20748 76468 20804 76478
rect 20076 76414 20078 76466
rect 20130 76414 20132 76466
rect 20076 76356 20132 76414
rect 20076 76290 20132 76300
rect 20300 76466 20804 76468
rect 20300 76414 20750 76466
rect 20802 76414 20804 76466
rect 20300 76412 20804 76414
rect 19068 75796 19124 75806
rect 20076 75796 20132 75806
rect 19124 75740 19236 75796
rect 19068 75702 19124 75740
rect 17052 75458 17108 75470
rect 17052 75406 17054 75458
rect 17106 75406 17108 75458
rect 17052 74900 17108 75406
rect 19068 75236 19124 75246
rect 17388 74900 17444 74910
rect 17052 74898 17444 74900
rect 17052 74846 17390 74898
rect 17442 74846 17444 74898
rect 17052 74844 17444 74846
rect 16828 74734 16830 74786
rect 16882 74734 16884 74786
rect 16828 74722 16884 74734
rect 16380 74114 16436 74126
rect 16380 74062 16382 74114
rect 16434 74062 16436 74114
rect 16380 74004 16436 74062
rect 16380 73938 16436 73948
rect 16828 74004 16884 74014
rect 16828 73910 16884 73948
rect 17388 74004 17444 74844
rect 18172 74788 18228 74798
rect 18172 74694 18228 74732
rect 18172 74228 18228 74238
rect 17388 73938 17444 73948
rect 17612 74114 17668 74126
rect 17612 74062 17614 74114
rect 17666 74062 17668 74114
rect 16604 73220 16660 73230
rect 16604 73126 16660 73164
rect 17164 73220 17220 73230
rect 17164 72658 17220 73164
rect 17612 73220 17668 74062
rect 18172 74114 18228 74172
rect 18172 74062 18174 74114
rect 18226 74062 18228 74114
rect 18172 74050 18228 74062
rect 18844 74002 18900 74014
rect 18844 73950 18846 74002
rect 18898 73950 18900 74002
rect 17612 73154 17668 73164
rect 17948 73332 18004 73342
rect 17948 73218 18004 73276
rect 18620 73332 18676 73342
rect 18620 73238 18676 73276
rect 17948 73166 17950 73218
rect 18002 73166 18004 73218
rect 17164 72606 17166 72658
rect 17218 72606 17220 72658
rect 17164 72594 17220 72606
rect 17052 72324 17108 72334
rect 17948 72324 18004 73166
rect 18844 72884 18900 73950
rect 19068 74004 19124 75180
rect 18844 72818 18900 72828
rect 18956 73332 19012 73342
rect 18172 72660 18228 72670
rect 18172 72566 18228 72604
rect 18956 72660 19012 73276
rect 18956 72566 19012 72604
rect 18732 72548 18788 72558
rect 17052 72322 17444 72324
rect 17052 72270 17054 72322
rect 17106 72270 17444 72322
rect 17052 72268 17444 72270
rect 17052 72258 17108 72268
rect 16604 71428 16660 71438
rect 16604 71090 16660 71372
rect 16604 71038 16606 71090
rect 16658 71038 16660 71090
rect 16604 71026 16660 71038
rect 16716 71316 16772 71326
rect 16268 70130 16324 70140
rect 15260 70082 15428 70084
rect 15260 70030 15262 70082
rect 15314 70030 15428 70082
rect 15260 70028 15428 70030
rect 15260 70018 15316 70028
rect 14924 69298 14980 69310
rect 14924 69246 14926 69298
rect 14978 69246 14980 69298
rect 14812 67060 14868 67070
rect 14812 66966 14868 67004
rect 14700 66780 14868 66836
rect 14140 66446 14142 66498
rect 14194 66446 14196 66498
rect 14140 66434 14196 66446
rect 14476 66556 14644 66612
rect 14476 66274 14532 66556
rect 14700 66500 14756 66510
rect 14476 66222 14478 66274
rect 14530 66222 14532 66274
rect 13804 66162 13860 66174
rect 13804 66110 13806 66162
rect 13858 66110 13860 66162
rect 13692 65716 13748 65726
rect 13468 65714 13748 65716
rect 13468 65662 13694 65714
rect 13746 65662 13748 65714
rect 13468 65660 13748 65662
rect 13692 65650 13748 65660
rect 13580 65492 13636 65502
rect 13468 65380 13524 65390
rect 13468 64372 13524 65324
rect 13580 64484 13636 65436
rect 13804 65380 13860 66110
rect 13916 66052 13972 66062
rect 13916 65602 13972 65996
rect 14028 66052 14084 66062
rect 14028 66050 14308 66052
rect 14028 65998 14030 66050
rect 14082 65998 14308 66050
rect 14028 65996 14308 65998
rect 14028 65986 14084 65996
rect 14252 65828 14308 65996
rect 14252 65762 14308 65772
rect 13916 65550 13918 65602
rect 13970 65550 13972 65602
rect 13916 65538 13972 65550
rect 14140 65604 14196 65614
rect 14140 65510 14196 65548
rect 14252 65492 14308 65502
rect 14476 65492 14532 66222
rect 14308 65436 14532 65492
rect 14588 66498 14756 66500
rect 14588 66446 14702 66498
rect 14754 66446 14756 66498
rect 14588 66444 14756 66446
rect 14252 65426 14308 65436
rect 13804 65324 13972 65380
rect 13692 65268 13748 65278
rect 13692 65266 13860 65268
rect 13692 65214 13694 65266
rect 13746 65214 13860 65266
rect 13692 65212 13860 65214
rect 13692 65202 13748 65212
rect 13692 64484 13748 64494
rect 13580 64482 13748 64484
rect 13580 64430 13694 64482
rect 13746 64430 13748 64482
rect 13580 64428 13748 64430
rect 13468 64316 13636 64372
rect 13132 64204 13412 64260
rect 13020 64148 13076 64158
rect 13132 64148 13188 64204
rect 12796 64146 13188 64148
rect 12796 64094 13022 64146
rect 13074 64094 13188 64146
rect 12796 64092 13188 64094
rect 13020 64082 13076 64092
rect 13244 64036 13300 64046
rect 13132 63252 13188 63262
rect 13132 62580 13188 63196
rect 12684 61478 12740 61516
rect 12796 62578 13188 62580
rect 12796 62526 13134 62578
rect 13186 62526 13188 62578
rect 12796 62524 13188 62526
rect 12796 61346 12852 62524
rect 13132 62514 13188 62524
rect 12796 61294 12798 61346
rect 12850 61294 12852 61346
rect 12796 61124 12852 61294
rect 12796 61058 12852 61068
rect 12908 62244 12964 62254
rect 13244 62188 13300 63980
rect 12236 58370 12292 58380
rect 12684 60004 12740 60014
rect 12348 58212 12404 58222
rect 11676 57698 11732 57708
rect 12236 58156 12348 58212
rect 11676 57538 11732 57550
rect 11676 57486 11678 57538
rect 11730 57486 11732 57538
rect 11676 57092 11732 57486
rect 11676 57036 12180 57092
rect 12124 56978 12180 57036
rect 12124 56926 12126 56978
rect 12178 56926 12180 56978
rect 12124 56914 12180 56926
rect 11452 56754 11508 56766
rect 11452 56702 11454 56754
rect 11506 56702 11508 56754
rect 11452 56082 11508 56702
rect 11788 56756 11844 56766
rect 12012 56756 12068 56766
rect 11788 56754 12068 56756
rect 11788 56702 11790 56754
rect 11842 56702 12014 56754
rect 12066 56702 12068 56754
rect 11788 56700 12068 56702
rect 11788 56690 11844 56700
rect 12012 56690 12068 56700
rect 12124 56756 12180 56766
rect 11564 56644 11620 56654
rect 11564 56550 11620 56588
rect 11564 56196 11620 56206
rect 11564 56102 11620 56140
rect 12124 56196 12180 56700
rect 12124 56102 12180 56140
rect 11452 56030 11454 56082
rect 11506 56030 11508 56082
rect 11452 54068 11508 56030
rect 11788 56082 11844 56094
rect 11788 56030 11790 56082
rect 11842 56030 11844 56082
rect 11788 54626 11844 56030
rect 12124 55524 12180 55534
rect 11900 55188 11956 55198
rect 11900 54738 11956 55132
rect 11900 54686 11902 54738
rect 11954 54686 11956 54738
rect 11900 54674 11956 54686
rect 11788 54574 11790 54626
rect 11842 54574 11844 54626
rect 11788 54562 11844 54574
rect 12124 54626 12180 55468
rect 12124 54574 12126 54626
rect 12178 54574 12180 54626
rect 12124 54562 12180 54574
rect 12236 54404 12292 58156
rect 12348 58146 12404 58156
rect 12572 57652 12628 57662
rect 12572 56868 12628 57596
rect 12460 56866 12628 56868
rect 12460 56814 12574 56866
rect 12626 56814 12628 56866
rect 12460 56812 12628 56814
rect 12348 56756 12404 56766
rect 12348 56662 12404 56700
rect 12348 54628 12404 54638
rect 12460 54628 12516 56812
rect 12572 56802 12628 56812
rect 12684 56644 12740 59948
rect 12908 57540 12964 62188
rect 13132 62132 13300 62188
rect 13020 61460 13076 61470
rect 13020 61366 13076 61404
rect 12684 56578 12740 56588
rect 12796 57484 12964 57540
rect 12348 54626 12740 54628
rect 12348 54574 12350 54626
rect 12402 54574 12740 54626
rect 12348 54572 12740 54574
rect 12348 54562 12404 54572
rect 12236 54348 12628 54404
rect 11452 54002 11508 54012
rect 11900 54068 11956 54078
rect 11564 53620 11620 53630
rect 11564 53170 11620 53564
rect 11564 53118 11566 53170
rect 11618 53118 11620 53170
rect 11564 53106 11620 53118
rect 11900 52948 11956 54012
rect 12012 53172 12068 53182
rect 12572 53172 12628 54348
rect 12012 53170 12628 53172
rect 12012 53118 12014 53170
rect 12066 53118 12574 53170
rect 12626 53118 12628 53170
rect 12012 53116 12628 53118
rect 12012 53106 12068 53116
rect 11900 52946 12180 52948
rect 11900 52894 11902 52946
rect 11954 52894 12180 52946
rect 11900 52892 12180 52894
rect 11900 52882 11956 52892
rect 11788 51940 11844 51950
rect 11788 51490 11844 51884
rect 11788 51438 11790 51490
rect 11842 51438 11844 51490
rect 11788 51426 11844 51438
rect 11340 50194 11396 50204
rect 11564 50148 11620 50158
rect 11228 48738 11284 48748
rect 11452 50036 11508 50046
rect 11004 48354 11172 48356
rect 11004 48302 11006 48354
rect 11058 48302 11172 48354
rect 11004 48300 11172 48302
rect 11004 48290 11060 48300
rect 11228 48244 11284 48254
rect 10668 48242 10948 48244
rect 10668 48190 10670 48242
rect 10722 48190 10948 48242
rect 10668 48188 10948 48190
rect 11116 48242 11396 48244
rect 11116 48190 11230 48242
rect 11282 48190 11396 48242
rect 11116 48188 11396 48190
rect 10668 48178 10724 48188
rect 10780 48020 10836 48030
rect 10556 47460 10612 47470
rect 10556 47366 10612 47404
rect 10668 46900 10724 46910
rect 10556 46786 10612 46798
rect 10556 46734 10558 46786
rect 10610 46734 10612 46786
rect 10556 46340 10612 46734
rect 10556 46274 10612 46284
rect 10556 45780 10612 45790
rect 10668 45780 10724 46844
rect 10556 45778 10724 45780
rect 10556 45726 10558 45778
rect 10610 45726 10724 45778
rect 10556 45724 10724 45726
rect 10556 45714 10612 45724
rect 10444 44370 10500 44380
rect 10780 43764 10836 47964
rect 11004 47458 11060 47470
rect 11004 47406 11006 47458
rect 11058 47406 11060 47458
rect 10892 47236 10948 47246
rect 11004 47236 11060 47406
rect 10948 47180 11060 47236
rect 10892 47170 10948 47180
rect 11116 46340 11172 48188
rect 11228 48178 11284 48188
rect 11340 48130 11396 48188
rect 11340 48078 11342 48130
rect 11394 48078 11396 48130
rect 11340 48066 11396 48078
rect 11228 46788 11284 46798
rect 11228 46450 11284 46732
rect 11228 46398 11230 46450
rect 11282 46398 11284 46450
rect 11228 46386 11284 46398
rect 11116 46274 11172 46284
rect 11452 46116 11508 49980
rect 11564 46900 11620 50092
rect 12124 49812 12180 52892
rect 12236 52946 12292 52958
rect 12236 52894 12238 52946
rect 12290 52894 12292 52946
rect 12236 52162 12292 52894
rect 12236 52110 12238 52162
rect 12290 52110 12292 52162
rect 12236 52098 12292 52110
rect 12348 51940 12404 51950
rect 12348 51846 12404 51884
rect 12236 50372 12292 50382
rect 12236 50034 12292 50316
rect 12236 49982 12238 50034
rect 12290 49982 12292 50034
rect 12236 49970 12292 49982
rect 12348 49924 12404 49934
rect 12348 49830 12404 49868
rect 12124 48468 12180 49756
rect 12236 49588 12292 49598
rect 12236 49494 12292 49532
rect 12236 48468 12292 48478
rect 12124 48466 12292 48468
rect 12124 48414 12238 48466
rect 12290 48414 12292 48466
rect 12124 48412 12292 48414
rect 12236 48402 12292 48412
rect 11676 48130 11732 48142
rect 11676 48078 11678 48130
rect 11730 48078 11732 48130
rect 11676 48018 11732 48078
rect 11676 47966 11678 48018
rect 11730 47966 11732 48018
rect 11676 47954 11732 47966
rect 11676 46900 11732 46910
rect 11620 46898 11732 46900
rect 11620 46846 11678 46898
rect 11730 46846 11732 46898
rect 11620 46844 11732 46846
rect 11564 46806 11620 46844
rect 11676 46834 11732 46844
rect 11004 46060 11508 46116
rect 11676 46564 11732 46574
rect 11676 46450 11732 46508
rect 11676 46398 11678 46450
rect 11730 46398 11732 46450
rect 11004 45778 11060 46060
rect 11564 46004 11620 46014
rect 11340 46002 11620 46004
rect 11340 45950 11566 46002
rect 11618 45950 11620 46002
rect 11340 45948 11620 45950
rect 11004 45726 11006 45778
rect 11058 45726 11060 45778
rect 11004 45556 11060 45726
rect 11228 45780 11284 45790
rect 11228 45686 11284 45724
rect 11004 45490 11060 45500
rect 11116 45666 11172 45678
rect 11116 45614 11118 45666
rect 11170 45614 11172 45666
rect 10892 44436 10948 44446
rect 10948 44380 11060 44436
rect 10892 44370 10948 44380
rect 10220 43650 10388 43652
rect 10220 43598 10222 43650
rect 10274 43598 10388 43650
rect 10220 43596 10388 43598
rect 10220 43586 10276 43596
rect 9884 43540 9940 43550
rect 9772 43538 10052 43540
rect 9772 43486 9886 43538
rect 9938 43486 10052 43538
rect 9772 43484 10052 43486
rect 9548 43204 9604 43484
rect 9884 43474 9940 43484
rect 9548 43138 9604 43148
rect 9660 43428 9716 43438
rect 9548 42756 9604 42766
rect 9436 42754 9604 42756
rect 9436 42702 9550 42754
rect 9602 42702 9604 42754
rect 9436 42700 9604 42702
rect 9548 42690 9604 42700
rect 9548 42530 9604 42542
rect 9548 42478 9550 42530
rect 9602 42478 9604 42530
rect 9548 40068 9604 42478
rect 9660 41970 9716 43372
rect 9884 43314 9940 43326
rect 9884 43262 9886 43314
rect 9938 43262 9940 43314
rect 9884 42978 9940 43262
rect 9884 42926 9886 42978
rect 9938 42926 9940 42978
rect 9884 42914 9940 42926
rect 9996 42420 10052 43484
rect 10332 42754 10388 43596
rect 10332 42702 10334 42754
rect 10386 42702 10388 42754
rect 10332 42690 10388 42702
rect 10444 43708 10836 43764
rect 10892 43762 10948 43774
rect 10892 43710 10894 43762
rect 10946 43710 10948 43762
rect 9996 42354 10052 42364
rect 10108 42642 10164 42654
rect 10108 42590 10110 42642
rect 10162 42590 10164 42642
rect 9660 41918 9662 41970
rect 9714 41918 9716 41970
rect 9660 41906 9716 41918
rect 9996 41860 10052 41870
rect 10108 41860 10164 42590
rect 10220 42532 10276 42542
rect 10220 42194 10276 42476
rect 10220 42142 10222 42194
rect 10274 42142 10276 42194
rect 10220 42130 10276 42142
rect 10052 41804 10164 41860
rect 9996 41794 10052 41804
rect 9772 40964 9828 40974
rect 9660 40628 9716 40638
rect 9660 40534 9716 40572
rect 9548 40012 9716 40068
rect 9548 38722 9604 38734
rect 9548 38670 9550 38722
rect 9602 38670 9604 38722
rect 9436 38164 9492 38174
rect 9436 37380 9492 38108
rect 9548 37492 9604 38670
rect 9660 38162 9716 40012
rect 9660 38110 9662 38162
rect 9714 38110 9716 38162
rect 9660 38098 9716 38110
rect 9548 37436 9716 37492
rect 9436 36484 9492 37324
rect 9548 37268 9604 37278
rect 9548 37174 9604 37212
rect 9660 36708 9716 37436
rect 9772 37266 9828 40908
rect 10108 40292 10164 40302
rect 10108 40198 10164 40236
rect 10444 37716 10500 43708
rect 10892 43652 10948 43710
rect 10780 43596 10948 43652
rect 11004 43652 11060 44380
rect 10556 43540 10612 43550
rect 10556 42532 10612 43484
rect 10556 42466 10612 42476
rect 10556 40068 10612 40078
rect 10556 39618 10612 40012
rect 10556 39566 10558 39618
rect 10610 39566 10612 39618
rect 10556 39554 10612 39566
rect 9772 37214 9774 37266
rect 9826 37214 9828 37266
rect 9772 37202 9828 37214
rect 10332 37660 10500 37716
rect 10108 37042 10164 37054
rect 10108 36990 10110 37042
rect 10162 36990 10164 37042
rect 9660 36652 9940 36708
rect 9660 36484 9716 36494
rect 9436 36482 9716 36484
rect 9436 36430 9662 36482
rect 9714 36430 9716 36482
rect 9436 36428 9716 36430
rect 9660 36418 9716 36428
rect 9548 36036 9604 36046
rect 9212 34860 9380 34916
rect 9436 35980 9548 36036
rect 9100 34356 9156 34366
rect 9100 34262 9156 34300
rect 9100 33906 9156 33918
rect 9100 33854 9102 33906
rect 9154 33854 9156 33906
rect 9100 31892 9156 33854
rect 9100 31826 9156 31836
rect 8988 29820 9156 29876
rect 8988 29652 9044 29662
rect 8652 29650 9044 29652
rect 8652 29598 8990 29650
rect 9042 29598 9044 29650
rect 8652 29596 9044 29598
rect 8988 29204 9044 29596
rect 8988 29138 9044 29148
rect 8540 28140 9044 28196
rect 8540 28082 8596 28140
rect 8540 28030 8542 28082
rect 8594 28030 8596 28082
rect 8540 28018 8596 28030
rect 8876 27972 8932 27982
rect 8764 27970 8932 27972
rect 8764 27918 8878 27970
rect 8930 27918 8932 27970
rect 8764 27916 8932 27918
rect 8652 27860 8708 27870
rect 7420 25454 7422 25506
rect 7474 25454 7476 25506
rect 7420 25284 7476 25454
rect 7420 25218 7476 25228
rect 7532 26852 7700 26908
rect 7756 26962 7812 26974
rect 7756 26910 7758 26962
rect 7810 26910 7812 26962
rect 7084 24724 7140 24734
rect 7308 24724 7364 24734
rect 7084 24722 7364 24724
rect 7084 24670 7086 24722
rect 7138 24670 7310 24722
rect 7362 24670 7364 24722
rect 7084 24668 7364 24670
rect 7084 24658 7140 24668
rect 7308 24658 7364 24668
rect 7084 22372 7140 22382
rect 7420 22372 7476 22382
rect 7532 22372 7588 26852
rect 7756 25620 7812 26910
rect 8204 26962 8260 27132
rect 8428 27858 8708 27860
rect 8428 27806 8654 27858
rect 8706 27806 8708 27858
rect 8428 27804 8708 27806
rect 8428 27074 8484 27804
rect 8652 27794 8708 27804
rect 8764 27076 8820 27916
rect 8876 27906 8932 27916
rect 8988 27972 9044 28140
rect 9100 27972 9156 29820
rect 8988 27970 9156 27972
rect 8988 27918 8990 27970
rect 9042 27918 9156 27970
rect 8988 27916 9156 27918
rect 8988 27906 9044 27916
rect 8876 27188 8932 27198
rect 9212 27188 9268 34860
rect 9324 34692 9380 34702
rect 9436 34692 9492 35980
rect 9548 35970 9604 35980
rect 9324 34690 9492 34692
rect 9324 34638 9326 34690
rect 9378 34638 9492 34690
rect 9324 34636 9492 34638
rect 9772 34690 9828 34702
rect 9772 34638 9774 34690
rect 9826 34638 9828 34690
rect 9324 34356 9380 34636
rect 9772 34580 9828 34638
rect 9772 34514 9828 34524
rect 9324 34290 9380 34300
rect 9884 33460 9940 36652
rect 9772 33404 9940 33460
rect 9548 33348 9604 33386
rect 9604 33292 9716 33348
rect 9548 33282 9604 33292
rect 9324 33236 9380 33246
rect 9324 33142 9380 33180
rect 9548 33124 9604 33134
rect 9548 33030 9604 33068
rect 9548 32676 9604 32686
rect 9324 32620 9548 32676
rect 9324 31778 9380 32620
rect 9548 32582 9604 32620
rect 9660 32564 9716 33292
rect 9660 32498 9716 32508
rect 9772 31892 9828 33404
rect 9884 33234 9940 33246
rect 9884 33182 9886 33234
rect 9938 33182 9940 33234
rect 9884 32786 9940 33182
rect 9884 32734 9886 32786
rect 9938 32734 9940 32786
rect 9884 32722 9940 32734
rect 9996 33236 10052 33246
rect 9996 32004 10052 33180
rect 9996 31938 10052 31948
rect 10108 32788 10164 36990
rect 10332 33572 10388 37660
rect 10780 37492 10836 43596
rect 11004 43540 11060 43596
rect 10892 43538 11060 43540
rect 10892 43486 11006 43538
rect 11058 43486 11060 43538
rect 10892 43484 11060 43486
rect 10892 42756 10948 43484
rect 11004 43474 11060 43484
rect 11004 42980 11060 42990
rect 11116 42980 11172 45614
rect 11228 43540 11284 43550
rect 11340 43540 11396 45948
rect 11564 45938 11620 45948
rect 11676 45778 11732 46398
rect 12460 45892 12516 53116
rect 12572 53106 12628 53116
rect 12572 52164 12628 52174
rect 12572 52070 12628 52108
rect 12684 52162 12740 54572
rect 12796 52836 12852 57484
rect 12908 55410 12964 55422
rect 12908 55358 12910 55410
rect 12962 55358 12964 55410
rect 12908 54964 12964 55358
rect 12908 54898 12964 54908
rect 13020 54740 13076 54750
rect 13132 54740 13188 62132
rect 13356 59668 13412 64204
rect 13468 63924 13524 63934
rect 13468 63830 13524 63868
rect 13580 62188 13636 64316
rect 13692 63588 13748 64428
rect 13804 63810 13860 65212
rect 13916 64930 13972 65324
rect 14588 65268 14644 66444
rect 14700 66434 14756 66444
rect 14812 65714 14868 66780
rect 14924 66050 14980 69246
rect 15260 67620 15316 67630
rect 15260 67526 15316 67564
rect 15036 67060 15092 67070
rect 15036 67058 15316 67060
rect 15036 67006 15038 67058
rect 15090 67006 15316 67058
rect 15036 67004 15316 67006
rect 15036 66994 15092 67004
rect 15036 66276 15092 66286
rect 15036 66182 15092 66220
rect 15260 66274 15316 67004
rect 15372 66948 15428 70028
rect 15484 66948 15540 66958
rect 15372 66946 15540 66948
rect 15372 66894 15486 66946
rect 15538 66894 15540 66946
rect 15372 66892 15540 66894
rect 15484 66836 15540 66892
rect 15932 66948 15988 66958
rect 15932 66854 15988 66892
rect 15484 66780 15764 66836
rect 15260 66222 15262 66274
rect 15314 66222 15316 66274
rect 14924 65998 14926 66050
rect 14978 65998 14980 66050
rect 14924 65986 14980 65998
rect 14812 65662 14814 65714
rect 14866 65662 14868 65714
rect 14812 65650 14868 65662
rect 14924 65828 14980 65838
rect 13916 64878 13918 64930
rect 13970 64878 13972 64930
rect 13916 64596 13972 64878
rect 14252 65212 14644 65268
rect 14700 65492 14756 65502
rect 14252 64930 14308 65212
rect 14252 64878 14254 64930
rect 14306 64878 14308 64930
rect 14252 64866 14308 64878
rect 14252 64706 14308 64718
rect 14252 64654 14254 64706
rect 14306 64654 14308 64706
rect 13972 64540 14084 64596
rect 13916 64530 13972 64540
rect 13916 64034 13972 64046
rect 13916 63982 13918 64034
rect 13970 63982 13972 64034
rect 13916 63924 13972 63982
rect 14028 64036 14084 64540
rect 14140 64036 14196 64046
rect 14028 64034 14196 64036
rect 14028 63982 14142 64034
rect 14194 63982 14196 64034
rect 14028 63980 14196 63982
rect 14140 63970 14196 63980
rect 14252 64036 14308 64654
rect 14588 64596 14644 64606
rect 14588 64502 14644 64540
rect 14588 64036 14644 64046
rect 14308 64034 14644 64036
rect 14308 63982 14590 64034
rect 14642 63982 14644 64034
rect 14308 63980 14644 63982
rect 14252 63970 14308 63980
rect 14588 63970 14644 63980
rect 13916 63858 13972 63868
rect 13804 63758 13806 63810
rect 13858 63758 13860 63810
rect 13804 63746 13860 63758
rect 13692 63532 14420 63588
rect 14028 63028 14084 63038
rect 14252 63028 14308 63038
rect 14028 63026 14308 63028
rect 14028 62974 14030 63026
rect 14082 62974 14254 63026
rect 14306 62974 14308 63026
rect 14028 62972 14308 62974
rect 14028 62580 14084 62972
rect 14252 62962 14308 62972
rect 14028 62514 14084 62524
rect 14252 62242 14308 62254
rect 14252 62190 14254 62242
rect 14306 62190 14308 62242
rect 14252 62188 14308 62190
rect 13580 62132 13972 62188
rect 13692 61570 13748 61582
rect 13692 61518 13694 61570
rect 13746 61518 13748 61570
rect 13468 61458 13524 61470
rect 13468 61406 13470 61458
rect 13522 61406 13524 61458
rect 13468 61236 13524 61406
rect 13692 61460 13748 61518
rect 13692 61394 13748 61404
rect 13580 61348 13636 61358
rect 13580 61254 13636 61292
rect 13804 61348 13860 61358
rect 13468 61170 13524 61180
rect 13356 59602 13412 59612
rect 13468 58434 13524 58446
rect 13468 58382 13470 58434
rect 13522 58382 13524 58434
rect 13356 56756 13412 56766
rect 13356 56662 13412 56700
rect 13468 56532 13524 58382
rect 13804 58212 13860 61292
rect 13804 58146 13860 58156
rect 13804 57764 13860 57774
rect 13804 57540 13860 57708
rect 13580 57538 13860 57540
rect 13580 57486 13806 57538
rect 13858 57486 13860 57538
rect 13580 57484 13860 57486
rect 13580 56754 13636 57484
rect 13804 57474 13860 57484
rect 13580 56702 13582 56754
rect 13634 56702 13636 56754
rect 13580 56690 13636 56702
rect 13692 56754 13748 56766
rect 13692 56702 13694 56754
rect 13746 56702 13748 56754
rect 13356 56476 13524 56532
rect 13356 55972 13412 56476
rect 13468 56196 13524 56206
rect 13468 56102 13524 56140
rect 13356 55906 13412 55916
rect 13580 55524 13636 55534
rect 13580 55430 13636 55468
rect 13692 55300 13748 56702
rect 13916 56196 13972 62132
rect 14028 62132 14308 62188
rect 14364 62188 14420 63532
rect 14588 63028 14644 63038
rect 14700 63028 14756 65436
rect 14812 65268 14868 65278
rect 14812 65174 14868 65212
rect 14924 65044 14980 65772
rect 14812 64988 14980 65044
rect 15036 65716 15092 65726
rect 15036 65490 15092 65660
rect 15260 65716 15316 66222
rect 15708 66162 15764 66780
rect 16268 66276 16324 66286
rect 16268 66274 16660 66276
rect 16268 66222 16270 66274
rect 16322 66222 16660 66274
rect 16268 66220 16660 66222
rect 16268 66210 16324 66220
rect 15708 66110 15710 66162
rect 15762 66110 15764 66162
rect 15596 66052 15652 66062
rect 15596 65958 15652 65996
rect 15596 65716 15652 65726
rect 15260 65714 15652 65716
rect 15260 65662 15598 65714
rect 15650 65662 15652 65714
rect 15260 65660 15652 65662
rect 15260 65604 15316 65660
rect 15596 65650 15652 65660
rect 15260 65510 15316 65548
rect 15036 65438 15038 65490
rect 15090 65438 15092 65490
rect 14812 64484 14868 64988
rect 15036 64932 15092 65438
rect 15596 65492 15652 65502
rect 15596 65156 15652 65436
rect 15596 65090 15652 65100
rect 15036 64876 15316 64932
rect 14924 64708 14980 64718
rect 15148 64708 15204 64718
rect 14924 64706 15148 64708
rect 14924 64654 14926 64706
rect 14978 64654 15148 64706
rect 14924 64652 15148 64654
rect 14924 64642 14980 64652
rect 15148 64642 15204 64652
rect 15260 64484 15316 64876
rect 15484 64484 15540 64494
rect 14812 64428 15092 64484
rect 15260 64428 15484 64484
rect 14588 63026 14756 63028
rect 14588 62974 14590 63026
rect 14642 62974 14756 63026
rect 14588 62972 14756 62974
rect 14924 63588 14980 63598
rect 14588 62962 14644 62972
rect 14700 62580 14756 62590
rect 14700 62486 14756 62524
rect 14924 62356 14980 63532
rect 14924 62290 14980 62300
rect 14364 62132 14532 62188
rect 14028 61458 14084 62132
rect 14028 61406 14030 61458
rect 14082 61406 14084 61458
rect 14028 60900 14084 61406
rect 14364 61572 14420 61582
rect 14364 61458 14420 61516
rect 14364 61406 14366 61458
rect 14418 61406 14420 61458
rect 14364 61394 14420 61406
rect 14028 60834 14084 60844
rect 14140 61124 14196 61134
rect 14140 60674 14196 61068
rect 14140 60622 14142 60674
rect 14194 60622 14196 60674
rect 14140 60610 14196 60622
rect 14252 58322 14308 58334
rect 14252 58270 14254 58322
rect 14306 58270 14308 58322
rect 14252 57876 14308 58270
rect 14364 57876 14420 57886
rect 14252 57874 14420 57876
rect 14252 57822 14366 57874
rect 14418 57822 14420 57874
rect 14252 57820 14420 57822
rect 14364 57810 14420 57820
rect 14140 57650 14196 57662
rect 14140 57598 14142 57650
rect 14194 57598 14196 57650
rect 14140 56306 14196 57598
rect 14140 56254 14142 56306
rect 14194 56254 14196 56306
rect 14140 56242 14196 56254
rect 13972 56140 14084 56196
rect 13916 56102 13972 56140
rect 13804 56084 13860 56094
rect 13804 55990 13860 56028
rect 13916 55972 13972 55982
rect 13692 55298 13860 55300
rect 13692 55246 13694 55298
rect 13746 55246 13860 55298
rect 13692 55244 13860 55246
rect 13692 55234 13748 55244
rect 13580 55074 13636 55086
rect 13580 55022 13582 55074
rect 13634 55022 13636 55074
rect 13580 54964 13636 55022
rect 13580 54898 13636 54908
rect 13468 54740 13524 54750
rect 13020 54738 13524 54740
rect 13020 54686 13022 54738
rect 13074 54686 13470 54738
rect 13522 54686 13524 54738
rect 13020 54684 13524 54686
rect 12908 52836 12964 52846
rect 12796 52780 12908 52836
rect 12908 52770 12964 52780
rect 12684 52110 12686 52162
rect 12738 52110 12740 52162
rect 12684 51044 12740 52110
rect 12684 50978 12740 50988
rect 13020 50428 13076 54684
rect 13468 54674 13524 54684
rect 13580 54628 13636 54638
rect 13580 54534 13636 54572
rect 13244 54514 13300 54526
rect 13244 54462 13246 54514
rect 13298 54462 13300 54514
rect 12684 50372 12740 50382
rect 12684 49138 12740 50316
rect 12684 49086 12686 49138
rect 12738 49086 12740 49138
rect 12684 49074 12740 49086
rect 12796 50372 13076 50428
rect 13132 53844 13188 53854
rect 12572 48356 12628 48366
rect 12572 48262 12628 48300
rect 12124 45836 12516 45892
rect 12572 46116 12628 46126
rect 11676 45726 11678 45778
rect 11730 45726 11732 45778
rect 11676 45714 11732 45726
rect 11900 45780 11956 45790
rect 11900 45686 11956 45724
rect 11452 43652 11844 43708
rect 11452 43650 11508 43652
rect 11452 43598 11454 43650
rect 11506 43598 11508 43650
rect 11452 43586 11508 43598
rect 11228 43538 11396 43540
rect 11228 43486 11230 43538
rect 11282 43486 11396 43538
rect 11228 43484 11396 43486
rect 11676 43540 11732 43550
rect 11228 43474 11284 43484
rect 11004 42978 11172 42980
rect 11004 42926 11006 42978
rect 11058 42926 11172 42978
rect 11004 42924 11172 42926
rect 11004 42914 11060 42924
rect 11228 42868 11284 42878
rect 10892 42754 11060 42756
rect 10892 42702 10894 42754
rect 10946 42702 11060 42754
rect 10892 42700 11060 42702
rect 10892 42690 10948 42700
rect 10892 42532 10948 42542
rect 10892 42194 10948 42476
rect 10892 42142 10894 42194
rect 10946 42142 10948 42194
rect 10892 42130 10948 42142
rect 11004 41746 11060 42700
rect 11004 41694 11006 41746
rect 11058 41694 11060 41746
rect 11004 41682 11060 41694
rect 11228 42754 11284 42812
rect 11228 42702 11230 42754
rect 11282 42702 11284 42754
rect 11228 40628 11284 42702
rect 11452 42756 11508 42766
rect 11676 42756 11732 43484
rect 11452 42754 11732 42756
rect 11452 42702 11454 42754
rect 11506 42702 11732 42754
rect 11452 42700 11732 42702
rect 11452 42690 11508 42700
rect 11340 42530 11396 42542
rect 11788 42532 11844 43652
rect 12012 43652 12068 43662
rect 12012 43538 12068 43596
rect 12012 43486 12014 43538
rect 12066 43486 12068 43538
rect 12012 43474 12068 43486
rect 12124 43316 12180 45836
rect 12236 45668 12292 45678
rect 12236 45218 12292 45612
rect 12348 45668 12404 45678
rect 12572 45668 12628 46060
rect 12348 45666 12628 45668
rect 12348 45614 12350 45666
rect 12402 45614 12628 45666
rect 12348 45612 12628 45614
rect 12348 45556 12404 45612
rect 12348 45490 12404 45500
rect 12236 45166 12238 45218
rect 12290 45166 12292 45218
rect 12236 45154 12292 45166
rect 12796 45108 12852 50372
rect 12348 45052 12852 45108
rect 13020 48468 13076 48478
rect 13020 47796 13076 48412
rect 13020 45106 13076 47740
rect 13020 45054 13022 45106
rect 13074 45054 13076 45106
rect 12348 44996 12404 45052
rect 13020 45042 13076 45054
rect 12012 43260 12180 43316
rect 12236 44940 12404 44996
rect 11900 42532 11956 42542
rect 11340 42478 11342 42530
rect 11394 42478 11396 42530
rect 11340 42084 11396 42478
rect 11676 42530 11956 42532
rect 11676 42478 11902 42530
rect 11954 42478 11956 42530
rect 11676 42476 11956 42478
rect 11340 42028 11620 42084
rect 11340 41858 11396 41870
rect 11340 41806 11342 41858
rect 11394 41806 11396 41858
rect 11340 41746 11396 41806
rect 11340 41694 11342 41746
rect 11394 41694 11396 41746
rect 11340 41682 11396 41694
rect 11228 40572 11396 40628
rect 11228 40402 11284 40414
rect 11228 40350 11230 40402
rect 11282 40350 11284 40402
rect 11228 39732 11284 40350
rect 11116 39396 11172 39406
rect 11116 39302 11172 39340
rect 10444 37436 10836 37492
rect 10444 36594 10500 37436
rect 10444 36542 10446 36594
rect 10498 36542 10500 36594
rect 10444 36530 10500 36542
rect 11228 35588 11284 39676
rect 10332 33506 10388 33516
rect 11116 35586 11284 35588
rect 11116 35534 11230 35586
rect 11282 35534 11284 35586
rect 11116 35532 11284 35534
rect 10332 33236 10388 33246
rect 10332 33142 10388 33180
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 9324 31714 9380 31726
rect 9436 31836 9828 31892
rect 9436 28756 9492 31836
rect 9548 31668 9604 31678
rect 9548 31574 9604 31612
rect 9996 31556 10052 31566
rect 9884 31500 9996 31556
rect 9660 31220 9716 31230
rect 9548 30996 9604 31006
rect 9548 29426 9604 30940
rect 9660 30994 9716 31164
rect 9660 30942 9662 30994
rect 9714 30942 9716 30994
rect 9660 30930 9716 30942
rect 9884 30996 9940 31500
rect 9996 31462 10052 31500
rect 10108 31332 10164 32732
rect 10220 33124 10276 33134
rect 10220 32340 10276 33068
rect 10444 33124 10500 33134
rect 10668 33124 10724 33134
rect 10444 33122 10612 33124
rect 10444 33070 10446 33122
rect 10498 33070 10612 33122
rect 10444 33068 10612 33070
rect 10444 33058 10500 33068
rect 10556 32788 10612 33068
rect 10668 33030 10724 33068
rect 10556 32732 11060 32788
rect 11004 32676 11060 32732
rect 11004 32582 11060 32620
rect 10220 32274 10276 32284
rect 10668 32564 10724 32574
rect 10668 31778 10724 32508
rect 11116 32452 11172 35532
rect 11228 35522 11284 35532
rect 11004 32396 11172 32452
rect 10668 31726 10670 31778
rect 10722 31726 10724 31778
rect 10668 31714 10724 31726
rect 10892 32004 10948 32014
rect 10892 31778 10948 31948
rect 10892 31726 10894 31778
rect 10946 31726 10948 31778
rect 10892 31714 10948 31726
rect 9884 30902 9940 30940
rect 9996 31276 10164 31332
rect 9548 29374 9550 29426
rect 9602 29374 9604 29426
rect 9548 29362 9604 29374
rect 9660 29986 9716 29998
rect 9660 29934 9662 29986
rect 9714 29934 9716 29986
rect 9436 28644 9492 28700
rect 9548 28644 9604 28654
rect 9436 28642 9604 28644
rect 9436 28590 9550 28642
rect 9602 28590 9604 28642
rect 9436 28588 9604 28590
rect 9548 28578 9604 28588
rect 8876 27094 8932 27132
rect 8988 27132 9268 27188
rect 8428 27022 8430 27074
rect 8482 27022 8484 27074
rect 8428 27010 8484 27022
rect 8652 27020 8820 27076
rect 8204 26910 8206 26962
rect 8258 26910 8260 26962
rect 8204 26898 8260 26910
rect 8652 26908 8708 27020
rect 8988 26908 9044 27132
rect 9660 26908 9716 29934
rect 9772 29428 9828 29438
rect 9996 29428 10052 31276
rect 10108 31108 10164 31118
rect 10108 30210 10164 31052
rect 10892 31106 10948 31118
rect 10892 31054 10894 31106
rect 10946 31054 10948 31106
rect 10108 30158 10110 30210
rect 10162 30158 10164 30210
rect 10108 30146 10164 30158
rect 10556 30882 10612 30894
rect 10556 30830 10558 30882
rect 10610 30830 10612 30882
rect 10556 29652 10612 30830
rect 10556 29586 10612 29596
rect 10780 30884 10836 30894
rect 9772 29426 10052 29428
rect 9772 29374 9774 29426
rect 9826 29374 10052 29426
rect 9772 29372 10052 29374
rect 10444 29428 10500 29438
rect 10668 29428 10724 29438
rect 10444 29426 10724 29428
rect 10444 29374 10446 29426
rect 10498 29374 10670 29426
rect 10722 29374 10724 29426
rect 10444 29372 10724 29374
rect 9772 29362 9828 29372
rect 10444 29362 10500 29372
rect 10668 29362 10724 29372
rect 9772 29204 9828 29214
rect 9996 29204 10052 29214
rect 9828 29202 10052 29204
rect 9828 29150 9998 29202
rect 10050 29150 10052 29202
rect 9828 29148 10052 29150
rect 9772 29138 9828 29148
rect 9996 29138 10052 29148
rect 10780 28866 10836 30828
rect 10892 29426 10948 31054
rect 10892 29374 10894 29426
rect 10946 29374 10948 29426
rect 10892 29362 10948 29374
rect 10780 28814 10782 28866
rect 10834 28814 10836 28866
rect 10780 28802 10836 28814
rect 10780 28644 10836 28654
rect 9884 28532 9940 28542
rect 8540 26852 8708 26908
rect 8764 26852 9044 26908
rect 9100 26852 9716 26908
rect 9772 28418 9828 28430
rect 9772 28366 9774 28418
rect 9826 28366 9828 28418
rect 8540 26178 8596 26852
rect 8540 26126 8542 26178
rect 8594 26126 8596 26178
rect 8540 26114 8596 26126
rect 7756 25526 7812 25564
rect 8092 25508 8148 25518
rect 8540 25508 8596 25518
rect 8092 25506 8596 25508
rect 8092 25454 8094 25506
rect 8146 25454 8542 25506
rect 8594 25454 8596 25506
rect 8092 25452 8596 25454
rect 8092 25442 8148 25452
rect 8204 24610 8260 25452
rect 8540 25442 8596 25452
rect 8316 25284 8372 25294
rect 8316 24722 8372 25228
rect 8316 24670 8318 24722
rect 8370 24670 8372 24722
rect 8316 24658 8372 24670
rect 8204 24558 8206 24610
rect 8258 24558 8260 24610
rect 8204 24546 8260 24558
rect 8316 24498 8372 24510
rect 8316 24446 8318 24498
rect 8370 24446 8372 24498
rect 7084 22370 7588 22372
rect 7084 22318 7086 22370
rect 7138 22318 7422 22370
rect 7474 22318 7588 22370
rect 7084 22316 7588 22318
rect 7644 23044 7700 23054
rect 7644 22484 7700 22988
rect 7644 22372 7700 22428
rect 7756 22372 7812 22382
rect 7644 22370 7812 22372
rect 7644 22318 7758 22370
rect 7810 22318 7812 22370
rect 7644 22316 7812 22318
rect 8316 22372 8372 24446
rect 8540 22484 8596 22494
rect 8540 22390 8596 22428
rect 8428 22372 8484 22382
rect 8316 22316 8428 22372
rect 7084 22306 7140 22316
rect 7420 22306 7476 22316
rect 7756 22306 7812 22316
rect 8428 22278 8484 22316
rect 7532 22148 7588 22158
rect 7532 22146 7700 22148
rect 7532 22094 7534 22146
rect 7586 22094 7700 22146
rect 7532 22092 7700 22094
rect 7532 22082 7588 22092
rect 6972 21746 7028 21756
rect 7644 21476 7700 22092
rect 8316 21588 8372 21598
rect 8316 21494 8372 21532
rect 7868 21476 7924 21486
rect 7644 21474 7924 21476
rect 7644 21422 7870 21474
rect 7922 21422 7924 21474
rect 7644 21420 7924 21422
rect 7868 21410 7924 21420
rect 6412 18050 6468 18060
rect 5516 17444 5572 17454
rect 5404 17388 5516 17444
rect 5516 17378 5572 17388
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 3276 3390 3278 3442
rect 3330 3390 3332 3442
rect 3276 3378 3332 3390
rect 6748 3444 6804 3454
rect 6972 3444 7028 3454
rect 6748 3442 7028 3444
rect 6748 3390 6750 3442
rect 6802 3390 6974 3442
rect 7026 3390 7028 3442
rect 6748 3388 7028 3390
rect 6748 800 6804 3388
rect 6972 3378 7028 3388
rect 7308 3444 7364 3454
rect 7308 3350 7364 3388
rect 8764 3444 8820 26852
rect 8988 26292 9044 26302
rect 8988 26198 9044 26236
rect 9100 25506 9156 26852
rect 9772 26180 9828 28366
rect 9884 27858 9940 28476
rect 10108 28530 10164 28542
rect 10108 28478 10110 28530
rect 10162 28478 10164 28530
rect 10108 28308 10164 28478
rect 10668 28532 10724 28542
rect 10668 28438 10724 28476
rect 10780 28532 10836 28588
rect 10780 28530 10948 28532
rect 10780 28478 10782 28530
rect 10834 28478 10948 28530
rect 10780 28476 10948 28478
rect 10780 28466 10836 28476
rect 10108 28252 10388 28308
rect 9884 27806 9886 27858
rect 9938 27806 9940 27858
rect 9884 27794 9940 27806
rect 10108 27970 10164 27982
rect 10108 27918 10110 27970
rect 10162 27918 10164 27970
rect 10108 27860 10164 27918
rect 10332 27860 10388 28252
rect 10780 28196 10836 28206
rect 10444 27860 10500 27870
rect 10332 27858 10500 27860
rect 10332 27806 10446 27858
rect 10498 27806 10500 27858
rect 10332 27804 10500 27806
rect 10108 27794 10164 27804
rect 10332 26964 10388 26974
rect 10444 26964 10500 27804
rect 10668 26964 10724 26974
rect 10332 26962 10724 26964
rect 10332 26910 10334 26962
rect 10386 26910 10670 26962
rect 10722 26910 10724 26962
rect 10332 26908 10724 26910
rect 9996 26852 10052 26862
rect 9884 26850 10052 26852
rect 9884 26798 9998 26850
rect 10050 26798 10052 26850
rect 9884 26796 10052 26798
rect 9884 26290 9940 26796
rect 9996 26786 10052 26796
rect 9884 26238 9886 26290
rect 9938 26238 9940 26290
rect 9884 26226 9940 26238
rect 9996 26628 10052 26638
rect 9772 26114 9828 26124
rect 9996 25618 10052 26572
rect 10332 26628 10388 26908
rect 10668 26898 10724 26908
rect 10780 26740 10836 28140
rect 10332 26562 10388 26572
rect 10668 26684 10836 26740
rect 9996 25566 9998 25618
rect 10050 25566 10052 25618
rect 9996 25554 10052 25566
rect 10108 26402 10164 26414
rect 10108 26350 10110 26402
rect 10162 26350 10164 26402
rect 9100 25454 9102 25506
rect 9154 25454 9156 25506
rect 8988 25396 9044 25406
rect 8988 16100 9044 25340
rect 9100 25284 9156 25454
rect 9100 25218 9156 25228
rect 10108 24164 10164 26350
rect 10556 26180 10612 26190
rect 10556 26086 10612 26124
rect 10108 24108 10388 24164
rect 10108 23940 10164 23950
rect 9660 23714 9716 23726
rect 9660 23662 9662 23714
rect 9714 23662 9716 23714
rect 9548 23268 9604 23278
rect 9660 23268 9716 23662
rect 9548 23266 9716 23268
rect 9548 23214 9550 23266
rect 9602 23214 9716 23266
rect 9548 23212 9716 23214
rect 9324 22372 9380 22382
rect 9548 22372 9604 23212
rect 9996 22484 10052 22494
rect 9324 22370 9604 22372
rect 9324 22318 9326 22370
rect 9378 22318 9604 22370
rect 9324 22316 9604 22318
rect 9772 22372 9828 22382
rect 9324 22306 9380 22316
rect 9772 22278 9828 22316
rect 9996 22370 10052 22428
rect 9996 22318 9998 22370
rect 10050 22318 10052 22370
rect 9996 22306 10052 22318
rect 9884 21812 9940 21822
rect 10108 21812 10164 23884
rect 10220 23826 10276 23838
rect 10220 23774 10222 23826
rect 10274 23774 10276 23826
rect 10220 23156 10276 23774
rect 10332 23268 10388 24108
rect 10668 24052 10724 26684
rect 10892 26628 10948 28476
rect 11004 28308 11060 32396
rect 11228 32340 11284 32350
rect 11228 32246 11284 32284
rect 11116 32004 11172 32014
rect 11172 31948 11284 32004
rect 11116 31938 11172 31948
rect 11116 31668 11172 31678
rect 11116 31574 11172 31612
rect 11228 31106 11284 31948
rect 11340 31780 11396 40572
rect 11564 38948 11620 42028
rect 11676 40514 11732 42476
rect 11900 42196 11956 42476
rect 11900 42130 11956 42140
rect 11788 42084 11844 42094
rect 11788 41858 11844 42028
rect 11788 41806 11790 41858
rect 11842 41806 11844 41858
rect 11788 41746 11844 41806
rect 11788 41694 11790 41746
rect 11842 41694 11844 41746
rect 11788 41682 11844 41694
rect 11676 40462 11678 40514
rect 11730 40462 11732 40514
rect 11676 40450 11732 40462
rect 11900 39732 11956 39742
rect 11900 39638 11956 39676
rect 11676 38948 11732 38958
rect 11564 38946 11732 38948
rect 11564 38894 11678 38946
rect 11730 38894 11732 38946
rect 11564 38892 11732 38894
rect 11676 38882 11732 38892
rect 11788 38162 11844 38174
rect 11788 38110 11790 38162
rect 11842 38110 11844 38162
rect 11564 37380 11620 37390
rect 11564 37266 11620 37324
rect 11564 37214 11566 37266
rect 11618 37214 11620 37266
rect 11564 37202 11620 37214
rect 11564 36596 11620 36606
rect 11564 35810 11620 36540
rect 11788 36036 11844 38110
rect 12012 36484 12068 43260
rect 12124 40402 12180 40414
rect 12124 40350 12126 40402
rect 12178 40350 12180 40402
rect 12124 39172 12180 40350
rect 12124 39106 12180 39116
rect 12012 36418 12068 36428
rect 11788 35970 11844 35980
rect 11564 35758 11566 35810
rect 11618 35758 11620 35810
rect 11564 34914 11620 35758
rect 11564 34862 11566 34914
rect 11618 34862 11620 34914
rect 11564 34850 11620 34862
rect 11900 34692 11956 34702
rect 11900 34690 12068 34692
rect 11900 34638 11902 34690
rect 11954 34638 12068 34690
rect 11900 34636 12068 34638
rect 11900 34626 11956 34636
rect 12012 34130 12068 34636
rect 12012 34078 12014 34130
rect 12066 34078 12068 34130
rect 11900 33348 11956 33358
rect 11676 33124 11732 33134
rect 11452 32676 11508 32686
rect 11452 32002 11508 32620
rect 11452 31950 11454 32002
rect 11506 31950 11508 32002
rect 11452 31938 11508 31950
rect 11564 32338 11620 32350
rect 11564 32286 11566 32338
rect 11618 32286 11620 32338
rect 11340 31724 11508 31780
rect 11228 31054 11230 31106
rect 11282 31054 11284 31106
rect 11228 31042 11284 31054
rect 11340 30100 11396 30110
rect 11340 30006 11396 30044
rect 11452 29988 11508 31724
rect 11452 29922 11508 29932
rect 11564 29764 11620 32286
rect 11004 28242 11060 28252
rect 11116 29708 11620 29764
rect 11116 28532 11172 29708
rect 11676 29652 11732 33068
rect 11900 31780 11956 33292
rect 12012 32564 12068 34078
rect 12236 34132 12292 44940
rect 12908 44324 12964 44334
rect 12908 44230 12964 44268
rect 12348 44100 12404 44110
rect 12348 43538 12404 44044
rect 12348 43486 12350 43538
rect 12402 43486 12404 43538
rect 12348 43474 12404 43486
rect 12460 43762 12516 43774
rect 12460 43710 12462 43762
rect 12514 43710 12516 43762
rect 12348 42530 12404 42542
rect 12348 42478 12350 42530
rect 12402 42478 12404 42530
rect 12348 42084 12404 42478
rect 12348 42018 12404 42028
rect 12348 39172 12404 39182
rect 12348 38834 12404 39116
rect 12348 38782 12350 38834
rect 12402 38782 12404 38834
rect 12348 38770 12404 38782
rect 12460 38668 12516 43710
rect 12348 38612 12516 38668
rect 12572 43538 12628 43550
rect 12572 43486 12574 43538
rect 12626 43486 12628 43538
rect 12572 42978 12628 43486
rect 12796 43540 12852 43550
rect 12796 43446 12852 43484
rect 13132 43204 13188 53788
rect 13244 53732 13300 54462
rect 13244 53666 13300 53676
rect 13804 53396 13860 55244
rect 13916 54514 13972 55916
rect 13916 54462 13918 54514
rect 13970 54462 13972 54514
rect 13916 53620 13972 54462
rect 14028 54180 14084 56140
rect 14476 54852 14532 62132
rect 14924 62132 14980 62142
rect 14700 61458 14756 61470
rect 14700 61406 14702 61458
rect 14754 61406 14756 61458
rect 14700 61012 14756 61406
rect 14812 61012 14868 61022
rect 14700 61010 14868 61012
rect 14700 60958 14814 61010
rect 14866 60958 14868 61010
rect 14700 60956 14868 60958
rect 14812 60676 14868 60956
rect 14812 60610 14868 60620
rect 14588 57650 14644 57662
rect 14588 57598 14590 57650
rect 14642 57598 14644 57650
rect 14588 57092 14644 57598
rect 14700 57652 14756 57662
rect 14700 57558 14756 57596
rect 14588 57026 14644 57036
rect 14924 56420 14980 62076
rect 14924 56354 14980 56364
rect 14476 54786 14532 54796
rect 14252 54628 14308 54638
rect 14140 54180 14196 54190
rect 14028 54124 14140 54180
rect 14140 54114 14196 54124
rect 14028 53620 14084 53630
rect 13916 53564 14028 53620
rect 14028 53554 14084 53564
rect 13692 53340 13860 53396
rect 13580 53172 13636 53182
rect 13356 52164 13412 52174
rect 13356 52070 13412 52108
rect 13580 52164 13636 53116
rect 13580 52050 13636 52108
rect 13580 51998 13582 52050
rect 13634 51998 13636 52050
rect 13580 51986 13636 51998
rect 13692 52162 13748 53340
rect 13804 53172 13860 53182
rect 14252 53172 14308 54572
rect 15036 54628 15092 64428
rect 15484 64390 15540 64428
rect 15596 63700 15652 63710
rect 15260 62692 15316 62702
rect 15260 62578 15316 62636
rect 15260 62526 15262 62578
rect 15314 62526 15316 62578
rect 15260 62514 15316 62526
rect 15596 62578 15652 63644
rect 15596 62526 15598 62578
rect 15650 62526 15652 62578
rect 15596 62356 15652 62526
rect 15596 62290 15652 62300
rect 15372 62244 15428 62254
rect 15372 61348 15428 62188
rect 15484 61572 15540 61582
rect 15484 61478 15540 61516
rect 15372 61292 15540 61348
rect 15372 61124 15428 61134
rect 15260 60788 15316 60798
rect 15260 60674 15316 60732
rect 15260 60622 15262 60674
rect 15314 60622 15316 60674
rect 15260 57988 15316 60622
rect 15260 57922 15316 57932
rect 15260 57652 15316 57662
rect 15036 54562 15092 54572
rect 15148 57540 15204 57550
rect 14700 54404 14756 54414
rect 14700 54402 15092 54404
rect 14700 54350 14702 54402
rect 14754 54350 15092 54402
rect 14700 54348 15092 54350
rect 14700 54338 14756 54348
rect 14924 54180 14980 54190
rect 14812 53732 14868 53742
rect 14812 53638 14868 53676
rect 13804 53170 14308 53172
rect 13804 53118 13806 53170
rect 13858 53118 14254 53170
rect 14306 53118 14308 53170
rect 13804 53116 14308 53118
rect 13804 53106 13860 53116
rect 13692 52110 13694 52162
rect 13746 52110 13748 52162
rect 13468 50036 13524 50046
rect 13692 50036 13748 52110
rect 13916 52164 13972 52174
rect 13916 51266 13972 52108
rect 13916 51214 13918 51266
rect 13970 51214 13972 51266
rect 13916 51202 13972 51214
rect 13468 50034 13748 50036
rect 13468 49982 13470 50034
rect 13522 49982 13748 50034
rect 13468 49980 13748 49982
rect 13916 51044 13972 51054
rect 13468 49924 13524 49980
rect 13468 49858 13524 49868
rect 13804 49812 13860 49822
rect 13804 49718 13860 49756
rect 13580 49026 13636 49038
rect 13580 48974 13582 49026
rect 13634 48974 13636 49026
rect 13580 48356 13636 48974
rect 13804 48916 13860 48954
rect 13804 48850 13860 48860
rect 13580 48290 13636 48300
rect 13804 48692 13860 48702
rect 13468 48242 13524 48254
rect 13468 48190 13470 48242
rect 13522 48190 13524 48242
rect 13356 47796 13412 47806
rect 13468 47796 13524 48190
rect 13412 47740 13524 47796
rect 13580 48132 13636 48142
rect 13356 47730 13412 47740
rect 13356 47124 13412 47134
rect 13356 45332 13412 47068
rect 13468 46900 13524 46910
rect 13468 46806 13524 46844
rect 13356 45106 13412 45276
rect 13356 45054 13358 45106
rect 13410 45054 13412 45106
rect 13356 45042 13412 45054
rect 13580 46002 13636 48076
rect 13804 47012 13860 48636
rect 13916 47572 13972 50988
rect 14028 48132 14084 53116
rect 14252 53106 14308 53116
rect 14700 53620 14756 53630
rect 14140 52948 14196 52958
rect 14140 49026 14196 52892
rect 14476 52948 14532 52958
rect 14476 52854 14532 52892
rect 14700 52164 14756 53564
rect 14812 52164 14868 52174
rect 14700 52162 14868 52164
rect 14700 52110 14814 52162
rect 14866 52110 14868 52162
rect 14700 52108 14868 52110
rect 14812 52098 14868 52108
rect 14140 48974 14142 49026
rect 14194 48974 14196 49026
rect 14140 48916 14196 48974
rect 14140 48850 14196 48860
rect 14252 49698 14308 49710
rect 14252 49646 14254 49698
rect 14306 49646 14308 49698
rect 14252 48804 14308 49646
rect 14812 49698 14868 49710
rect 14812 49646 14814 49698
rect 14866 49646 14868 49698
rect 14812 49586 14868 49646
rect 14812 49534 14814 49586
rect 14866 49534 14868 49586
rect 14812 49522 14868 49534
rect 14476 48916 14532 48926
rect 14700 48916 14756 48926
rect 14476 48914 14756 48916
rect 14476 48862 14478 48914
rect 14530 48862 14702 48914
rect 14754 48862 14756 48914
rect 14476 48860 14756 48862
rect 14476 48850 14532 48860
rect 14700 48850 14756 48860
rect 14252 48710 14308 48748
rect 14812 48802 14868 48814
rect 14812 48750 14814 48802
rect 14866 48750 14868 48802
rect 14812 48468 14868 48750
rect 14140 48412 14868 48468
rect 14140 48354 14196 48412
rect 14140 48302 14142 48354
rect 14194 48302 14196 48354
rect 14140 48290 14196 48302
rect 14028 48076 14756 48132
rect 13916 47516 14420 47572
rect 14364 47346 14420 47516
rect 14588 47460 14644 47470
rect 14364 47294 14366 47346
rect 14418 47294 14420 47346
rect 14364 47282 14420 47294
rect 14476 47458 14644 47460
rect 14476 47406 14590 47458
rect 14642 47406 14644 47458
rect 14476 47404 14644 47406
rect 13804 46956 14196 47012
rect 13692 46900 13748 46910
rect 14140 46900 14196 46956
rect 13748 46844 13860 46900
rect 13692 46834 13748 46844
rect 13804 46786 13860 46844
rect 14140 46898 14420 46900
rect 14140 46846 14142 46898
rect 14194 46846 14420 46898
rect 14140 46844 14420 46846
rect 14140 46834 14196 46844
rect 13804 46734 13806 46786
rect 13858 46734 13860 46786
rect 13804 46722 13860 46734
rect 13580 45950 13582 46002
rect 13634 45950 13636 46002
rect 13356 44882 13412 44894
rect 13356 44830 13358 44882
rect 13410 44830 13412 44882
rect 13356 44100 13412 44830
rect 13580 44324 13636 45950
rect 14140 45892 14196 45902
rect 14140 45798 14196 45836
rect 13692 45780 13748 45790
rect 13692 45218 13748 45724
rect 14364 45556 14420 46844
rect 14476 45780 14532 47404
rect 14588 47394 14644 47404
rect 14476 45686 14532 45724
rect 14364 45500 14532 45556
rect 13692 45166 13694 45218
rect 13746 45166 13748 45218
rect 13692 44660 13748 45166
rect 14140 44994 14196 45006
rect 14140 44942 14142 44994
rect 14194 44942 14196 44994
rect 14140 44884 14196 44942
rect 14140 44818 14196 44828
rect 13692 44604 14420 44660
rect 13692 44546 13748 44604
rect 13692 44494 13694 44546
rect 13746 44494 13748 44546
rect 13692 44482 13748 44494
rect 13580 44258 13636 44268
rect 13916 44436 13972 44446
rect 13356 44034 13412 44044
rect 13804 44212 13860 44222
rect 13356 43764 13412 43774
rect 12572 42926 12574 42978
rect 12626 42926 12628 42978
rect 12572 38668 12628 42926
rect 12796 43148 13188 43204
rect 13244 43426 13300 43438
rect 13244 43374 13246 43426
rect 13298 43374 13300 43426
rect 12796 42868 12852 43148
rect 13020 42980 13076 42990
rect 13244 42980 13300 43374
rect 13020 42978 13300 42980
rect 13020 42926 13022 42978
rect 13074 42926 13300 42978
rect 13020 42924 13300 42926
rect 13020 42914 13076 42924
rect 12796 42774 12852 42812
rect 12908 42084 12964 42094
rect 12908 40514 12964 42028
rect 12908 40462 12910 40514
rect 12962 40462 12964 40514
rect 12908 40450 12964 40462
rect 13356 38668 13412 43708
rect 13468 43540 13524 43550
rect 13692 43540 13748 43550
rect 13524 43538 13748 43540
rect 13524 43486 13694 43538
rect 13746 43486 13748 43538
rect 13524 43484 13748 43486
rect 13468 42642 13524 43484
rect 13692 43474 13748 43484
rect 13804 42754 13860 44156
rect 13916 44210 13972 44380
rect 14028 44436 14084 44446
rect 14028 44434 14196 44436
rect 14028 44382 14030 44434
rect 14082 44382 14196 44434
rect 14028 44380 14196 44382
rect 14028 44370 14084 44380
rect 13916 44158 13918 44210
rect 13970 44158 13972 44210
rect 13916 44146 13972 44158
rect 14028 43540 14084 43550
rect 14028 43446 14084 43484
rect 14140 43538 14196 44380
rect 14364 44210 14420 44604
rect 14364 44158 14366 44210
rect 14418 44158 14420 44210
rect 14364 44146 14420 44158
rect 14476 43988 14532 45500
rect 14588 45332 14644 45342
rect 14588 44660 14644 45276
rect 14588 44594 14644 44604
rect 14588 44322 14644 44334
rect 14588 44270 14590 44322
rect 14642 44270 14644 44322
rect 14588 44212 14644 44270
rect 14588 44146 14644 44156
rect 14700 43988 14756 48076
rect 14812 45892 14868 45902
rect 14812 45798 14868 45836
rect 14140 43486 14142 43538
rect 14194 43486 14196 43538
rect 14140 43474 14196 43486
rect 14252 43932 14476 43988
rect 14252 43538 14308 43932
rect 14476 43922 14532 43932
rect 14588 43932 14756 43988
rect 14476 43764 14532 43774
rect 14252 43486 14254 43538
rect 14306 43486 14308 43538
rect 14252 43474 14308 43486
rect 14364 43762 14532 43764
rect 14364 43710 14478 43762
rect 14530 43710 14532 43762
rect 14364 43708 14532 43710
rect 13804 42702 13806 42754
rect 13858 42702 13860 42754
rect 13804 42690 13860 42702
rect 13468 42590 13470 42642
rect 13522 42590 13524 42642
rect 13468 42578 13524 42590
rect 14252 39732 14308 39742
rect 14364 39732 14420 43708
rect 14476 43698 14532 43708
rect 14252 39730 14420 39732
rect 14252 39678 14254 39730
rect 14306 39678 14420 39730
rect 14252 39676 14420 39678
rect 14252 39666 14308 39676
rect 13468 39620 13524 39630
rect 13468 38948 13524 39564
rect 13468 38882 13524 38892
rect 12572 38612 12852 38668
rect 12348 37378 12404 38612
rect 12348 37326 12350 37378
rect 12402 37326 12404 37378
rect 12348 37314 12404 37326
rect 12572 36596 12628 36606
rect 12572 36502 12628 36540
rect 12236 34066 12292 34076
rect 12460 34692 12516 34702
rect 12460 34130 12516 34636
rect 12460 34078 12462 34130
rect 12514 34078 12516 34130
rect 12236 33348 12292 33358
rect 12236 33254 12292 33292
rect 12124 33124 12180 33134
rect 12460 33124 12516 34078
rect 12684 34244 12740 34254
rect 12684 33570 12740 34188
rect 12684 33518 12686 33570
rect 12738 33518 12740 33570
rect 12684 33506 12740 33518
rect 12572 33460 12628 33470
rect 12572 33346 12628 33404
rect 12572 33294 12574 33346
rect 12626 33294 12628 33346
rect 12572 33282 12628 33294
rect 12684 33348 12740 33358
rect 12684 33234 12740 33292
rect 12684 33182 12686 33234
rect 12738 33182 12740 33234
rect 12684 33170 12740 33182
rect 12460 33068 12628 33124
rect 12124 32786 12180 33068
rect 12124 32734 12126 32786
rect 12178 32734 12180 32786
rect 12124 32722 12180 32734
rect 12348 32564 12404 32574
rect 12012 32508 12348 32564
rect 12348 32470 12404 32508
rect 12348 32004 12404 32014
rect 11900 31724 12068 31780
rect 11900 31554 11956 31566
rect 11900 31502 11902 31554
rect 11954 31502 11956 31554
rect 11788 30884 11844 30894
rect 11788 30790 11844 30828
rect 11900 30212 11956 31502
rect 11340 29596 11732 29652
rect 11788 30156 11956 30212
rect 11228 29540 11284 29550
rect 11228 29446 11284 29484
rect 11228 28756 11284 28766
rect 11228 28642 11284 28700
rect 11228 28590 11230 28642
rect 11282 28590 11284 28642
rect 11228 28578 11284 28590
rect 11004 28084 11060 28094
rect 11004 27858 11060 28028
rect 11004 27806 11006 27858
rect 11058 27806 11060 27858
rect 11004 27794 11060 27806
rect 11116 27188 11172 28476
rect 11116 27122 11172 27132
rect 11340 27970 11396 29596
rect 11340 27918 11342 27970
rect 11394 27918 11396 27970
rect 11004 26964 11060 27002
rect 11004 26898 11060 26908
rect 10556 23996 10724 24052
rect 10780 26572 10948 26628
rect 10780 24722 10836 26572
rect 10780 24670 10782 24722
rect 10834 24670 10836 24722
rect 10556 23268 10612 23996
rect 10780 23940 10836 24670
rect 10780 23874 10836 23884
rect 10892 26402 10948 26414
rect 10892 26350 10894 26402
rect 10946 26350 10948 26402
rect 10892 25284 10948 26350
rect 10668 23826 10724 23838
rect 10668 23774 10670 23826
rect 10722 23774 10724 23826
rect 10668 23716 10724 23774
rect 10780 23716 10836 23726
rect 10668 23660 10780 23716
rect 10780 23650 10836 23660
rect 10892 23714 10948 25228
rect 11116 24948 11172 24958
rect 11172 24892 11284 24948
rect 11116 24854 11172 24892
rect 11116 24500 11172 24510
rect 11116 24052 11172 24444
rect 11228 24164 11284 24892
rect 11340 24276 11396 27918
rect 11452 29204 11508 29214
rect 11452 24500 11508 29148
rect 11788 28868 11844 30156
rect 12012 29650 12068 31724
rect 12236 31556 12292 31566
rect 12348 31556 12404 31948
rect 12236 31554 12404 31556
rect 12236 31502 12238 31554
rect 12290 31502 12404 31554
rect 12236 31500 12404 31502
rect 12236 31490 12292 31500
rect 12124 30996 12180 31006
rect 12124 30210 12180 30940
rect 12124 30158 12126 30210
rect 12178 30158 12180 30210
rect 12124 30146 12180 30158
rect 12236 30994 12292 31006
rect 12236 30942 12238 30994
rect 12290 30942 12292 30994
rect 12012 29598 12014 29650
rect 12066 29598 12068 29650
rect 11900 29428 11956 29438
rect 11900 29334 11956 29372
rect 11564 28812 11844 28868
rect 11564 28644 11620 28812
rect 12012 28756 12068 29598
rect 12236 29426 12292 30942
rect 12572 30996 12628 33068
rect 12796 31668 12852 38612
rect 13132 38612 13412 38668
rect 13804 38612 13860 38622
rect 13132 33348 13188 38612
rect 13132 33282 13188 33292
rect 13468 38556 13804 38612
rect 12796 31602 12852 31612
rect 13356 32004 13412 32014
rect 13244 30996 13300 31006
rect 12572 30940 12740 30996
rect 12572 30100 12628 30110
rect 12236 29374 12238 29426
rect 12290 29374 12292 29426
rect 12236 29092 12292 29374
rect 12460 30098 12628 30100
rect 12460 30046 12574 30098
rect 12626 30046 12628 30098
rect 12460 30044 12628 30046
rect 12460 29428 12516 30044
rect 12572 30034 12628 30044
rect 12684 30098 12740 30940
rect 12908 30994 13300 30996
rect 12908 30942 13246 30994
rect 13298 30942 13300 30994
rect 12908 30940 13300 30942
rect 12908 30210 12964 30940
rect 13244 30930 13300 30940
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30146 12964 30158
rect 12684 30046 12686 30098
rect 12738 30046 12740 30098
rect 12572 29652 12628 29662
rect 12684 29652 12740 30046
rect 12572 29650 13188 29652
rect 12572 29598 12574 29650
rect 12626 29598 13188 29650
rect 12572 29596 13188 29598
rect 12572 29586 12628 29596
rect 12460 29372 12852 29428
rect 12236 29036 12516 29092
rect 11564 28530 11620 28588
rect 11564 28478 11566 28530
rect 11618 28478 11620 28530
rect 11564 28466 11620 28478
rect 11900 28754 12068 28756
rect 11900 28702 12014 28754
rect 12066 28702 12068 28754
rect 11900 28700 12068 28702
rect 11564 28196 11620 28206
rect 11564 28082 11620 28140
rect 11788 28084 11844 28094
rect 11564 28030 11566 28082
rect 11618 28030 11620 28082
rect 11564 28018 11620 28030
rect 11676 28028 11788 28084
rect 11676 27970 11732 28028
rect 11788 28018 11844 28028
rect 11676 27918 11678 27970
rect 11730 27918 11732 27970
rect 11676 27906 11732 27918
rect 11788 27858 11844 27870
rect 11788 27806 11790 27858
rect 11842 27806 11844 27858
rect 11788 27636 11844 27806
rect 11788 27570 11844 27580
rect 11676 27300 11788 27412
rect 11900 27300 11956 28700
rect 12012 28690 12068 28700
rect 12236 28196 12292 28206
rect 12124 28140 12236 28196
rect 12124 27972 12180 28140
rect 12236 28130 12292 28140
rect 12348 28084 12404 28094
rect 12460 28084 12516 29036
rect 12796 28196 12852 29372
rect 12796 28130 12852 28140
rect 12572 28084 12628 28094
rect 12460 28082 12628 28084
rect 12460 28030 12574 28082
rect 12626 28030 12628 28082
rect 12460 28028 12628 28030
rect 12348 27990 12404 28028
rect 12572 28018 12628 28028
rect 12124 27916 12292 27972
rect 12012 27860 12068 27870
rect 12012 27766 12068 27804
rect 11676 27244 11956 27300
rect 11676 26908 11732 27244
rect 12012 27188 12068 27198
rect 11676 26852 11844 26908
rect 11788 25618 11844 26852
rect 12012 26516 12068 27132
rect 12124 26962 12180 26974
rect 12124 26910 12126 26962
rect 12178 26910 12180 26962
rect 12124 26908 12180 26910
rect 12124 26842 12180 26852
rect 12012 26460 12180 26516
rect 11788 25566 11790 25618
rect 11842 25566 11844 25618
rect 11788 25396 11844 25566
rect 12124 25506 12180 26460
rect 12124 25454 12126 25506
rect 12178 25454 12180 25506
rect 12124 25442 12180 25454
rect 12236 25508 12292 27916
rect 12348 27860 12404 27870
rect 12348 27188 12404 27804
rect 12908 27858 12964 27870
rect 12908 27806 12910 27858
rect 12962 27806 12964 27858
rect 12460 27748 12516 27758
rect 12460 27654 12516 27692
rect 12348 27074 12404 27132
rect 12348 27022 12350 27074
rect 12402 27022 12404 27074
rect 12348 27010 12404 27022
rect 12796 27636 12852 27646
rect 12796 27074 12852 27580
rect 12908 27186 12964 27806
rect 12908 27134 12910 27186
rect 12962 27134 12964 27186
rect 12908 27122 12964 27134
rect 13020 27188 13076 27198
rect 12796 27022 12798 27074
rect 12850 27022 12852 27074
rect 12796 27010 12852 27022
rect 12684 26964 12740 26974
rect 12572 26852 12628 26862
rect 12572 26758 12628 26796
rect 12460 26404 12516 26414
rect 12460 26402 12628 26404
rect 12460 26350 12462 26402
rect 12514 26350 12628 26402
rect 12460 26348 12628 26350
rect 12460 26338 12516 26348
rect 12236 25452 12404 25508
rect 11788 25284 11844 25340
rect 12236 25284 12292 25294
rect 11788 25282 12292 25284
rect 11788 25230 12238 25282
rect 12290 25230 12292 25282
rect 11788 25228 12292 25230
rect 12236 25218 12292 25228
rect 11452 24434 11508 24444
rect 11788 24948 11844 24958
rect 11340 24220 11732 24276
rect 11228 24108 11508 24164
rect 11116 23996 11284 24052
rect 10892 23662 10894 23714
rect 10946 23662 10948 23714
rect 10892 23650 10948 23662
rect 11004 23714 11060 23726
rect 11004 23662 11006 23714
rect 11058 23662 11060 23714
rect 10556 23212 10948 23268
rect 10332 23202 10388 23212
rect 10220 23090 10276 23100
rect 10780 23044 10836 23054
rect 10556 22930 10612 22942
rect 10556 22878 10558 22930
rect 10610 22878 10612 22930
rect 10556 22260 10612 22878
rect 9772 21756 9884 21812
rect 9660 21476 9716 21486
rect 9548 21474 9716 21476
rect 9548 21422 9662 21474
rect 9714 21422 9716 21474
rect 9548 21420 9716 21422
rect 9212 19010 9268 19022
rect 9212 18958 9214 19010
rect 9266 18958 9268 19010
rect 9212 18452 9268 18958
rect 9212 18386 9268 18396
rect 9548 17556 9604 21420
rect 9660 21410 9716 21420
rect 9772 19234 9828 21756
rect 9884 21746 9940 21756
rect 9996 21756 10164 21812
rect 10220 22204 10612 22260
rect 10668 22258 10724 22270
rect 10668 22206 10670 22258
rect 10722 22206 10724 22258
rect 10220 21810 10276 22204
rect 10220 21758 10222 21810
rect 10274 21758 10276 21810
rect 9884 20132 9940 20142
rect 9996 20132 10052 21756
rect 10220 21746 10276 21758
rect 10668 21362 10724 22206
rect 10780 21810 10836 22988
rect 10780 21758 10782 21810
rect 10834 21758 10836 21810
rect 10780 21746 10836 21758
rect 10892 21812 10948 23212
rect 10892 21718 10948 21756
rect 10668 21310 10670 21362
rect 10722 21310 10724 21362
rect 10668 20916 10724 21310
rect 9884 20130 10052 20132
rect 9884 20078 9886 20130
rect 9938 20078 10052 20130
rect 9884 20076 10052 20078
rect 10108 20860 10724 20916
rect 10108 20802 10164 20860
rect 10108 20750 10110 20802
rect 10162 20750 10164 20802
rect 9884 20066 9940 20076
rect 9772 19182 9774 19234
rect 9826 19182 9828 19234
rect 9772 18674 9828 19182
rect 9772 18622 9774 18674
rect 9826 18622 9828 18674
rect 9772 18452 9828 18622
rect 9884 19908 9940 19918
rect 9884 19122 9940 19852
rect 9996 19796 10052 19806
rect 9996 19702 10052 19740
rect 9884 19070 9886 19122
rect 9938 19070 9940 19122
rect 9884 18564 9940 19070
rect 9884 18498 9940 18508
rect 9772 18386 9828 18396
rect 10108 18450 10164 20750
rect 10556 20692 10612 20702
rect 10332 20690 10612 20692
rect 10332 20638 10558 20690
rect 10610 20638 10612 20690
rect 10332 20636 10612 20638
rect 10332 19234 10388 20636
rect 10556 20626 10612 20636
rect 11004 20132 11060 23662
rect 11116 23714 11172 23726
rect 11116 23662 11118 23714
rect 11170 23662 11172 23714
rect 11116 22484 11172 23662
rect 11116 22418 11172 22428
rect 11228 20804 11284 23996
rect 11452 23938 11508 24108
rect 11452 23886 11454 23938
rect 11506 23886 11508 23938
rect 11452 23874 11508 23886
rect 11340 23716 11396 23726
rect 11340 23622 11396 23660
rect 11004 20066 11060 20076
rect 11116 20748 11284 20804
rect 11340 23268 11396 23278
rect 10556 20018 10612 20030
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 10556 19796 10612 19966
rect 11116 19908 11172 20748
rect 11116 19814 11172 19852
rect 11228 20580 11284 20590
rect 10332 19182 10334 19234
rect 10386 19182 10388 19234
rect 10332 18676 10388 19182
rect 10444 19236 10500 19246
rect 10444 19010 10500 19180
rect 10444 18958 10446 19010
rect 10498 18958 10500 19010
rect 10444 18946 10500 18958
rect 10444 18676 10500 18686
rect 10332 18620 10444 18676
rect 10444 18610 10500 18620
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18386 10164 18398
rect 10332 18452 10388 18462
rect 10332 18358 10388 18396
rect 10556 18450 10612 19740
rect 11228 19234 11284 20524
rect 11340 19460 11396 23212
rect 11564 22370 11620 24220
rect 11676 23938 11732 24220
rect 11676 23886 11678 23938
rect 11730 23886 11732 23938
rect 11676 23874 11732 23886
rect 11564 22318 11566 22370
rect 11618 22318 11620 22370
rect 11564 22306 11620 22318
rect 11676 23156 11732 23166
rect 11676 22370 11732 23100
rect 11788 23154 11844 24892
rect 12348 24276 12404 25452
rect 12460 25284 12516 25294
rect 12460 25190 12516 25228
rect 11900 24220 12404 24276
rect 11900 23938 11956 24220
rect 11900 23886 11902 23938
rect 11954 23886 11956 23938
rect 11900 23874 11956 23886
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 23090 11844 23102
rect 11788 22484 11844 22494
rect 11788 22390 11844 22428
rect 11676 22318 11678 22370
rect 11730 22318 11732 22370
rect 11676 22306 11732 22318
rect 11900 22372 11956 22382
rect 11900 22278 11956 22316
rect 12012 22370 12068 24220
rect 12236 24052 12292 24062
rect 12124 23940 12180 23950
rect 12124 23846 12180 23884
rect 12236 23042 12292 23996
rect 12572 23548 12628 26348
rect 12684 26402 12740 26908
rect 13020 26964 13076 27132
rect 13020 26898 13076 26908
rect 12684 26350 12686 26402
rect 12738 26350 12740 26402
rect 12684 26338 12740 26350
rect 12796 24834 12852 24846
rect 12796 24782 12798 24834
rect 12850 24782 12852 24834
rect 12796 23940 12852 24782
rect 12572 23492 12740 23548
rect 12236 22990 12238 23042
rect 12290 22990 12292 23042
rect 12236 22978 12292 22990
rect 12684 23044 12740 23492
rect 12796 23156 12852 23884
rect 13132 23268 13188 29596
rect 13244 27748 13300 27758
rect 13244 26290 13300 27692
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 26226 13300 26238
rect 12796 23062 12852 23100
rect 12908 23212 13132 23268
rect 12684 22978 12740 22988
rect 12012 22318 12014 22370
rect 12066 22318 12068 22370
rect 12012 22306 12068 22318
rect 12124 22930 12180 22942
rect 12124 22878 12126 22930
rect 12178 22878 12180 22930
rect 11452 21812 11508 21822
rect 11452 21718 11508 21756
rect 12124 20580 12180 22878
rect 12908 22482 12964 23212
rect 13132 23202 13188 23212
rect 13356 23266 13412 31948
rect 13468 31780 13524 38556
rect 13804 38546 13860 38556
rect 14252 37156 14308 37166
rect 14476 37156 14532 37166
rect 14252 36594 14308 37100
rect 14252 36542 14254 36594
rect 14306 36542 14308 36594
rect 14252 36530 14308 36542
rect 14364 37154 14532 37156
rect 14364 37102 14478 37154
rect 14530 37102 14532 37154
rect 14364 37100 14532 37102
rect 14364 34356 14420 37100
rect 14476 37090 14532 37100
rect 14588 37044 14644 43932
rect 14700 39060 14756 39070
rect 14700 38050 14756 39004
rect 14924 38612 14980 54124
rect 15036 53842 15092 54348
rect 15036 53790 15038 53842
rect 15090 53790 15092 53842
rect 15036 53778 15092 53790
rect 15148 53284 15204 57484
rect 15260 57204 15316 57596
rect 15372 57428 15428 61068
rect 15484 57652 15540 61292
rect 15596 61124 15652 61134
rect 15596 60788 15652 61068
rect 15596 60694 15652 60732
rect 15484 57558 15540 57596
rect 15708 57652 15764 66110
rect 16492 65602 16548 65614
rect 16492 65550 16494 65602
rect 16546 65550 16548 65602
rect 15932 65492 15988 65502
rect 16492 65492 16548 65550
rect 15932 65490 16100 65492
rect 15932 65438 15934 65490
rect 15986 65438 16100 65490
rect 15932 65436 16100 65438
rect 15932 65426 15988 65436
rect 15820 65380 15876 65390
rect 15820 64820 15876 65324
rect 15932 64820 15988 64830
rect 15820 64818 15988 64820
rect 15820 64766 15934 64818
rect 15986 64766 15988 64818
rect 15820 64764 15988 64766
rect 15932 64754 15988 64764
rect 16044 64708 16100 65436
rect 16492 65426 16548 65436
rect 16380 65380 16436 65390
rect 16380 65286 16436 65324
rect 16044 64036 16100 64652
rect 16268 65266 16324 65278
rect 16268 65214 16270 65266
rect 16322 65214 16324 65266
rect 16268 64596 16324 65214
rect 16268 64530 16324 64540
rect 16044 63970 16100 63980
rect 16380 62916 16436 62926
rect 16380 62804 16436 62860
rect 15820 62748 16436 62804
rect 15820 60004 15876 62748
rect 15932 62580 15988 62590
rect 15932 62354 15988 62524
rect 16604 62580 16660 66220
rect 16716 64820 16772 71260
rect 17052 71316 17108 71326
rect 16716 64754 16772 64764
rect 16828 70084 16884 70094
rect 16828 63252 16884 70028
rect 17052 69524 17108 71260
rect 17164 70754 17220 70766
rect 17164 70702 17166 70754
rect 17218 70702 17220 70754
rect 17164 70644 17220 70702
rect 17164 70578 17220 70588
rect 17388 69748 17444 72268
rect 17948 72258 18004 72268
rect 18620 72546 18788 72548
rect 18620 72494 18734 72546
rect 18786 72494 18788 72546
rect 18620 72492 18788 72494
rect 18508 71650 18564 71662
rect 18508 71598 18510 71650
rect 18562 71598 18564 71650
rect 17724 71428 17780 71438
rect 17724 70420 17780 71372
rect 17836 70978 17892 70990
rect 17836 70926 17838 70978
rect 17890 70926 17892 70978
rect 17836 70644 17892 70926
rect 17836 70578 17892 70588
rect 18284 70978 18340 70990
rect 18284 70926 18286 70978
rect 18338 70926 18340 70978
rect 18284 70420 18340 70926
rect 18508 70756 18564 71598
rect 18508 70690 18564 70700
rect 17724 70364 17892 70420
rect 17724 70194 17780 70206
rect 17724 70142 17726 70194
rect 17778 70142 17780 70194
rect 17612 70084 17668 70094
rect 17724 70084 17780 70142
rect 17668 70028 17780 70084
rect 17612 70018 17668 70028
rect 17388 69692 17668 69748
rect 17052 69522 17444 69524
rect 17052 69470 17054 69522
rect 17106 69470 17444 69522
rect 17052 69468 17444 69470
rect 17052 69458 17108 69468
rect 17388 67842 17444 69468
rect 17388 67790 17390 67842
rect 17442 67790 17444 67842
rect 17388 67778 17444 67790
rect 17500 69522 17556 69534
rect 17500 69470 17502 69522
rect 17554 69470 17556 69522
rect 17388 67620 17444 67630
rect 17276 66948 17332 66958
rect 16940 66164 16996 66174
rect 16940 66162 17108 66164
rect 16940 66110 16942 66162
rect 16994 66110 17108 66162
rect 16940 66108 17108 66110
rect 16940 66098 16996 66108
rect 16940 64482 16996 64494
rect 16940 64430 16942 64482
rect 16994 64430 16996 64482
rect 16940 64036 16996 64430
rect 17052 64484 17108 66108
rect 17276 65380 17332 66892
rect 17388 66276 17444 67564
rect 17500 66948 17556 69470
rect 17500 66882 17556 66892
rect 17388 66210 17444 66220
rect 17612 65716 17668 69692
rect 17724 69524 17780 69534
rect 17836 69524 17892 70364
rect 18284 70194 18340 70364
rect 18396 70644 18452 70654
rect 18396 70306 18452 70588
rect 18396 70254 18398 70306
rect 18450 70254 18452 70306
rect 18396 70242 18452 70254
rect 18284 70142 18286 70194
rect 18338 70142 18340 70194
rect 18284 70130 18340 70142
rect 17724 69522 17892 69524
rect 17724 69470 17726 69522
rect 17778 69470 17892 69522
rect 17724 69468 17892 69470
rect 17724 69458 17780 69468
rect 18620 68068 18676 72492
rect 18732 72482 18788 72492
rect 18732 71874 18788 71886
rect 18732 71822 18734 71874
rect 18786 71822 18788 71874
rect 18732 71092 18788 71822
rect 18956 71092 19012 71102
rect 18732 71090 19012 71092
rect 18732 71038 18958 71090
rect 19010 71038 19012 71090
rect 18732 71036 19012 71038
rect 18956 71026 19012 71036
rect 18732 70420 18788 70430
rect 19068 70420 19124 73948
rect 19180 74228 19236 75740
rect 20076 75460 20132 75740
rect 20076 75404 20244 75460
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19180 73330 19236 74172
rect 19404 74788 19460 74798
rect 19404 74002 19460 74732
rect 20188 74226 20244 75404
rect 20300 74786 20356 76412
rect 20748 76402 20804 76412
rect 22428 76466 22484 76478
rect 22428 76414 22430 76466
rect 22482 76414 22484 76466
rect 22092 76356 22148 76366
rect 22092 76262 22148 76300
rect 20300 74734 20302 74786
rect 20354 74734 20356 74786
rect 20300 74722 20356 74734
rect 20524 75682 20580 75694
rect 20524 75630 20526 75682
rect 20578 75630 20580 75682
rect 20524 75460 20580 75630
rect 20188 74174 20190 74226
rect 20242 74174 20244 74226
rect 20188 74162 20244 74174
rect 20524 74228 20580 75404
rect 20636 75684 20692 75694
rect 20636 74786 20692 75628
rect 22428 75684 22484 76414
rect 23100 76354 23156 76974
rect 23100 76302 23102 76354
rect 23154 76302 23156 76354
rect 23100 76290 23156 76302
rect 24332 76580 24388 76590
rect 22428 75618 22484 75628
rect 23548 74900 23604 74910
rect 23212 74844 23548 74900
rect 20636 74734 20638 74786
rect 20690 74734 20692 74786
rect 20636 74722 20692 74734
rect 22764 74788 22820 74798
rect 22764 74694 22820 74732
rect 22764 74452 22820 74462
rect 20524 74162 20580 74172
rect 22316 74228 22372 74238
rect 22764 74228 22820 74396
rect 23212 74228 23268 74844
rect 23548 74806 23604 74844
rect 23996 74900 24052 74910
rect 23996 74806 24052 74844
rect 24332 74452 24388 76524
rect 24444 75794 24500 77420
rect 25788 77026 25844 79200
rect 25788 76974 25790 77026
rect 25842 76974 25844 77026
rect 25788 76962 25844 76974
rect 26348 77026 26404 77038
rect 26348 76974 26350 77026
rect 26402 76974 26404 77026
rect 26348 76578 26404 76974
rect 27580 76692 27636 79200
rect 29372 77252 29428 79200
rect 29372 77186 29428 77196
rect 30380 77252 30436 77262
rect 27580 76626 27636 76636
rect 29260 76692 29316 76702
rect 26348 76526 26350 76578
rect 26402 76526 26404 76578
rect 26348 76514 26404 76526
rect 27244 76468 27300 76478
rect 27244 76374 27300 76412
rect 28812 76466 28868 76478
rect 28812 76414 28814 76466
rect 28866 76414 28868 76466
rect 24444 75742 24446 75794
rect 24498 75742 24500 75794
rect 24444 75730 24500 75742
rect 24780 75908 24836 75918
rect 24668 74900 24724 74910
rect 24668 74806 24724 74844
rect 24332 74386 24388 74396
rect 22316 74134 22372 74172
rect 22428 74226 23156 74228
rect 22428 74174 22766 74226
rect 22818 74174 23156 74226
rect 22428 74172 23156 74174
rect 19404 73950 19406 74002
rect 19458 73950 19460 74002
rect 19404 73938 19460 73950
rect 19740 74004 19796 74014
rect 19740 73910 19796 73948
rect 20748 74004 20804 74014
rect 20804 73948 20916 74004
rect 20748 73910 20804 73948
rect 20860 73892 21252 73948
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 20636 73668 20692 73678
rect 19180 73278 19182 73330
rect 19234 73278 19236 73330
rect 19180 73266 19236 73278
rect 20300 73332 20356 73342
rect 20300 73330 20468 73332
rect 20300 73278 20302 73330
rect 20354 73278 20468 73330
rect 20300 73276 20468 73278
rect 20300 73266 20356 73276
rect 19292 73218 19348 73230
rect 19292 73166 19294 73218
rect 19346 73166 19348 73218
rect 19180 72660 19236 72670
rect 19180 70532 19236 72604
rect 19292 71316 19348 73166
rect 20300 72546 20356 72558
rect 20300 72494 20302 72546
rect 20354 72494 20356 72546
rect 19404 72434 19460 72446
rect 19404 72382 19406 72434
rect 19458 72382 19460 72434
rect 19404 71876 19460 72382
rect 19740 72436 19796 72446
rect 19740 72434 20132 72436
rect 19740 72382 19742 72434
rect 19794 72382 20132 72434
rect 19740 72380 20132 72382
rect 19740 72370 19796 72380
rect 20076 72324 20132 72380
rect 20076 72268 20244 72324
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 20188 71876 20244 72268
rect 19404 71820 19796 71876
rect 19740 71762 19796 71820
rect 19740 71710 19742 71762
rect 19794 71710 19796 71762
rect 19740 71698 19796 71710
rect 19964 71820 20244 71876
rect 19292 71260 19796 71316
rect 19628 70978 19684 70990
rect 19628 70926 19630 70978
rect 19682 70926 19684 70978
rect 19404 70866 19460 70878
rect 19404 70814 19406 70866
rect 19458 70814 19460 70866
rect 19404 70644 19460 70814
rect 19404 70578 19460 70588
rect 19180 70476 19348 70532
rect 19068 70364 19236 70420
rect 18732 69522 18788 70364
rect 18732 69470 18734 69522
rect 18786 69470 18788 69522
rect 18732 69458 18788 69470
rect 19068 70194 19124 70206
rect 19068 70142 19070 70194
rect 19122 70142 19124 70194
rect 18620 68012 19012 68068
rect 17948 67842 18004 67854
rect 17948 67790 17950 67842
rect 18002 67790 18004 67842
rect 17948 67172 18004 67790
rect 18620 67732 18676 67742
rect 18620 67730 18788 67732
rect 18620 67678 18622 67730
rect 18674 67678 18788 67730
rect 18620 67676 18788 67678
rect 18620 67666 18676 67676
rect 18172 67284 18228 67294
rect 17948 67106 18004 67116
rect 18060 67228 18172 67284
rect 17612 65650 17668 65660
rect 17276 65324 17444 65380
rect 17276 64596 17332 64606
rect 17276 64502 17332 64540
rect 17052 64418 17108 64428
rect 16940 63970 16996 63980
rect 16828 63186 16884 63196
rect 17276 63140 17332 63150
rect 17276 63046 17332 63084
rect 16828 62916 16884 62926
rect 16828 62822 16884 62860
rect 16268 62466 16324 62478
rect 16268 62414 16270 62466
rect 16322 62414 16324 62466
rect 15932 62302 15934 62354
rect 15986 62302 15988 62354
rect 15932 61124 15988 62302
rect 15932 61058 15988 61068
rect 16044 62356 16100 62366
rect 15820 59938 15876 59948
rect 15932 60900 15988 60910
rect 16044 60900 16100 62300
rect 16268 62188 16324 62414
rect 16604 62466 16660 62524
rect 16604 62414 16606 62466
rect 16658 62414 16660 62466
rect 16604 62402 16660 62414
rect 16716 62356 16772 62366
rect 17276 62356 17332 62366
rect 16716 62188 16772 62300
rect 16268 62132 16548 62188
rect 16492 61572 16548 62132
rect 16156 61460 16212 61470
rect 16156 61458 16436 61460
rect 16156 61406 16158 61458
rect 16210 61406 16436 61458
rect 16156 61404 16436 61406
rect 16156 61394 16212 61404
rect 16268 60900 16324 60910
rect 16044 60898 16324 60900
rect 16044 60846 16270 60898
rect 16322 60846 16324 60898
rect 16044 60844 16324 60846
rect 15708 57586 15764 57596
rect 15820 57762 15876 57774
rect 15820 57710 15822 57762
rect 15874 57710 15876 57762
rect 15820 57540 15876 57710
rect 15820 57474 15876 57484
rect 15372 57372 15540 57428
rect 15260 56978 15316 57148
rect 15260 56926 15262 56978
rect 15314 56926 15316 56978
rect 15260 56914 15316 56926
rect 15484 54628 15540 57372
rect 15708 57092 15764 57102
rect 15708 56998 15764 57036
rect 15932 57092 15988 60844
rect 16268 60834 16324 60844
rect 16380 60564 16436 61404
rect 16492 60788 16548 61516
rect 16492 60722 16548 60732
rect 16604 62132 16772 62188
rect 16940 62354 17332 62356
rect 16940 62302 17278 62354
rect 17330 62302 17332 62354
rect 16940 62300 17332 62302
rect 16604 60786 16660 62132
rect 16604 60734 16606 60786
rect 16658 60734 16660 60786
rect 16604 60722 16660 60734
rect 16940 60786 16996 62300
rect 17276 62290 17332 62300
rect 17388 62188 17444 65324
rect 17612 65156 17668 65166
rect 17612 64706 17668 65100
rect 17836 64932 17892 64942
rect 17612 64654 17614 64706
rect 17666 64654 17668 64706
rect 17612 64642 17668 64654
rect 17724 64930 17892 64932
rect 17724 64878 17838 64930
rect 17890 64878 17892 64930
rect 17724 64876 17892 64878
rect 17612 64484 17668 64494
rect 17612 64390 17668 64428
rect 17724 63250 17780 64876
rect 17836 64866 17892 64876
rect 17836 63364 17892 63374
rect 17836 63270 17892 63308
rect 17724 63198 17726 63250
rect 17778 63198 17780 63250
rect 17724 63186 17780 63198
rect 17500 63138 17556 63150
rect 17500 63086 17502 63138
rect 17554 63086 17556 63138
rect 17500 62916 17556 63086
rect 17500 62578 17556 62860
rect 17500 62526 17502 62578
rect 17554 62526 17556 62578
rect 17500 62514 17556 62526
rect 17836 62804 17892 62814
rect 17276 62132 17444 62188
rect 17612 62354 17668 62366
rect 17612 62302 17614 62354
rect 17666 62302 17668 62354
rect 16940 60734 16942 60786
rect 16994 60734 16996 60786
rect 16940 60722 16996 60734
rect 17164 61236 17220 61246
rect 16716 60674 16772 60686
rect 16716 60622 16718 60674
rect 16770 60622 16772 60674
rect 16716 60564 16772 60622
rect 16380 60508 16772 60564
rect 16940 60564 16996 60574
rect 16940 60002 16996 60508
rect 16940 59950 16942 60002
rect 16994 59950 16996 60002
rect 16492 59332 16548 59342
rect 16380 58548 16436 58558
rect 16380 58454 16436 58492
rect 16492 57650 16548 59276
rect 16716 58548 16772 58558
rect 16716 57764 16772 58492
rect 16940 57988 16996 59950
rect 17164 59890 17220 61180
rect 17164 59838 17166 59890
rect 17218 59838 17220 59890
rect 17164 59826 17220 59838
rect 16940 57922 16996 57932
rect 16492 57598 16494 57650
rect 16546 57598 16548 57650
rect 16492 57586 16548 57598
rect 16604 57762 16772 57764
rect 16604 57710 16718 57762
rect 16770 57710 16772 57762
rect 16604 57708 16772 57710
rect 15932 57026 15988 57036
rect 15708 56756 15764 56766
rect 15708 56662 15764 56700
rect 15820 56756 15876 56766
rect 16492 56756 16548 56766
rect 16604 56756 16660 57708
rect 16716 57698 16772 57708
rect 16828 57652 16884 57690
rect 16828 57586 16884 57596
rect 16828 57428 16884 57438
rect 15820 56754 16100 56756
rect 15820 56702 15822 56754
rect 15874 56702 16100 56754
rect 15820 56700 16100 56702
rect 15820 56690 15876 56700
rect 16044 55298 16100 56700
rect 16548 56700 16660 56756
rect 16716 57204 16772 57214
rect 16492 56690 16548 56700
rect 16716 56420 16772 57148
rect 16044 55246 16046 55298
rect 16098 55246 16100 55298
rect 15932 55188 15988 55198
rect 15932 55094 15988 55132
rect 15708 55076 15764 55086
rect 15484 54562 15540 54572
rect 15596 55074 15764 55076
rect 15596 55022 15710 55074
rect 15762 55022 15764 55074
rect 15596 55020 15764 55022
rect 15596 54404 15652 55020
rect 15708 55010 15764 55020
rect 15260 54348 15652 54404
rect 15260 53730 15316 54348
rect 15260 53678 15262 53730
rect 15314 53678 15316 53730
rect 15260 53666 15316 53678
rect 15484 53620 15540 53630
rect 15820 53620 15876 53630
rect 15484 53618 15820 53620
rect 15484 53566 15486 53618
rect 15538 53566 15820 53618
rect 15484 53564 15820 53566
rect 15484 53554 15540 53564
rect 15148 53228 15540 53284
rect 15260 52948 15316 52958
rect 15260 52854 15316 52892
rect 15260 52724 15316 52734
rect 15260 50428 15316 52668
rect 15372 52052 15428 52062
rect 15372 50708 15428 51996
rect 15372 50614 15428 50652
rect 15260 50372 15428 50428
rect 15148 49812 15204 49822
rect 15148 49810 15316 49812
rect 15148 49758 15150 49810
rect 15202 49758 15316 49810
rect 15148 49756 15316 49758
rect 15148 49746 15204 49756
rect 15260 49700 15316 49756
rect 15260 49634 15316 49644
rect 15036 49588 15092 49598
rect 15036 49026 15092 49532
rect 15036 48974 15038 49026
rect 15090 48974 15092 49026
rect 15036 48962 15092 48974
rect 15148 49586 15204 49598
rect 15148 49534 15150 49586
rect 15202 49534 15204 49586
rect 15148 48916 15204 49534
rect 15260 48916 15316 48926
rect 15148 48914 15316 48916
rect 15148 48862 15262 48914
rect 15314 48862 15316 48914
rect 15148 48860 15316 48862
rect 15260 48804 15316 48860
rect 15260 48738 15316 48748
rect 15148 47458 15204 47470
rect 15148 47406 15150 47458
rect 15202 47406 15204 47458
rect 15036 45892 15092 45902
rect 15148 45892 15204 47406
rect 15372 47346 15428 50372
rect 15372 47294 15374 47346
rect 15426 47294 15428 47346
rect 15372 47282 15428 47294
rect 15484 46900 15540 53228
rect 15596 53170 15652 53182
rect 15596 53118 15598 53170
rect 15650 53118 15652 53170
rect 15596 52274 15652 53118
rect 15708 52948 15764 52958
rect 15708 52854 15764 52892
rect 15820 52946 15876 53564
rect 16044 53060 16100 55246
rect 16604 56364 16772 56420
rect 16828 56866 16884 57372
rect 16828 56814 16830 56866
rect 16882 56814 16884 56866
rect 16604 53732 16660 56364
rect 16828 55300 16884 56814
rect 16940 56420 16996 56430
rect 16940 56306 16996 56364
rect 16940 56254 16942 56306
rect 16994 56254 16996 56306
rect 16940 56242 16996 56254
rect 17164 56196 17220 56206
rect 17052 56140 17164 56196
rect 16940 55300 16996 55310
rect 16828 55244 16940 55300
rect 16940 55206 16996 55244
rect 17052 55188 17108 56140
rect 17164 56130 17220 56140
rect 16828 54404 16884 54414
rect 17052 54404 17108 55132
rect 16828 54402 17108 54404
rect 16828 54350 16830 54402
rect 16882 54350 17108 54402
rect 16828 54348 17108 54350
rect 17164 55636 17220 55646
rect 16828 54338 16884 54348
rect 17164 54180 17220 55580
rect 17276 54628 17332 62132
rect 17612 61236 17668 62302
rect 17836 62188 17892 62748
rect 18060 62580 18116 67228
rect 18172 67218 18228 67228
rect 18620 67172 18676 67182
rect 18620 67078 18676 67116
rect 18284 67058 18340 67070
rect 18284 67006 18286 67058
rect 18338 67006 18340 67058
rect 18172 65268 18228 65278
rect 18172 64594 18228 65212
rect 18172 64542 18174 64594
rect 18226 64542 18228 64594
rect 18172 63700 18228 64542
rect 18172 63634 18228 63644
rect 18284 63588 18340 67006
rect 18620 65378 18676 65390
rect 18620 65326 18622 65378
rect 18674 65326 18676 65378
rect 18396 64596 18452 64606
rect 18396 64502 18452 64540
rect 18284 63522 18340 63532
rect 18396 64036 18452 64046
rect 18172 63364 18228 63374
rect 18172 63026 18228 63308
rect 18172 62974 18174 63026
rect 18226 62974 18228 63026
rect 18172 62962 18228 62974
rect 18396 63138 18452 63980
rect 18396 63086 18398 63138
rect 18450 63086 18452 63138
rect 18172 62804 18228 62814
rect 18396 62804 18452 63086
rect 18228 62748 18452 62804
rect 18620 64036 18676 65326
rect 18732 65044 18788 67676
rect 18956 66388 19012 68012
rect 19068 67284 19124 70142
rect 19180 69524 19236 70364
rect 19292 70308 19348 70476
rect 19628 70308 19684 70926
rect 19740 70980 19796 71260
rect 19852 71204 19908 71214
rect 19964 71204 20020 71820
rect 19852 71202 20020 71204
rect 19852 71150 19854 71202
rect 19906 71150 20020 71202
rect 19852 71148 20020 71150
rect 19852 71138 19908 71148
rect 20076 70980 20132 70990
rect 19740 70978 20132 70980
rect 19740 70926 20078 70978
rect 20130 70926 20132 70978
rect 19740 70924 20132 70926
rect 20076 70914 20132 70924
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19740 70308 19796 70318
rect 19628 70306 19796 70308
rect 19628 70254 19742 70306
rect 19794 70254 19796 70306
rect 19628 70252 19796 70254
rect 19292 70082 19348 70252
rect 19740 70242 19796 70252
rect 20188 70308 20244 70318
rect 20188 70214 20244 70252
rect 19292 70030 19294 70082
rect 19346 70030 19348 70082
rect 19292 70018 19348 70030
rect 19180 69468 19684 69524
rect 19068 67218 19124 67228
rect 19068 66388 19124 66398
rect 18956 66386 19124 66388
rect 18956 66334 19070 66386
rect 19122 66334 19124 66386
rect 18956 66332 19124 66334
rect 18956 65602 19012 66332
rect 19068 66322 19124 66332
rect 18956 65550 18958 65602
rect 19010 65550 19012 65602
rect 18956 65538 19012 65550
rect 18844 65268 18900 65278
rect 18844 65174 18900 65212
rect 18732 64988 19012 65044
rect 18956 64482 19012 64988
rect 18956 64430 18958 64482
rect 19010 64430 19012 64482
rect 18956 64418 19012 64430
rect 19068 64706 19124 64718
rect 19068 64654 19070 64706
rect 19122 64654 19124 64706
rect 19068 64260 19124 64654
rect 18956 64204 19124 64260
rect 19292 64706 19348 64718
rect 19292 64654 19294 64706
rect 19346 64654 19348 64706
rect 18956 64036 19012 64204
rect 18620 63980 19012 64036
rect 18172 62738 18228 62748
rect 18172 62580 18228 62590
rect 18060 62578 18452 62580
rect 18060 62526 18174 62578
rect 18226 62526 18452 62578
rect 18060 62524 18452 62526
rect 18172 62514 18228 62524
rect 17948 62356 18004 62366
rect 17948 62262 18004 62300
rect 18284 62354 18340 62366
rect 18284 62302 18286 62354
rect 18338 62302 18340 62354
rect 17836 62132 18004 62188
rect 17612 61170 17668 61180
rect 17836 60786 17892 60798
rect 17836 60734 17838 60786
rect 17890 60734 17892 60786
rect 17612 60676 17668 60686
rect 17612 60114 17668 60620
rect 17836 60676 17892 60734
rect 17836 60610 17892 60620
rect 17612 60062 17614 60114
rect 17666 60062 17668 60114
rect 17276 54562 17332 54572
rect 17388 59780 17444 59790
rect 17388 54404 17444 59724
rect 17500 59668 17556 59678
rect 17500 58548 17556 59612
rect 17612 58772 17668 60062
rect 17948 59556 18004 62132
rect 18284 61908 18340 62302
rect 18060 61852 18340 61908
rect 18060 61012 18116 61852
rect 18284 61684 18340 61694
rect 18396 61684 18452 62524
rect 18508 62244 18564 62254
rect 18620 62244 18676 63980
rect 19292 63924 19348 64654
rect 19516 64594 19572 64606
rect 19516 64542 19518 64594
rect 19570 64542 19572 64594
rect 19516 64484 19572 64542
rect 19516 64418 19572 64428
rect 19628 64034 19684 69468
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 20300 67396 20356 72494
rect 20412 69412 20468 73276
rect 20636 73330 20692 73612
rect 20636 73278 20638 73330
rect 20690 73278 20692 73330
rect 20636 72658 20692 73278
rect 20636 72606 20638 72658
rect 20690 72606 20692 72658
rect 20636 72594 20692 72606
rect 20748 72884 20804 72894
rect 20748 71874 20804 72828
rect 20748 71822 20750 71874
rect 20802 71822 20804 71874
rect 20748 71810 20804 71822
rect 20524 70868 20580 70878
rect 20524 70774 20580 70812
rect 20636 70082 20692 70094
rect 20636 70030 20638 70082
rect 20690 70030 20692 70082
rect 20636 69636 20692 70030
rect 20636 69570 20692 69580
rect 20412 69356 20804 69412
rect 20748 67956 20804 69356
rect 20636 67954 20804 67956
rect 20636 67902 20750 67954
rect 20802 67902 20804 67954
rect 20636 67900 20804 67902
rect 20300 67340 20580 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 20188 65490 20244 65502
rect 20188 65438 20190 65490
rect 20242 65438 20244 65490
rect 19852 65378 19908 65390
rect 19852 65326 19854 65378
rect 19906 65326 19908 65378
rect 19852 64820 19908 65326
rect 20188 65156 20244 65438
rect 20188 65090 20244 65100
rect 20412 65266 20468 65278
rect 20412 65214 20414 65266
rect 20466 65214 20468 65266
rect 20412 64930 20468 65214
rect 20412 64878 20414 64930
rect 20466 64878 20468 64930
rect 20412 64866 20468 64878
rect 19852 64764 20244 64820
rect 20188 64708 20244 64764
rect 20412 64708 20468 64718
rect 20188 64706 20468 64708
rect 20188 64654 20414 64706
rect 20466 64654 20468 64706
rect 20188 64652 20468 64654
rect 19740 64596 19796 64606
rect 19740 64502 19796 64540
rect 20076 64594 20132 64606
rect 20076 64542 20078 64594
rect 20130 64542 20132 64594
rect 20076 64484 20132 64542
rect 20076 64428 20244 64484
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19628 63982 19630 64034
rect 19682 63982 19684 64034
rect 19628 63970 19684 63982
rect 18844 63868 19348 63924
rect 18844 63362 18900 63868
rect 20188 63476 20244 64428
rect 19964 63420 20244 63476
rect 18844 63310 18846 63362
rect 18898 63310 18900 63362
rect 18844 63298 18900 63310
rect 19180 63364 19236 63374
rect 19180 63270 19236 63308
rect 19964 63364 20020 63420
rect 19964 63270 20020 63308
rect 20300 63252 20356 63262
rect 20300 63158 20356 63196
rect 18844 63140 18900 63150
rect 18564 62188 18676 62244
rect 18732 63084 18844 63140
rect 18508 62178 18564 62188
rect 18284 61682 18452 61684
rect 18284 61630 18286 61682
rect 18338 61630 18452 61682
rect 18284 61628 18452 61630
rect 18284 61618 18340 61628
rect 18060 60918 18116 60956
rect 18284 60564 18340 60574
rect 18060 59780 18116 59790
rect 18284 59780 18340 60508
rect 18116 59778 18340 59780
rect 18116 59726 18286 59778
rect 18338 59726 18340 59778
rect 18116 59724 18340 59726
rect 18060 59714 18116 59724
rect 18284 59714 18340 59724
rect 17948 59500 18340 59556
rect 18060 59332 18116 59342
rect 18060 59238 18116 59276
rect 17948 59220 18004 59230
rect 17836 59218 18004 59220
rect 17836 59166 17950 59218
rect 18002 59166 18004 59218
rect 17836 59164 18004 59166
rect 17724 59108 17780 59118
rect 17724 59014 17780 59052
rect 17612 58716 17780 58772
rect 17612 58548 17668 58558
rect 17500 58546 17668 58548
rect 17500 58494 17502 58546
rect 17554 58494 17614 58546
rect 17666 58494 17668 58546
rect 17500 58492 17668 58494
rect 17500 58454 17556 58492
rect 17612 58482 17668 58492
rect 17500 57764 17556 57774
rect 17500 57670 17556 57708
rect 17612 57652 17668 57662
rect 17500 57426 17556 57438
rect 17500 57374 17502 57426
rect 17554 57374 17556 57426
rect 17500 56754 17556 57374
rect 17500 56702 17502 56754
rect 17554 56702 17556 56754
rect 17500 56690 17556 56702
rect 17500 56196 17556 56206
rect 17500 56102 17556 56140
rect 17612 56084 17668 57596
rect 17724 57428 17780 58716
rect 17836 57652 17892 59164
rect 17948 59154 18004 59164
rect 18172 59220 18228 59230
rect 17836 57586 17892 57596
rect 17948 58658 18004 58670
rect 17948 58606 17950 58658
rect 18002 58606 18004 58658
rect 17948 57650 18004 58606
rect 18060 58436 18116 58446
rect 18060 58342 18116 58380
rect 18172 57874 18228 59164
rect 18172 57822 18174 57874
rect 18226 57822 18228 57874
rect 18172 57810 18228 57822
rect 17948 57598 17950 57650
rect 18002 57598 18004 57650
rect 17948 57586 18004 57598
rect 18284 57652 18340 59500
rect 18396 58772 18452 61628
rect 18508 61908 18564 61918
rect 18508 61012 18564 61852
rect 18620 61458 18676 61470
rect 18620 61406 18622 61458
rect 18674 61406 18676 61458
rect 18620 61236 18676 61406
rect 18620 61170 18676 61180
rect 18732 61346 18788 63084
rect 18844 63046 18900 63084
rect 19404 62916 19460 62926
rect 19404 62578 19460 62860
rect 19740 62916 19796 62954
rect 20188 62916 20244 62926
rect 19796 62914 20244 62916
rect 19796 62862 20190 62914
rect 20242 62862 20244 62914
rect 19796 62860 20244 62862
rect 19740 62850 19796 62860
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19404 62526 19406 62578
rect 19458 62526 19460 62578
rect 18732 61294 18734 61346
rect 18786 61294 18788 61346
rect 18508 60956 18676 61012
rect 18508 60788 18564 60798
rect 18508 60694 18564 60732
rect 18396 58706 18452 58716
rect 18620 58660 18676 60956
rect 18732 60564 18788 61294
rect 18844 62244 18900 62254
rect 18844 61348 18900 62188
rect 19404 61908 19460 62526
rect 20188 62188 20244 62860
rect 20412 62468 20468 64652
rect 19404 61842 19460 61852
rect 19852 62132 20244 62188
rect 20300 62412 20468 62468
rect 20300 62244 20356 62412
rect 20524 62188 20580 67340
rect 20636 67058 20692 67900
rect 20748 67890 20804 67900
rect 20636 67006 20638 67058
rect 20690 67006 20692 67058
rect 20636 66994 20692 67006
rect 20748 66946 20804 66958
rect 20748 66894 20750 66946
rect 20802 66894 20804 66946
rect 20748 65716 20804 66894
rect 20636 65660 20804 65716
rect 20636 64484 20692 65660
rect 20860 65602 20916 65614
rect 20860 65550 20862 65602
rect 20914 65550 20916 65602
rect 20748 65490 20804 65502
rect 20748 65438 20750 65490
rect 20802 65438 20804 65490
rect 20748 65380 20804 65438
rect 20860 65492 20916 65550
rect 20860 65426 20916 65436
rect 20972 65602 21028 65614
rect 20972 65550 20974 65602
rect 21026 65550 21028 65602
rect 20748 65314 20804 65324
rect 20972 64596 21028 65550
rect 20972 64530 21028 64540
rect 20636 64418 20692 64428
rect 21196 62188 21252 73892
rect 21980 73330 22036 73342
rect 21980 73278 21982 73330
rect 22034 73278 22036 73330
rect 21308 73218 21364 73230
rect 21308 73166 21310 73218
rect 21362 73166 21364 73218
rect 21308 71764 21364 73166
rect 21644 72436 21700 72446
rect 21644 72342 21700 72380
rect 21868 71764 21924 71774
rect 21308 71762 21924 71764
rect 21308 71710 21870 71762
rect 21922 71710 21924 71762
rect 21308 71708 21924 71710
rect 21868 71698 21924 71708
rect 21980 71428 22036 73278
rect 22428 73330 22484 74172
rect 22764 74162 22820 74172
rect 23100 73554 23156 74172
rect 23212 74114 23268 74172
rect 23884 74228 23940 74238
rect 23884 74134 23940 74172
rect 23212 74062 23214 74114
rect 23266 74062 23268 74114
rect 23212 74050 23268 74062
rect 23100 73502 23102 73554
rect 23154 73502 23156 73554
rect 23100 73490 23156 73502
rect 22428 73278 22430 73330
rect 22482 73278 22484 73330
rect 22428 72658 22484 73278
rect 23884 73330 23940 73342
rect 23884 73278 23886 73330
rect 23938 73278 23940 73330
rect 22652 73220 22708 73230
rect 23660 73220 23716 73230
rect 22428 72606 22430 72658
rect 22482 72606 22484 72658
rect 22428 72594 22484 72606
rect 22540 73218 22708 73220
rect 22540 73166 22654 73218
rect 22706 73166 22708 73218
rect 22540 73164 22708 73166
rect 22204 72546 22260 72558
rect 22204 72494 22206 72546
rect 22258 72494 22260 72546
rect 22204 72436 22260 72494
rect 22204 72370 22260 72380
rect 22428 71764 22484 71774
rect 21980 71362 22036 71372
rect 22316 71708 22428 71764
rect 21420 70756 21476 70766
rect 21420 70420 21476 70700
rect 22316 70420 22372 71708
rect 22428 71698 22484 71708
rect 22428 70980 22484 70990
rect 22540 70980 22596 73164
rect 22652 73154 22708 73164
rect 23548 73218 23716 73220
rect 23548 73166 23662 73218
rect 23714 73166 23716 73218
rect 23548 73164 23716 73166
rect 22876 72434 22932 72446
rect 22876 72382 22878 72434
rect 22930 72382 22932 72434
rect 22652 71762 22708 71774
rect 22652 71710 22654 71762
rect 22706 71710 22708 71762
rect 22652 71316 22708 71710
rect 22764 71764 22820 71774
rect 22764 71650 22820 71708
rect 22764 71598 22766 71650
rect 22818 71598 22820 71650
rect 22764 71586 22820 71598
rect 22652 71250 22708 71260
rect 22876 70980 22932 72382
rect 23548 71764 23604 73164
rect 23660 73154 23716 73164
rect 22428 70978 22596 70980
rect 22428 70926 22430 70978
rect 22482 70926 22596 70978
rect 22428 70924 22596 70926
rect 22652 70924 22932 70980
rect 22988 71708 23604 71764
rect 23884 72324 23940 73278
rect 24332 73330 24388 73342
rect 24332 73278 24334 73330
rect 24386 73278 24388 73330
rect 24332 73108 24388 73278
rect 24780 73332 24836 75852
rect 25452 75684 25508 75694
rect 25452 75682 26180 75684
rect 25452 75630 25454 75682
rect 25506 75630 26180 75682
rect 25452 75628 26180 75630
rect 25452 75618 25508 75628
rect 26012 75460 26068 75470
rect 25788 75458 26068 75460
rect 25788 75406 26014 75458
rect 26066 75406 26068 75458
rect 25788 75404 26068 75406
rect 25228 75010 25284 75022
rect 25228 74958 25230 75010
rect 25282 74958 25284 75010
rect 25228 74228 25284 74958
rect 25228 74162 25284 74172
rect 25452 74900 25508 74910
rect 25788 74900 25844 75404
rect 26012 75394 26068 75404
rect 25452 74898 25844 74900
rect 25452 74846 25454 74898
rect 25506 74846 25844 74898
rect 25452 74844 25844 74846
rect 26012 74900 26068 74910
rect 25452 73948 25508 74844
rect 26012 74806 26068 74844
rect 26012 74228 26068 74238
rect 26124 74228 26180 75628
rect 26684 74786 26740 74798
rect 26684 74734 26686 74786
rect 26738 74734 26740 74786
rect 26012 74226 26180 74228
rect 26012 74174 26014 74226
rect 26066 74174 26180 74226
rect 26012 74172 26180 74174
rect 26348 74340 26404 74350
rect 26012 74162 26068 74172
rect 24780 73266 24836 73276
rect 25228 73892 25508 73948
rect 26348 74002 26404 74284
rect 26572 74116 26628 74126
rect 26348 73950 26350 74002
rect 26402 73950 26404 74002
rect 26348 73938 26404 73950
rect 26460 74114 26628 74116
rect 26460 74062 26574 74114
rect 26626 74062 26628 74114
rect 26460 74060 26628 74062
rect 24892 73108 24948 73118
rect 24332 73052 24892 73108
rect 24556 72660 24612 72670
rect 22428 70914 22484 70924
rect 22428 70420 22484 70430
rect 21420 70354 21476 70364
rect 21868 70418 22484 70420
rect 21868 70366 22430 70418
rect 22482 70366 22484 70418
rect 21868 70364 22484 70366
rect 21308 70194 21364 70206
rect 21308 70142 21310 70194
rect 21362 70142 21364 70194
rect 21308 69636 21364 70142
rect 21868 70194 21924 70364
rect 22428 70354 22484 70364
rect 21868 70142 21870 70194
rect 21922 70142 21924 70194
rect 21868 70130 21924 70142
rect 21980 70084 22036 70094
rect 21980 70082 22372 70084
rect 21980 70030 21982 70082
rect 22034 70030 22372 70082
rect 21980 70028 22372 70030
rect 21980 70018 22036 70028
rect 21308 69570 21364 69580
rect 22316 69410 22372 70028
rect 22540 69636 22596 69646
rect 22652 69636 22708 70924
rect 22988 70532 23044 71708
rect 23772 71652 23828 71662
rect 23548 71650 23828 71652
rect 23548 71598 23774 71650
rect 23826 71598 23828 71650
rect 23548 71596 23828 71598
rect 23100 71092 23156 71102
rect 23100 70998 23156 71036
rect 23548 70866 23604 71596
rect 23772 71586 23828 71596
rect 23548 70814 23550 70866
rect 23602 70814 23604 70866
rect 23548 70802 23604 70814
rect 23884 70644 23940 72268
rect 22540 69634 22708 69636
rect 22540 69582 22542 69634
rect 22594 69582 22708 69634
rect 22540 69580 22708 69582
rect 22764 70476 23044 70532
rect 23548 70588 23940 70644
rect 23996 72546 24052 72558
rect 24556 72548 24612 72604
rect 23996 72494 23998 72546
rect 24050 72494 24052 72546
rect 22764 69634 22820 70476
rect 23548 70082 23604 70588
rect 23548 70030 23550 70082
rect 23602 70030 23604 70082
rect 23548 70018 23604 70030
rect 23660 70194 23716 70206
rect 23660 70142 23662 70194
rect 23714 70142 23716 70194
rect 22764 69582 22766 69634
rect 22818 69582 22820 69634
rect 22540 69570 22596 69580
rect 22764 69570 22820 69582
rect 23436 69972 23492 69982
rect 23436 69634 23492 69916
rect 23436 69582 23438 69634
rect 23490 69582 23492 69634
rect 23436 69570 23492 69582
rect 22316 69358 22318 69410
rect 22370 69358 22372 69410
rect 22316 69346 22372 69358
rect 22988 69412 23044 69422
rect 22988 69410 23380 69412
rect 22988 69358 22990 69410
rect 23042 69358 23380 69410
rect 22988 69356 23380 69358
rect 22988 69346 23044 69356
rect 23324 68740 23380 69356
rect 23436 68740 23492 68750
rect 23324 68738 23492 68740
rect 23324 68686 23438 68738
rect 23490 68686 23492 68738
rect 23324 68684 23492 68686
rect 23436 68674 23492 68684
rect 23660 67508 23716 70142
rect 23660 67442 23716 67452
rect 23884 68626 23940 68638
rect 23884 68574 23886 68626
rect 23938 68574 23940 68626
rect 21308 67172 21364 67182
rect 21308 65490 21364 67116
rect 23324 67172 23380 67182
rect 23324 67078 23380 67116
rect 22988 66946 23044 66958
rect 22988 66894 22990 66946
rect 23042 66894 23044 66946
rect 21644 66276 21700 66286
rect 21308 65438 21310 65490
rect 21362 65438 21364 65490
rect 21308 65426 21364 65438
rect 21532 66274 21700 66276
rect 21532 66222 21646 66274
rect 21698 66222 21700 66274
rect 21532 66220 21700 66222
rect 21308 65156 21364 65166
rect 21308 64706 21364 65100
rect 21308 64654 21310 64706
rect 21362 64654 21364 64706
rect 21308 64642 21364 64654
rect 21532 62916 21588 66220
rect 21644 66210 21700 66220
rect 21756 66164 21812 66174
rect 21644 64706 21700 64718
rect 21644 64654 21646 64706
rect 21698 64654 21700 64706
rect 21644 63252 21700 64654
rect 21756 64482 21812 66108
rect 22428 66164 22484 66174
rect 22428 66070 22484 66108
rect 22092 65492 22148 65502
rect 22092 65398 22148 65436
rect 22988 65380 23044 66894
rect 22988 64820 23044 65324
rect 22652 64764 23044 64820
rect 22092 64708 22148 64718
rect 22092 64614 22148 64652
rect 21868 64596 21924 64606
rect 21868 64502 21924 64540
rect 21756 64430 21758 64482
rect 21810 64430 21812 64482
rect 21756 64418 21812 64430
rect 22652 63700 22708 64764
rect 23660 64484 23716 64494
rect 22764 64092 23268 64148
rect 22764 63922 22820 64092
rect 22764 63870 22766 63922
rect 22818 63870 22820 63922
rect 22764 63858 22820 63870
rect 23212 63922 23268 64092
rect 23212 63870 23214 63922
rect 23266 63870 23268 63922
rect 22652 63644 23044 63700
rect 21644 63186 21700 63196
rect 21532 62850 21588 62860
rect 21868 62356 21924 62366
rect 20300 62178 20356 62188
rect 20412 62132 20580 62188
rect 20860 62132 21252 62188
rect 21756 62354 21924 62356
rect 21756 62302 21870 62354
rect 21922 62302 21924 62354
rect 21756 62300 21924 62302
rect 18956 61572 19012 61582
rect 18956 61478 19012 61516
rect 18844 61282 18900 61292
rect 19180 61458 19236 61470
rect 19180 61406 19182 61458
rect 19234 61406 19236 61458
rect 19180 61236 19236 61406
rect 19516 61460 19572 61470
rect 19740 61460 19796 61470
rect 19516 61366 19572 61404
rect 19628 61458 19796 61460
rect 19628 61406 19742 61458
rect 19794 61406 19796 61458
rect 19628 61404 19796 61406
rect 19292 61348 19348 61358
rect 19292 61254 19348 61292
rect 19180 61170 19236 61180
rect 19516 61236 19572 61246
rect 19628 61236 19684 61404
rect 19740 61394 19796 61404
rect 19852 61458 19908 62132
rect 20076 61572 20132 61582
rect 20076 61570 20356 61572
rect 20076 61518 20078 61570
rect 20130 61518 20356 61570
rect 20076 61516 20356 61518
rect 20076 61506 20132 61516
rect 19852 61406 19854 61458
rect 19906 61406 19908 61458
rect 19852 61394 19908 61406
rect 19572 61180 19684 61236
rect 20188 61346 20244 61358
rect 20188 61294 20190 61346
rect 20242 61294 20244 61346
rect 19836 61180 20100 61190
rect 19516 61170 19572 61180
rect 18732 60498 18788 60508
rect 19068 61124 19124 61134
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 18508 58604 18676 58660
rect 18956 58772 19012 58782
rect 18284 57596 18452 57652
rect 17724 57372 18004 57428
rect 17612 56082 17780 56084
rect 17612 56030 17614 56082
rect 17666 56030 17780 56082
rect 17612 56028 17780 56030
rect 17612 56018 17668 56028
rect 17500 55858 17556 55870
rect 17500 55806 17502 55858
rect 17554 55806 17556 55858
rect 17500 55186 17556 55806
rect 17500 55134 17502 55186
rect 17554 55134 17556 55186
rect 17500 55122 17556 55134
rect 17612 54628 17668 54638
rect 17612 54534 17668 54572
rect 17724 54516 17780 56028
rect 17948 55636 18004 57372
rect 18284 57426 18340 57438
rect 18284 57374 18286 57426
rect 18338 57374 18340 57426
rect 17948 55570 18004 55580
rect 18172 56196 18228 56206
rect 17948 54740 18004 54750
rect 17948 54646 18004 54684
rect 18172 54738 18228 56140
rect 18284 55972 18340 57374
rect 18396 56196 18452 57596
rect 18508 56980 18564 58604
rect 18844 58546 18900 58558
rect 18844 58494 18846 58546
rect 18898 58494 18900 58546
rect 18620 58436 18676 58446
rect 18676 58380 18788 58436
rect 18620 58370 18676 58380
rect 18620 58210 18676 58222
rect 18620 58158 18622 58210
rect 18674 58158 18676 58210
rect 18620 57652 18676 58158
rect 18732 57874 18788 58380
rect 18732 57822 18734 57874
rect 18786 57822 18788 57874
rect 18732 57810 18788 57822
rect 18620 57596 18788 57652
rect 18508 56914 18564 56924
rect 18620 57426 18676 57438
rect 18620 57374 18622 57426
rect 18674 57374 18676 57426
rect 18396 56140 18564 56196
rect 18396 55972 18452 55982
rect 18284 55970 18452 55972
rect 18284 55918 18398 55970
rect 18450 55918 18452 55970
rect 18284 55916 18452 55918
rect 18396 55860 18452 55916
rect 18396 55794 18452 55804
rect 18172 54686 18174 54738
rect 18226 54686 18228 54738
rect 18172 54674 18228 54686
rect 18396 55300 18452 55310
rect 17836 54516 17892 54526
rect 17724 54514 17892 54516
rect 17724 54462 17838 54514
rect 17890 54462 17892 54514
rect 17724 54460 17892 54462
rect 17388 54348 17668 54404
rect 17164 54124 17556 54180
rect 16268 53676 16548 53732
rect 16604 53676 16884 53732
rect 16268 53620 16324 53676
rect 16268 53526 16324 53564
rect 16380 53508 16436 53518
rect 16492 53508 16548 53676
rect 16716 53508 16772 53518
rect 16492 53506 16772 53508
rect 16492 53454 16718 53506
rect 16770 53454 16772 53506
rect 16492 53452 16772 53454
rect 16380 53170 16436 53452
rect 16716 53442 16772 53452
rect 16380 53118 16382 53170
rect 16434 53118 16436 53170
rect 16380 53106 16436 53118
rect 16268 53060 16324 53070
rect 15820 52894 15822 52946
rect 15874 52894 15876 52946
rect 15596 52222 15598 52274
rect 15650 52222 15652 52274
rect 15596 52210 15652 52222
rect 15820 51380 15876 52894
rect 15708 51324 15876 51380
rect 15932 53058 16324 53060
rect 15932 53006 16270 53058
rect 16322 53006 16324 53058
rect 15932 53004 16324 53006
rect 15596 49812 15652 49822
rect 15708 49812 15764 51324
rect 15932 50148 15988 53004
rect 16268 52994 16324 53004
rect 16604 52948 16660 52958
rect 16604 52854 16660 52892
rect 16604 52612 16660 52622
rect 15820 50036 15876 50046
rect 15932 50036 15988 50092
rect 15820 50034 15988 50036
rect 15820 49982 15822 50034
rect 15874 49982 15988 50034
rect 15820 49980 15988 49982
rect 16156 52276 16212 52286
rect 15820 49970 15876 49980
rect 15708 49756 15876 49812
rect 15596 49718 15652 49756
rect 15484 46834 15540 46844
rect 15596 49364 15652 49374
rect 15092 45836 15204 45892
rect 15372 45890 15428 45902
rect 15596 45892 15652 49308
rect 15708 49028 15764 49038
rect 15708 48934 15764 48972
rect 15820 48804 15876 49756
rect 16156 49700 16212 52220
rect 16380 50148 16436 50158
rect 16380 49978 16436 50092
rect 16268 49922 16324 49934
rect 16268 49870 16270 49922
rect 16322 49870 16324 49922
rect 16380 49926 16382 49978
rect 16434 49926 16436 49978
rect 16380 49914 16436 49926
rect 16268 49812 16324 49870
rect 16268 49756 16436 49812
rect 15820 48738 15876 48748
rect 16044 49140 16100 49150
rect 15372 45838 15374 45890
rect 15426 45838 15428 45890
rect 15036 45826 15092 45836
rect 15148 45666 15204 45678
rect 15148 45614 15150 45666
rect 15202 45614 15204 45666
rect 15148 45332 15204 45614
rect 15148 45266 15204 45276
rect 15260 45444 15316 45454
rect 15260 45330 15316 45388
rect 15260 45278 15262 45330
rect 15314 45278 15316 45330
rect 15260 45266 15316 45278
rect 15372 45330 15428 45838
rect 15372 45278 15374 45330
rect 15426 45278 15428 45330
rect 15372 45266 15428 45278
rect 15484 45836 15652 45892
rect 15708 47012 15764 47022
rect 15708 46228 15764 46956
rect 15932 46900 15988 46910
rect 15260 44098 15316 44110
rect 15260 44046 15262 44098
rect 15314 44046 15316 44098
rect 15036 43988 15092 43998
rect 15036 42866 15092 43932
rect 15260 43540 15316 44046
rect 15372 43764 15428 43774
rect 15372 43650 15428 43708
rect 15372 43598 15374 43650
rect 15426 43598 15428 43650
rect 15372 43586 15428 43598
rect 15484 43652 15540 45836
rect 15596 45668 15652 45678
rect 15596 45574 15652 45612
rect 15708 45444 15764 46172
rect 15820 46452 15876 46462
rect 15820 45890 15876 46396
rect 15820 45838 15822 45890
rect 15874 45838 15876 45890
rect 15820 45826 15876 45838
rect 15932 46004 15988 46844
rect 15932 45890 15988 45948
rect 15932 45838 15934 45890
rect 15986 45838 15988 45890
rect 15932 45826 15988 45838
rect 16044 45556 16100 49084
rect 16156 49026 16212 49644
rect 16268 49588 16324 49598
rect 16268 49494 16324 49532
rect 16156 48974 16158 49026
rect 16210 48974 16212 49026
rect 16156 48962 16212 48974
rect 16268 48916 16324 48926
rect 16380 48916 16436 49756
rect 16324 48860 16436 48916
rect 16156 48804 16212 48814
rect 16156 45668 16212 48748
rect 16268 48130 16324 48860
rect 16268 48078 16270 48130
rect 16322 48078 16324 48130
rect 16268 48066 16324 48078
rect 16604 46116 16660 52556
rect 16828 52276 16884 53676
rect 16492 46060 16660 46116
rect 16716 52220 16884 52276
rect 16380 45668 16436 45678
rect 16156 45666 16436 45668
rect 16156 45614 16382 45666
rect 16434 45614 16436 45666
rect 16156 45612 16436 45614
rect 16044 45500 16324 45556
rect 15596 45332 15652 45342
rect 15708 45332 15764 45388
rect 15596 45330 15764 45332
rect 15596 45278 15598 45330
rect 15650 45278 15764 45330
rect 15596 45276 15764 45278
rect 15596 45266 15652 45276
rect 15708 45108 15764 45118
rect 15708 45014 15764 45052
rect 15932 44436 15988 44446
rect 16268 44436 16324 45500
rect 16380 44996 16436 45612
rect 16492 45108 16548 46060
rect 16604 45890 16660 45902
rect 16604 45838 16606 45890
rect 16658 45838 16660 45890
rect 16604 45780 16660 45838
rect 16604 45714 16660 45724
rect 16716 45332 16772 52220
rect 17052 50708 17108 50718
rect 17052 49026 17108 50652
rect 17052 48974 17054 49026
rect 17106 48974 17108 49026
rect 17052 48962 17108 48974
rect 17500 47348 17556 54124
rect 17612 50036 17668 54348
rect 17724 53508 17780 53518
rect 17724 52274 17780 53452
rect 17836 53172 17892 54460
rect 18396 54516 18452 55244
rect 18508 55076 18564 56140
rect 18620 55298 18676 57374
rect 18732 57428 18788 57596
rect 18732 57362 18788 57372
rect 18844 56866 18900 58494
rect 18956 58322 19012 58716
rect 18956 58270 18958 58322
rect 19010 58270 19012 58322
rect 18956 58258 19012 58270
rect 18844 56814 18846 56866
rect 18898 56814 18900 56866
rect 18844 56802 18900 56814
rect 18956 57428 19012 57438
rect 18956 56644 19012 57372
rect 19068 56868 19124 61068
rect 19180 60676 19236 60686
rect 19180 60582 19236 60620
rect 19964 60676 20020 60686
rect 20020 60620 20132 60676
rect 19964 60610 20020 60620
rect 19292 60116 19348 60126
rect 19180 58322 19236 58334
rect 19180 58270 19182 58322
rect 19234 58270 19236 58322
rect 19180 57426 19236 58270
rect 19180 57374 19182 57426
rect 19234 57374 19236 57426
rect 19180 57362 19236 57374
rect 19292 57204 19348 60060
rect 20076 60114 20132 60620
rect 20076 60062 20078 60114
rect 20130 60062 20132 60114
rect 20076 60050 20132 60062
rect 19852 60004 19908 60014
rect 19852 59910 19908 59948
rect 20188 60002 20244 61294
rect 20188 59950 20190 60002
rect 20242 59950 20244 60002
rect 20188 59938 20244 59950
rect 20300 60004 20356 61516
rect 20300 59938 20356 59948
rect 20412 61346 20468 62132
rect 20412 61294 20414 61346
rect 20466 61294 20468 61346
rect 20412 60676 20468 61294
rect 20524 61458 20580 61470
rect 20524 61406 20526 61458
rect 20578 61406 20580 61458
rect 20524 61348 20580 61406
rect 20524 61012 20580 61292
rect 20524 60946 20580 60956
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19628 59220 19684 59230
rect 19628 59126 19684 59164
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19964 57652 20020 57662
rect 19964 57558 20020 57596
rect 20188 57652 20244 57662
rect 20412 57652 20468 60620
rect 20524 59892 20580 59902
rect 20524 59798 20580 59836
rect 20636 59218 20692 59230
rect 20636 59166 20638 59218
rect 20690 59166 20692 59218
rect 20636 59108 20692 59166
rect 20636 59042 20692 59052
rect 20188 57650 20468 57652
rect 20188 57598 20190 57650
rect 20242 57598 20468 57650
rect 20188 57596 20468 57598
rect 20524 58212 20580 58222
rect 20524 57650 20580 58156
rect 20636 57764 20692 57774
rect 20636 57762 20804 57764
rect 20636 57710 20638 57762
rect 20690 57710 20804 57762
rect 20636 57708 20804 57710
rect 20636 57698 20692 57708
rect 20524 57598 20526 57650
rect 20578 57598 20580 57650
rect 20188 57586 20244 57596
rect 19404 57538 19460 57550
rect 19404 57486 19406 57538
rect 19458 57486 19460 57538
rect 19404 57428 19460 57486
rect 19404 57362 19460 57372
rect 19516 57426 19572 57438
rect 19516 57374 19518 57426
rect 19570 57374 19572 57426
rect 19292 57148 19460 57204
rect 19292 56868 19348 56878
rect 19068 56866 19348 56868
rect 19068 56814 19294 56866
rect 19346 56814 19348 56866
rect 19068 56812 19348 56814
rect 19292 56802 19348 56812
rect 18844 56588 19012 56644
rect 19180 56642 19236 56654
rect 19180 56590 19182 56642
rect 19234 56590 19236 56642
rect 18732 55860 18788 55870
rect 18844 55860 18900 56588
rect 18956 56420 19012 56430
rect 18956 56306 19012 56364
rect 18956 56254 18958 56306
rect 19010 56254 19012 56306
rect 18956 56242 19012 56254
rect 18788 55804 18900 55860
rect 19068 55860 19124 55870
rect 18732 55766 18788 55804
rect 19068 55766 19124 55804
rect 19180 55636 19236 56590
rect 19180 55570 19236 55580
rect 18620 55246 18622 55298
rect 18674 55246 18676 55298
rect 18620 55234 18676 55246
rect 19292 55300 19348 55310
rect 19404 55300 19460 57148
rect 19292 55298 19460 55300
rect 19292 55246 19294 55298
rect 19346 55246 19460 55298
rect 19292 55244 19460 55246
rect 19516 56980 19572 57374
rect 19852 57426 19908 57438
rect 19852 57374 19854 57426
rect 19906 57374 19908 57426
rect 19852 57092 19908 57374
rect 20188 57204 20244 57214
rect 19852 56980 19908 57036
rect 19516 56924 19908 56980
rect 20076 57148 20188 57204
rect 19292 55234 19348 55244
rect 18508 55020 19124 55076
rect 18620 54626 18676 54638
rect 18620 54574 18622 54626
rect 18674 54574 18676 54626
rect 18508 54516 18564 54526
rect 18396 54514 18564 54516
rect 18396 54462 18510 54514
rect 18562 54462 18564 54514
rect 18396 54460 18564 54462
rect 18284 53172 18340 53182
rect 17836 53170 18340 53172
rect 17836 53118 18286 53170
rect 18338 53118 18340 53170
rect 17836 53116 18340 53118
rect 18284 53106 18340 53116
rect 18396 52948 18452 54460
rect 18508 54450 18564 54460
rect 18620 53954 18676 54574
rect 18620 53902 18622 53954
rect 18674 53902 18676 53954
rect 18620 53890 18676 53902
rect 18732 53618 18788 53630
rect 18732 53566 18734 53618
rect 18786 53566 18788 53618
rect 18620 53508 18676 53518
rect 18620 53414 18676 53452
rect 18732 53060 18788 53566
rect 18620 53004 18788 53060
rect 17724 52222 17726 52274
rect 17778 52222 17780 52274
rect 17724 52210 17780 52222
rect 18284 52892 18452 52948
rect 18508 52948 18564 52958
rect 17836 51716 17892 51726
rect 17724 51660 17836 51716
rect 17724 50428 17780 51660
rect 17836 51650 17892 51660
rect 18172 50708 18228 50718
rect 18284 50708 18340 52892
rect 18508 52854 18564 52892
rect 18172 50706 18340 50708
rect 18172 50654 18174 50706
rect 18226 50654 18340 50706
rect 18172 50652 18340 50654
rect 18396 52500 18452 52510
rect 18172 50642 18228 50652
rect 17724 50372 17892 50428
rect 17612 49970 17668 49980
rect 17836 50034 17892 50372
rect 17836 49982 17838 50034
rect 17890 49982 17892 50034
rect 17836 49812 17892 49982
rect 17948 50036 18004 50046
rect 17948 49942 18004 49980
rect 18396 49812 18452 52444
rect 18620 50932 18676 53004
rect 18956 52948 19012 52958
rect 18732 52946 19012 52948
rect 18732 52894 18958 52946
rect 19010 52894 19012 52946
rect 18732 52892 19012 52894
rect 18732 51716 18788 52892
rect 18956 52882 19012 52892
rect 19068 52724 19124 55020
rect 19180 55074 19236 55086
rect 19180 55022 19182 55074
rect 19234 55022 19236 55074
rect 19180 53956 19236 55022
rect 19180 53890 19236 53900
rect 19292 53172 19348 53182
rect 19516 53172 19572 56924
rect 20076 56868 20132 57148
rect 20188 57138 20244 57148
rect 19628 56866 20132 56868
rect 19628 56814 20078 56866
rect 20130 56814 20132 56866
rect 19628 56812 20132 56814
rect 19628 55972 19684 56812
rect 20076 56802 20132 56812
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20188 56084 20244 56094
rect 20188 56082 20356 56084
rect 20188 56030 20190 56082
rect 20242 56030 20356 56082
rect 20188 56028 20356 56030
rect 20188 56018 20244 56028
rect 19628 55970 20132 55972
rect 19628 55918 19630 55970
rect 19682 55918 20132 55970
rect 19628 55916 20132 55918
rect 19628 55906 19684 55916
rect 20076 55298 20132 55916
rect 20076 55246 20078 55298
rect 20130 55246 20132 55298
rect 20076 55076 20132 55246
rect 20076 55010 20132 55020
rect 20188 55860 20244 55870
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54514 20244 55804
rect 20300 55412 20356 56028
rect 20524 56082 20580 57598
rect 20636 56196 20692 56206
rect 20636 56102 20692 56140
rect 20524 56030 20526 56082
rect 20578 56030 20580 56082
rect 20412 55412 20468 55422
rect 20300 55356 20412 55412
rect 20412 55346 20468 55356
rect 20188 54462 20190 54514
rect 20242 54462 20244 54514
rect 20188 54450 20244 54462
rect 20300 55188 20356 55198
rect 20188 54292 20244 54302
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19292 53170 19572 53172
rect 19292 53118 19294 53170
rect 19346 53118 19572 53170
rect 19292 53116 19572 53118
rect 19292 53106 19348 53116
rect 19852 52948 19908 52958
rect 18844 52668 19124 52724
rect 19180 52836 19236 52846
rect 18844 52386 18900 52668
rect 18844 52334 18846 52386
rect 18898 52334 18900 52386
rect 18844 52322 18900 52334
rect 19068 52164 19124 52174
rect 18844 52052 18900 52062
rect 18844 51958 18900 51996
rect 18956 52050 19012 52062
rect 18956 51998 18958 52050
rect 19010 51998 19012 52050
rect 18956 51828 19012 51998
rect 18956 51762 19012 51772
rect 18732 51650 18788 51660
rect 18956 51268 19012 51278
rect 18620 50866 18676 50876
rect 18844 51266 19012 51268
rect 18844 51214 18958 51266
rect 19010 51214 19012 51266
rect 18844 51212 19012 51214
rect 18508 50596 18564 50606
rect 18508 50034 18564 50540
rect 18508 49982 18510 50034
rect 18562 49982 18564 50034
rect 18508 49970 18564 49982
rect 18620 50372 18676 50382
rect 18844 50372 18900 51212
rect 18956 51202 19012 51212
rect 18620 50370 18900 50372
rect 18620 50318 18622 50370
rect 18674 50318 18900 50370
rect 18620 50316 18900 50318
rect 18956 51044 19012 51054
rect 17836 49756 18228 49812
rect 18396 49756 18564 49812
rect 18060 49586 18116 49598
rect 18060 49534 18062 49586
rect 18114 49534 18116 49586
rect 17724 49364 17780 49374
rect 18060 49364 18116 49534
rect 17724 49026 17780 49308
rect 17724 48974 17726 49026
rect 17778 48974 17780 49026
rect 17724 47572 17780 48974
rect 17724 47506 17780 47516
rect 17836 49308 18116 49364
rect 17836 48354 17892 49308
rect 17836 48302 17838 48354
rect 17890 48302 17892 48354
rect 17500 47292 17668 47348
rect 17500 46900 17556 46910
rect 17500 46806 17556 46844
rect 17388 46676 17444 46686
rect 16716 45266 16772 45276
rect 17052 46674 17444 46676
rect 17052 46622 17390 46674
rect 17442 46622 17444 46674
rect 17052 46620 17444 46622
rect 16716 45108 16772 45118
rect 16492 45052 16660 45108
rect 16380 44940 16548 44996
rect 15932 44434 16324 44436
rect 15932 44382 15934 44434
rect 15986 44382 16324 44434
rect 15932 44380 16324 44382
rect 15932 44370 15988 44380
rect 16268 44210 16324 44380
rect 16268 44158 16270 44210
rect 16322 44158 16324 44210
rect 16268 44146 16324 44158
rect 16380 44324 16436 44334
rect 16044 44098 16100 44110
rect 16044 44046 16046 44098
rect 16098 44046 16100 44098
rect 15596 43652 15652 43662
rect 16044 43652 16100 44046
rect 16380 43876 16436 44268
rect 15484 43650 15652 43652
rect 15484 43598 15598 43650
rect 15650 43598 15652 43650
rect 15484 43596 15652 43598
rect 15260 43474 15316 43484
rect 15036 42814 15038 42866
rect 15090 42814 15092 42866
rect 15036 42802 15092 42814
rect 15596 42868 15652 43596
rect 15932 43596 16100 43652
rect 16156 43820 16436 43876
rect 15932 43538 15988 43596
rect 15932 43486 15934 43538
rect 15986 43486 15988 43538
rect 15932 43474 15988 43486
rect 15036 42308 15092 42318
rect 15484 42308 15540 42318
rect 15036 41298 15092 42252
rect 15036 41246 15038 41298
rect 15090 41246 15092 41298
rect 15036 40964 15092 41246
rect 15372 42252 15484 42308
rect 15372 41186 15428 42252
rect 15484 42242 15540 42252
rect 15596 41860 15652 42812
rect 16044 43426 16100 43438
rect 16044 43374 16046 43426
rect 16098 43374 16100 43426
rect 15932 42420 15988 42430
rect 15932 41860 15988 42364
rect 16044 42084 16100 43374
rect 16044 42018 16100 42028
rect 16044 41860 16100 41870
rect 15932 41858 16100 41860
rect 15932 41806 16046 41858
rect 16098 41806 16100 41858
rect 15932 41804 16100 41806
rect 15596 41794 15652 41804
rect 16044 41794 16100 41804
rect 15372 41134 15374 41186
rect 15426 41134 15428 41186
rect 15372 41122 15428 41134
rect 15708 41076 15764 41086
rect 15932 41076 15988 41086
rect 15708 41074 15988 41076
rect 15708 41022 15710 41074
rect 15762 41022 15934 41074
rect 15986 41022 15988 41074
rect 15708 41020 15988 41022
rect 15708 41010 15764 41020
rect 15932 41010 15988 41020
rect 15484 40964 15540 40974
rect 15036 40908 15484 40964
rect 15484 40870 15540 40908
rect 16044 40962 16100 40974
rect 16044 40910 16046 40962
rect 16098 40910 16100 40962
rect 14924 38546 14980 38556
rect 15036 40290 15092 40302
rect 15036 40238 15038 40290
rect 15090 40238 15092 40290
rect 14700 37998 14702 38050
rect 14754 37998 14756 38050
rect 14700 37986 14756 37998
rect 15036 37380 15092 40238
rect 15484 38948 15540 38958
rect 15484 38854 15540 38892
rect 15820 38946 15876 38958
rect 15820 38894 15822 38946
rect 15874 38894 15876 38946
rect 15820 38836 15876 38894
rect 15820 38770 15876 38780
rect 16044 38668 16100 40910
rect 16156 40180 16212 43820
rect 16380 43652 16436 43662
rect 16268 43650 16436 43652
rect 16268 43598 16382 43650
rect 16434 43598 16436 43650
rect 16268 43596 16436 43598
rect 16268 43538 16324 43596
rect 16380 43586 16436 43596
rect 16268 43486 16270 43538
rect 16322 43486 16324 43538
rect 16268 43474 16324 43486
rect 16492 43316 16548 44940
rect 16604 44548 16660 45052
rect 16604 43764 16660 44492
rect 16604 43650 16660 43708
rect 16604 43598 16606 43650
rect 16658 43598 16660 43650
rect 16604 43586 16660 43598
rect 16716 43650 16772 45052
rect 16828 44322 16884 44334
rect 16828 44270 16830 44322
rect 16882 44270 16884 44322
rect 16828 44212 16884 44270
rect 16828 44146 16884 44156
rect 17052 44324 17108 46620
rect 17388 46610 17444 46620
rect 17500 46452 17556 46462
rect 17500 46358 17556 46396
rect 17500 46116 17556 46126
rect 17612 46116 17668 47292
rect 17500 46114 17668 46116
rect 17500 46062 17502 46114
rect 17554 46062 17668 46114
rect 17500 46060 17668 46062
rect 17500 46050 17556 46060
rect 17164 46004 17220 46014
rect 17164 45910 17220 45948
rect 17836 45892 17892 48302
rect 17948 48356 18004 48366
rect 17948 48262 18004 48300
rect 18060 48020 18116 48030
rect 18060 47926 18116 47964
rect 18060 46900 18116 46910
rect 18172 46900 18228 49756
rect 18396 49252 18452 49262
rect 18396 49138 18452 49196
rect 18396 49086 18398 49138
rect 18450 49086 18452 49138
rect 18396 49074 18452 49086
rect 18060 46898 18452 46900
rect 18060 46846 18062 46898
rect 18114 46846 18452 46898
rect 18060 46844 18452 46846
rect 18060 46834 18116 46844
rect 18284 46674 18340 46686
rect 18284 46622 18286 46674
rect 18338 46622 18340 46674
rect 17836 45890 18004 45892
rect 17836 45838 17838 45890
rect 17890 45838 18004 45890
rect 17836 45836 18004 45838
rect 17836 45826 17892 45836
rect 17836 45332 17892 45342
rect 17500 45108 17556 45118
rect 17500 45014 17556 45052
rect 17836 45106 17892 45276
rect 17836 45054 17838 45106
rect 17890 45054 17892 45106
rect 17836 45042 17892 45054
rect 17724 44994 17780 45006
rect 17724 44942 17726 44994
rect 17778 44942 17780 44994
rect 17724 44324 17780 44942
rect 17836 44324 17892 44334
rect 17724 44268 17836 44324
rect 17052 44210 17108 44268
rect 17836 44230 17892 44268
rect 17052 44158 17054 44210
rect 17106 44158 17108 44210
rect 17052 44146 17108 44158
rect 17500 44212 17556 44222
rect 17500 44098 17556 44156
rect 17500 44046 17502 44098
rect 17554 44046 17556 44098
rect 17500 44034 17556 44046
rect 17948 43764 18004 45836
rect 18060 45780 18116 45790
rect 18284 45780 18340 46622
rect 18060 45778 18340 45780
rect 18060 45726 18062 45778
rect 18114 45726 18340 45778
rect 18060 45724 18340 45726
rect 18060 44884 18116 45724
rect 18396 45332 18452 46844
rect 18508 46114 18564 49756
rect 18620 49364 18676 50316
rect 18844 50036 18900 50046
rect 18844 49942 18900 49980
rect 18620 49298 18676 49308
rect 18620 49028 18676 49038
rect 18620 48934 18676 48972
rect 18620 48132 18676 48142
rect 18620 48038 18676 48076
rect 18956 47068 19012 50988
rect 19068 50596 19124 52108
rect 19180 52162 19236 52780
rect 19180 52110 19182 52162
rect 19234 52110 19236 52162
rect 19180 52098 19236 52110
rect 19852 52164 19908 52892
rect 19852 52070 19908 52108
rect 19516 52050 19572 52062
rect 19516 51998 19518 52050
rect 19570 51998 19572 52050
rect 19404 51940 19460 51950
rect 19404 51846 19460 51884
rect 19516 51828 19572 51998
rect 19068 50530 19124 50540
rect 19404 50596 19460 50606
rect 19404 50034 19460 50540
rect 19404 49982 19406 50034
rect 19458 49982 19460 50034
rect 19404 49970 19460 49982
rect 19180 49812 19236 49822
rect 19516 49812 19572 51772
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20076 50932 20132 50942
rect 20076 50706 20132 50876
rect 20076 50654 20078 50706
rect 20130 50654 20132 50706
rect 20076 50642 20132 50654
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19180 49810 19572 49812
rect 19180 49758 19182 49810
rect 19234 49758 19572 49810
rect 19180 49756 19572 49758
rect 19628 49922 19684 49934
rect 19628 49870 19630 49922
rect 19682 49870 19684 49922
rect 19068 49588 19124 49598
rect 19068 49026 19124 49532
rect 19068 48974 19070 49026
rect 19122 48974 19124 49026
rect 19068 48962 19124 48974
rect 18508 46062 18510 46114
rect 18562 46062 18564 46114
rect 18508 46050 18564 46062
rect 18844 47012 19012 47068
rect 18620 45890 18676 45902
rect 18620 45838 18622 45890
rect 18674 45838 18676 45890
rect 18620 45556 18676 45838
rect 18620 45500 18788 45556
rect 18620 45332 18676 45342
rect 18452 45330 18676 45332
rect 18452 45278 18622 45330
rect 18674 45278 18676 45330
rect 18452 45276 18676 45278
rect 18396 45238 18452 45276
rect 18620 45266 18676 45276
rect 18060 44434 18116 44828
rect 18060 44382 18062 44434
rect 18114 44382 18116 44434
rect 18060 44370 18116 44382
rect 18732 44324 18788 45500
rect 18844 45220 18900 47012
rect 19068 46900 19124 46910
rect 18956 46564 19012 46574
rect 19068 46564 19124 46844
rect 18956 46562 19124 46564
rect 18956 46510 18958 46562
rect 19010 46510 19124 46562
rect 18956 46508 19124 46510
rect 18956 46498 19012 46508
rect 18956 45890 19012 45902
rect 18956 45838 18958 45890
rect 19010 45838 19012 45890
rect 18956 45668 19012 45838
rect 18956 45602 19012 45612
rect 18956 45220 19012 45230
rect 18844 45218 19012 45220
rect 18844 45166 18958 45218
rect 19010 45166 19012 45218
rect 18844 45164 19012 45166
rect 18732 44258 18788 44268
rect 18956 43876 19012 45164
rect 19180 44994 19236 49756
rect 19628 49364 19684 49870
rect 19740 49812 19796 49822
rect 19740 49718 19796 49756
rect 19628 49298 19684 49308
rect 19404 49028 19460 49038
rect 19404 45332 19460 48972
rect 20188 49028 20244 54236
rect 20300 52612 20356 55132
rect 20524 53732 20580 56030
rect 20524 53666 20580 53676
rect 20748 53396 20804 57708
rect 20748 53330 20804 53340
rect 20524 53172 20580 53182
rect 20748 53172 20804 53182
rect 20580 53170 20804 53172
rect 20580 53118 20750 53170
rect 20802 53118 20804 53170
rect 20580 53116 20804 53118
rect 20524 53106 20580 53116
rect 20748 53106 20804 53116
rect 20636 52948 20692 52958
rect 20300 52546 20356 52556
rect 20412 52946 20692 52948
rect 20412 52894 20638 52946
rect 20690 52894 20692 52946
rect 20412 52892 20692 52894
rect 20412 52050 20468 52892
rect 20636 52882 20692 52892
rect 20748 52948 20804 52958
rect 20860 52948 20916 62132
rect 20972 61684 21028 61694
rect 20972 54292 21028 61628
rect 21644 61570 21700 61582
rect 21644 61518 21646 61570
rect 21698 61518 21700 61570
rect 21644 61460 21700 61518
rect 21644 61394 21700 61404
rect 21756 60788 21812 62300
rect 21868 62290 21924 62300
rect 22540 62242 22596 62254
rect 22540 62190 22542 62242
rect 22594 62190 22596 62242
rect 22540 62188 22596 62190
rect 21868 62132 22596 62188
rect 22876 62244 22932 62254
rect 21868 61682 21924 62132
rect 22764 61794 22820 61806
rect 22764 61742 22766 61794
rect 22818 61742 22820 61794
rect 22764 61684 22820 61742
rect 21868 61630 21870 61682
rect 21922 61630 21924 61682
rect 21868 61618 21924 61630
rect 22204 61628 22820 61684
rect 22092 61572 22148 61582
rect 22204 61572 22260 61628
rect 22092 61570 22260 61572
rect 22092 61518 22094 61570
rect 22146 61518 22260 61570
rect 22092 61516 22260 61518
rect 22092 61506 22148 61516
rect 22316 61458 22372 61470
rect 22316 61406 22318 61458
rect 22370 61406 22372 61458
rect 22316 60900 22372 61406
rect 22652 61458 22708 61470
rect 22652 61406 22654 61458
rect 22706 61406 22708 61458
rect 22652 61348 22708 61406
rect 22540 60900 22596 60910
rect 22316 60844 22540 60900
rect 21756 60694 21812 60732
rect 21308 60676 21364 60686
rect 22428 60676 22484 60686
rect 21308 60582 21364 60620
rect 21868 60674 22484 60676
rect 21868 60622 22430 60674
rect 22482 60622 22484 60674
rect 21868 60620 22484 60622
rect 21868 60114 21924 60620
rect 22428 60610 22484 60620
rect 21868 60062 21870 60114
rect 21922 60062 21924 60114
rect 21868 60050 21924 60062
rect 22092 60116 22148 60126
rect 21644 60004 21700 60014
rect 21644 59910 21700 59948
rect 22092 60002 22148 60060
rect 22092 59950 22094 60002
rect 22146 59950 22148 60002
rect 22092 59938 22148 59950
rect 22316 59892 22372 59902
rect 22540 59892 22596 60844
rect 22372 59836 22596 59892
rect 22652 59890 22708 61292
rect 22764 61348 22820 61358
rect 22876 61348 22932 62188
rect 22764 61346 22932 61348
rect 22764 61294 22766 61346
rect 22818 61294 22932 61346
rect 22764 61292 22932 61294
rect 22764 61282 22820 61292
rect 22764 60226 22820 60238
rect 22764 60174 22766 60226
rect 22818 60174 22820 60226
rect 22764 60116 22820 60174
rect 22764 60050 22820 60060
rect 22652 59838 22654 59890
rect 22706 59838 22708 59890
rect 22316 59798 22372 59836
rect 22652 59826 22708 59838
rect 22764 59892 22820 59902
rect 21868 59444 21924 59454
rect 21868 59350 21924 59388
rect 21420 59218 21476 59230
rect 21420 59166 21422 59218
rect 21474 59166 21476 59218
rect 21420 57204 21476 59166
rect 22204 58658 22260 58670
rect 22204 58606 22206 58658
rect 22258 58606 22260 58658
rect 22204 58548 22260 58606
rect 22764 58658 22820 59836
rect 22764 58606 22766 58658
rect 22818 58606 22820 58658
rect 22764 58594 22820 58606
rect 21420 57138 21476 57148
rect 21980 58546 22260 58548
rect 21980 58494 22206 58546
rect 22258 58494 22260 58546
rect 21980 58492 22260 58494
rect 21756 57092 21812 57102
rect 21756 56998 21812 57036
rect 21980 56754 22036 58492
rect 22204 58482 22260 58492
rect 22652 58210 22708 58222
rect 22652 58158 22654 58210
rect 22706 58158 22708 58210
rect 22652 57876 22708 58158
rect 22652 57810 22708 57820
rect 22204 57652 22260 57662
rect 22204 57558 22260 57596
rect 22428 57092 22484 57102
rect 22428 56998 22484 57036
rect 21980 56702 21982 56754
rect 22034 56702 22036 56754
rect 21980 56690 22036 56702
rect 22092 56978 22148 56990
rect 22092 56926 22094 56978
rect 22146 56926 22148 56978
rect 21420 56642 21476 56654
rect 21420 56590 21422 56642
rect 21474 56590 21476 56642
rect 21420 55188 21476 56590
rect 22092 56084 22148 56926
rect 22764 56868 22820 56878
rect 22876 56868 22932 61292
rect 22764 56866 22932 56868
rect 22764 56814 22766 56866
rect 22818 56814 22932 56866
rect 22764 56812 22932 56814
rect 22764 56802 22820 56812
rect 22540 56642 22596 56654
rect 22540 56590 22542 56642
rect 22594 56590 22596 56642
rect 22204 56084 22260 56094
rect 22092 56082 22260 56084
rect 22092 56030 22206 56082
rect 22258 56030 22260 56082
rect 22092 56028 22260 56030
rect 22204 56018 22260 56028
rect 22428 55972 22484 55982
rect 21532 55412 21588 55422
rect 21532 55318 21588 55356
rect 22316 55300 22372 55310
rect 22316 55206 22372 55244
rect 21420 55122 21476 55132
rect 21980 55076 22036 55086
rect 22428 55076 22484 55916
rect 21196 54628 21252 54638
rect 21196 54514 21252 54572
rect 21196 54462 21198 54514
rect 21250 54462 21252 54514
rect 21196 54450 21252 54462
rect 21980 54514 22036 55020
rect 21980 54462 21982 54514
rect 22034 54462 22036 54514
rect 21980 54450 22036 54462
rect 22316 55020 22484 55076
rect 20972 54226 21028 54236
rect 22316 53844 22372 55020
rect 22540 54852 22596 56590
rect 22988 55300 23044 63644
rect 23212 62188 23268 63870
rect 23660 62188 23716 64428
rect 23884 62244 23940 68574
rect 23996 67172 24052 72494
rect 24444 72546 24612 72548
rect 24444 72494 24558 72546
rect 24610 72494 24612 72546
rect 24444 72492 24612 72494
rect 24332 71764 24388 71774
rect 24332 71670 24388 71708
rect 24444 70308 24500 72492
rect 24556 72482 24612 72492
rect 24332 70252 24500 70308
rect 24556 70978 24612 70990
rect 24556 70926 24558 70978
rect 24610 70926 24612 70978
rect 24556 70306 24612 70926
rect 24556 70254 24558 70306
rect 24610 70254 24612 70306
rect 24220 69188 24276 69198
rect 24220 69094 24276 69132
rect 24332 68626 24388 70252
rect 24556 70242 24612 70254
rect 24668 69188 24724 69198
rect 24668 69094 24724 69132
rect 24332 68574 24334 68626
rect 24386 68574 24388 68626
rect 24332 68066 24388 68574
rect 24332 68014 24334 68066
rect 24386 68014 24388 68066
rect 24332 68002 24388 68014
rect 24780 68066 24836 68078
rect 24780 68014 24782 68066
rect 24834 68014 24836 68066
rect 24780 67954 24836 68014
rect 24780 67902 24782 67954
rect 24834 67902 24836 67954
rect 24780 67890 24836 67902
rect 24444 67508 24500 67518
rect 24500 67452 24612 67508
rect 24444 67442 24500 67452
rect 24052 67116 24276 67172
rect 23996 67106 24052 67116
rect 24220 65378 24276 67116
rect 24556 66388 24612 67452
rect 24556 66386 24724 66388
rect 24556 66334 24558 66386
rect 24610 66334 24724 66386
rect 24556 66332 24724 66334
rect 24556 66322 24612 66332
rect 24668 65602 24724 66332
rect 24668 65550 24670 65602
rect 24722 65550 24724 65602
rect 24668 65538 24724 65550
rect 24220 65326 24222 65378
rect 24274 65326 24276 65378
rect 24220 65314 24276 65326
rect 23212 62132 23492 62188
rect 23660 62132 23828 62188
rect 23884 62178 23940 62188
rect 24556 65266 24612 65278
rect 24556 65214 24558 65266
rect 24610 65214 24612 65266
rect 24556 64596 24612 65214
rect 23324 60676 23380 60686
rect 23324 60114 23380 60620
rect 23324 60062 23326 60114
rect 23378 60062 23380 60114
rect 23324 59892 23380 60062
rect 23324 59826 23380 59836
rect 23100 59106 23156 59118
rect 23100 59054 23102 59106
rect 23154 59054 23156 59106
rect 23100 58884 23156 59054
rect 23100 58818 23156 58828
rect 23100 58324 23156 58334
rect 23156 58268 23380 58324
rect 23100 58230 23156 58268
rect 22988 55234 23044 55244
rect 23100 56980 23156 56990
rect 23324 56980 23380 58268
rect 23436 57092 23492 62132
rect 23548 59106 23604 59118
rect 23548 59054 23550 59106
rect 23602 59054 23604 59106
rect 23548 58996 23604 59054
rect 23548 58930 23604 58940
rect 23772 57762 23828 62132
rect 24444 61572 24500 61582
rect 24108 60788 24164 60798
rect 23996 59330 24052 59342
rect 23996 59278 23998 59330
rect 24050 59278 24052 59330
rect 23884 59218 23940 59230
rect 23884 59166 23886 59218
rect 23938 59166 23940 59218
rect 23884 58436 23940 59166
rect 23996 58884 24052 59278
rect 24108 59220 24164 60732
rect 24444 60676 24500 61516
rect 24556 60900 24612 64540
rect 24668 62244 24724 62282
rect 24668 62178 24724 62188
rect 24892 61572 24948 73052
rect 25116 72436 25172 72446
rect 25004 72434 25172 72436
rect 25004 72382 25118 72434
rect 25170 72382 25172 72434
rect 25004 72380 25172 72382
rect 25004 70866 25060 72380
rect 25116 72370 25172 72380
rect 25004 70814 25006 70866
rect 25058 70814 25060 70866
rect 25004 70802 25060 70814
rect 25004 70196 25060 70206
rect 25004 69522 25060 70140
rect 25004 69470 25006 69522
rect 25058 69470 25060 69522
rect 25004 69458 25060 69470
rect 25228 63588 25284 73892
rect 25452 73444 25508 73454
rect 25452 73350 25508 73388
rect 25676 73332 25732 73342
rect 25564 73330 25732 73332
rect 25564 73278 25678 73330
rect 25730 73278 25732 73330
rect 25564 73276 25732 73278
rect 25340 72324 25396 72334
rect 25340 71986 25396 72268
rect 25340 71934 25342 71986
rect 25394 71934 25396 71986
rect 25340 71922 25396 71934
rect 25452 70084 25508 70094
rect 25452 69990 25508 70028
rect 25452 68740 25508 68750
rect 25564 68740 25620 73276
rect 25676 73266 25732 73276
rect 26236 73220 26292 73230
rect 25676 72660 25732 72670
rect 25676 72566 25732 72604
rect 26236 72324 26292 73164
rect 26236 72258 26292 72268
rect 26460 71090 26516 74060
rect 26572 74050 26628 74060
rect 26684 73556 26740 74734
rect 27244 74788 27300 74798
rect 27244 74002 27300 74732
rect 28588 74788 28644 74798
rect 27244 73950 27246 74002
rect 27298 73950 27300 74002
rect 27244 73938 27300 73950
rect 27580 74002 27636 74014
rect 27580 73950 27582 74002
rect 27634 73950 27636 74002
rect 26684 73490 26740 73500
rect 26684 73218 26740 73230
rect 26684 73166 26686 73218
rect 26738 73166 26740 73218
rect 26684 73108 26740 73166
rect 26684 73042 26740 73052
rect 27580 71876 27636 73950
rect 28252 74002 28308 74014
rect 28252 73950 28254 74002
rect 28306 73950 28308 74002
rect 27692 73556 27748 73566
rect 27692 73462 27748 73500
rect 28028 73330 28084 73342
rect 28028 73278 28030 73330
rect 28082 73278 28084 73330
rect 28028 72100 28084 73278
rect 28028 72034 28084 72044
rect 28140 71876 28196 71886
rect 27580 71820 28140 71876
rect 26460 71038 26462 71090
rect 26514 71038 26516 71090
rect 26460 71026 26516 71038
rect 25900 70980 25956 70990
rect 25900 70418 25956 70924
rect 25900 70366 25902 70418
rect 25954 70366 25956 70418
rect 25900 70354 25956 70366
rect 26572 70978 26628 70990
rect 26908 70980 26964 70990
rect 26572 70926 26574 70978
rect 26626 70926 26628 70978
rect 26012 70306 26068 70318
rect 26012 70254 26014 70306
rect 26066 70254 26068 70306
rect 26012 70196 26068 70254
rect 26460 70308 26516 70318
rect 26572 70308 26628 70926
rect 26460 70306 26628 70308
rect 26460 70254 26462 70306
rect 26514 70254 26628 70306
rect 26460 70252 26628 70254
rect 26460 70242 26516 70252
rect 25452 68738 25620 68740
rect 25452 68686 25454 68738
rect 25506 68686 25620 68738
rect 25452 68684 25620 68686
rect 25676 70140 26068 70196
rect 25676 69410 25732 70140
rect 25788 69970 25844 69982
rect 25788 69918 25790 69970
rect 25842 69918 25844 69970
rect 25788 69636 25844 69918
rect 25900 69636 25956 69646
rect 25788 69580 25900 69636
rect 25900 69522 25956 69580
rect 25900 69470 25902 69522
rect 25954 69470 25956 69522
rect 25900 69458 25956 69470
rect 25676 69358 25678 69410
rect 25730 69358 25732 69410
rect 25676 69188 25732 69358
rect 26572 69410 26628 70252
rect 26572 69358 26574 69410
rect 26626 69358 26628 69410
rect 26572 69346 26628 69358
rect 26796 70924 26908 70980
rect 26796 69410 26852 70924
rect 26908 70886 26964 70924
rect 27356 70308 27412 70318
rect 27132 70194 27188 70206
rect 27132 70142 27134 70194
rect 27186 70142 27188 70194
rect 27132 69860 27188 70142
rect 27356 70194 27412 70252
rect 27356 70142 27358 70194
rect 27410 70142 27412 70194
rect 27356 70130 27412 70142
rect 27804 70308 27860 70318
rect 26796 69358 26798 69410
rect 26850 69358 26852 69410
rect 26796 69346 26852 69358
rect 27020 69804 27132 69860
rect 26684 69188 26740 69198
rect 25452 68674 25508 68684
rect 25676 68068 25732 69132
rect 26124 69186 26740 69188
rect 26124 69134 26686 69186
rect 26738 69134 26740 69186
rect 26124 69132 26740 69134
rect 26124 68626 26180 69132
rect 26124 68574 26126 68626
rect 26178 68574 26180 68626
rect 26124 68562 26180 68574
rect 25564 68012 25732 68068
rect 26236 68514 26292 68526
rect 26236 68462 26238 68514
rect 26290 68462 26292 68514
rect 25452 66948 25508 66958
rect 25452 66854 25508 66892
rect 25340 64820 25396 64830
rect 25340 64726 25396 64764
rect 25452 63922 25508 63934
rect 25452 63870 25454 63922
rect 25506 63870 25508 63922
rect 25340 63588 25396 63598
rect 25228 63532 25340 63588
rect 25340 63522 25396 63532
rect 25452 63364 25508 63870
rect 25452 63298 25508 63308
rect 25340 63028 25396 63038
rect 25340 61684 25396 62972
rect 25564 62188 25620 68012
rect 26236 67842 26292 68462
rect 26236 67790 26238 67842
rect 26290 67790 26292 67842
rect 26236 66834 26292 67790
rect 26460 67842 26516 69132
rect 26684 69122 26740 69132
rect 27020 68852 27076 69804
rect 27132 69794 27188 69804
rect 27804 69634 27860 70252
rect 27804 69582 27806 69634
rect 27858 69582 27860 69634
rect 27804 69570 27860 69582
rect 28028 69860 28084 69870
rect 28028 69522 28084 69804
rect 28028 69470 28030 69522
rect 28082 69470 28084 69522
rect 28028 69458 28084 69470
rect 27132 69300 27188 69310
rect 27468 69300 27524 69310
rect 27132 69298 27524 69300
rect 27132 69246 27134 69298
rect 27186 69246 27470 69298
rect 27522 69246 27524 69298
rect 27132 69244 27524 69246
rect 27132 69234 27188 69244
rect 27468 69234 27524 69244
rect 27132 68852 27188 68862
rect 27020 68850 27188 68852
rect 27020 68798 27134 68850
rect 27186 68798 27188 68850
rect 27020 68796 27188 68798
rect 26460 67790 26462 67842
rect 26514 67790 26516 67842
rect 26460 67778 26516 67790
rect 26796 67844 26852 67854
rect 27020 67844 27076 67854
rect 26796 67842 27076 67844
rect 26796 67790 26798 67842
rect 26850 67790 27022 67842
rect 27074 67790 27076 67842
rect 26796 67788 27076 67790
rect 26796 67778 26852 67788
rect 27020 67778 27076 67788
rect 26236 66782 26238 66834
rect 26290 66782 26292 66834
rect 26236 66770 26292 66782
rect 26348 67618 26404 67630
rect 26348 67566 26350 67618
rect 26402 67566 26404 67618
rect 26348 65380 26404 67566
rect 26572 67060 26628 67070
rect 26572 66946 26628 67004
rect 26572 66894 26574 66946
rect 26626 66894 26628 66946
rect 26572 66882 26628 66894
rect 26684 67058 26740 67070
rect 26684 67006 26686 67058
rect 26738 67006 26740 67058
rect 26684 66948 26740 67006
rect 25900 65324 26404 65380
rect 26460 66052 26516 66062
rect 26684 66052 26740 66892
rect 26796 66052 26852 66062
rect 26460 66050 26852 66052
rect 26460 65998 26462 66050
rect 26514 65998 26798 66050
rect 26850 65998 26852 66050
rect 26460 65996 26852 65998
rect 25900 64708 25956 65324
rect 26124 64820 26180 64830
rect 25676 64706 25956 64708
rect 25676 64654 25902 64706
rect 25954 64654 25956 64706
rect 25676 64652 25956 64654
rect 25676 63922 25732 64652
rect 25900 64642 25956 64652
rect 26012 64818 26180 64820
rect 26012 64766 26126 64818
rect 26178 64766 26180 64818
rect 26012 64764 26180 64766
rect 26012 63924 26068 64764
rect 26124 64754 26180 64764
rect 26236 64148 26292 64158
rect 26236 64034 26292 64092
rect 26236 63982 26238 64034
rect 26290 63982 26292 64034
rect 26236 63970 26292 63982
rect 25676 63870 25678 63922
rect 25730 63870 25732 63922
rect 25676 63858 25732 63870
rect 25900 63922 26068 63924
rect 25900 63870 26014 63922
rect 26066 63870 26068 63922
rect 25900 63868 26068 63870
rect 25788 63812 25844 63822
rect 25788 63718 25844 63756
rect 25900 63588 25956 63868
rect 26012 63858 26068 63868
rect 25676 63532 25956 63588
rect 25676 63250 25732 63532
rect 25676 63198 25678 63250
rect 25730 63198 25732 63250
rect 25676 63186 25732 63198
rect 26348 63138 26404 63150
rect 26348 63086 26350 63138
rect 26402 63086 26404 63138
rect 26348 63028 26404 63086
rect 26348 62962 26404 62972
rect 25340 61618 25396 61628
rect 25452 62132 25620 62188
rect 25676 62916 25732 62926
rect 24892 61506 24948 61516
rect 24892 61346 24948 61358
rect 24892 61294 24894 61346
rect 24946 61294 24948 61346
rect 24556 60844 24836 60900
rect 24556 60676 24612 60686
rect 24500 60674 24612 60676
rect 24500 60622 24558 60674
rect 24610 60622 24612 60674
rect 24500 60620 24612 60622
rect 24444 60582 24500 60620
rect 24556 60610 24612 60620
rect 24668 60004 24724 60014
rect 24220 60002 24724 60004
rect 24220 59950 24670 60002
rect 24722 59950 24724 60002
rect 24220 59948 24724 59950
rect 24220 59442 24276 59948
rect 24668 59938 24724 59948
rect 24220 59390 24222 59442
rect 24274 59390 24276 59442
rect 24220 59378 24276 59390
rect 24556 59220 24612 59230
rect 24108 59218 24612 59220
rect 24108 59166 24558 59218
rect 24610 59166 24612 59218
rect 24108 59164 24612 59166
rect 23996 58818 24052 58828
rect 24220 58996 24276 59006
rect 24108 58436 24164 58446
rect 23884 58434 24164 58436
rect 23884 58382 24110 58434
rect 24162 58382 24164 58434
rect 23884 58380 24164 58382
rect 23884 58212 23940 58222
rect 23884 58118 23940 58156
rect 23772 57710 23774 57762
rect 23826 57710 23828 57762
rect 23772 57698 23828 57710
rect 23884 57876 23940 57886
rect 23436 57036 23828 57092
rect 23324 56924 23604 56980
rect 23100 55300 23156 56924
rect 23212 56642 23268 56654
rect 23212 56590 23214 56642
rect 23266 56590 23268 56642
rect 23212 56420 23268 56590
rect 23212 56354 23268 56364
rect 23100 55298 23380 55300
rect 23100 55246 23102 55298
rect 23154 55246 23380 55298
rect 23100 55244 23380 55246
rect 23100 55234 23156 55244
rect 22876 55188 22932 55198
rect 22764 55076 22820 55086
rect 22876 55076 22932 55132
rect 22988 55076 23044 55086
rect 22876 55074 23044 55076
rect 22876 55022 22990 55074
rect 23042 55022 23044 55074
rect 22876 55020 23044 55022
rect 22764 54982 22820 55020
rect 22988 55010 23044 55020
rect 22540 54796 23156 54852
rect 22428 54740 22484 54750
rect 22428 54646 22484 54684
rect 22988 54516 23044 54526
rect 22316 53778 22372 53788
rect 22428 54514 23044 54516
rect 22428 54462 22990 54514
rect 23042 54462 23044 54514
rect 22428 54460 23044 54462
rect 21532 53732 21588 53742
rect 21532 53638 21588 53676
rect 21420 53620 21476 53630
rect 20972 53618 21476 53620
rect 20972 53566 21422 53618
rect 21474 53566 21476 53618
rect 20972 53564 21476 53566
rect 20972 53170 21028 53564
rect 21420 53554 21476 53564
rect 20972 53118 20974 53170
rect 21026 53118 21028 53170
rect 20972 53106 21028 53118
rect 21868 53060 21924 53070
rect 21756 53058 21924 53060
rect 21756 53006 21870 53058
rect 21922 53006 21924 53058
rect 21756 53004 21924 53006
rect 20860 52892 21140 52948
rect 20412 51998 20414 52050
rect 20466 51998 20468 52050
rect 20412 51492 20468 51998
rect 20748 51604 20804 52892
rect 20860 51604 20916 51614
rect 20748 51602 20916 51604
rect 20748 51550 20862 51602
rect 20914 51550 20916 51602
rect 20748 51548 20916 51550
rect 20860 51538 20916 51548
rect 20524 51492 20580 51502
rect 20412 51436 20524 51492
rect 20524 51398 20580 51436
rect 20636 51492 20692 51502
rect 20636 51490 20804 51492
rect 20636 51438 20638 51490
rect 20690 51438 20804 51490
rect 20636 51436 20804 51438
rect 20636 51426 20692 51436
rect 20748 50932 20804 51436
rect 20636 50876 20804 50932
rect 20636 50372 20692 50876
rect 20636 50306 20692 50316
rect 20748 50370 20804 50382
rect 20972 50372 21028 50382
rect 20748 50318 20750 50370
rect 20802 50318 20804 50370
rect 20412 50036 20468 50046
rect 20748 50036 20804 50318
rect 20300 49698 20356 49710
rect 20300 49646 20302 49698
rect 20354 49646 20356 49698
rect 20300 49364 20356 49646
rect 20300 49298 20356 49308
rect 20188 48962 20244 48972
rect 19516 48916 19572 48926
rect 19516 48822 19572 48860
rect 20188 48804 20244 48814
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19516 48020 19572 48030
rect 19516 45332 19572 47964
rect 19740 47572 19796 47582
rect 20188 47572 20244 48748
rect 20300 48020 20356 48030
rect 20300 47682 20356 47964
rect 20300 47630 20302 47682
rect 20354 47630 20356 47682
rect 20300 47618 20356 47630
rect 19740 47478 19796 47516
rect 20076 47516 20244 47572
rect 20076 47236 20132 47516
rect 20412 47458 20468 49980
rect 20636 49980 20804 50036
rect 20860 50316 20972 50372
rect 20636 49588 20692 49980
rect 20636 49522 20692 49532
rect 20748 49810 20804 49822
rect 20748 49758 20750 49810
rect 20802 49758 20804 49810
rect 20412 47406 20414 47458
rect 20466 47406 20468 47458
rect 20300 47236 20356 47246
rect 20076 47180 20244 47236
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20188 47068 20244 47180
rect 20300 47142 20356 47180
rect 20412 47068 20468 47406
rect 20748 49028 20804 49758
rect 20748 47236 20804 48972
rect 20748 47170 20804 47180
rect 20188 47012 20356 47068
rect 19836 47002 20100 47012
rect 19628 45668 19684 45678
rect 19628 45574 19684 45612
rect 20188 45668 20244 45678
rect 20188 45574 20244 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19516 45276 20132 45332
rect 19404 45266 19460 45276
rect 19180 44942 19182 44994
rect 19234 44942 19236 44994
rect 19180 44930 19236 44942
rect 19628 44996 19684 45006
rect 19628 44902 19684 44940
rect 18956 43810 19012 43820
rect 19516 44882 19572 44894
rect 19516 44830 19518 44882
rect 19570 44830 19572 44882
rect 18284 43764 18340 43774
rect 17948 43762 18340 43764
rect 17948 43710 18286 43762
rect 18338 43710 18340 43762
rect 17948 43708 18340 43710
rect 18284 43698 18340 43708
rect 19516 43762 19572 44830
rect 19852 44884 19908 44894
rect 19852 44790 19908 44828
rect 20076 44546 20132 45276
rect 20300 45220 20356 47012
rect 20412 47012 20692 47068
rect 20412 46004 20468 47012
rect 20636 46898 20692 47012
rect 20636 46846 20638 46898
rect 20690 46846 20692 46898
rect 20636 46834 20692 46846
rect 20748 46676 20804 46686
rect 20748 46582 20804 46620
rect 20412 45938 20468 45948
rect 20636 46452 20692 46462
rect 20636 45890 20692 46396
rect 20636 45838 20638 45890
rect 20690 45838 20692 45890
rect 20412 45220 20468 45230
rect 20300 45218 20468 45220
rect 20300 45166 20414 45218
rect 20466 45166 20468 45218
rect 20300 45164 20468 45166
rect 20412 44996 20468 45164
rect 20412 44930 20468 44940
rect 20524 45220 20580 45230
rect 20636 45220 20692 45838
rect 20748 45780 20804 45790
rect 20748 45686 20804 45724
rect 20748 45220 20804 45230
rect 20636 45218 20804 45220
rect 20636 45166 20750 45218
rect 20802 45166 20804 45218
rect 20636 45164 20804 45166
rect 20188 44884 20244 44894
rect 20188 44790 20244 44828
rect 20076 44494 20078 44546
rect 20130 44494 20132 44546
rect 20076 44482 20132 44494
rect 20188 44660 20244 44670
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43876 20244 44604
rect 20412 44436 20468 44446
rect 20412 44342 20468 44380
rect 20188 43810 20244 43820
rect 20300 44324 20356 44334
rect 20300 44098 20356 44268
rect 20300 44046 20302 44098
rect 20354 44046 20356 44098
rect 19516 43710 19518 43762
rect 19570 43710 19572 43762
rect 19516 43698 19572 43710
rect 20300 43762 20356 44046
rect 20300 43710 20302 43762
rect 20354 43710 20356 43762
rect 20300 43698 20356 43710
rect 16716 43598 16718 43650
rect 16770 43598 16772 43650
rect 16268 43260 16548 43316
rect 16268 41748 16324 43260
rect 16380 42868 16436 42878
rect 16380 42774 16436 42812
rect 16716 42644 16772 43598
rect 18508 43650 18564 43662
rect 18508 43598 18510 43650
rect 18562 43598 18564 43650
rect 16380 42588 16772 42644
rect 16828 43540 16884 43550
rect 16380 42308 16436 42588
rect 16380 42082 16436 42252
rect 16380 42030 16382 42082
rect 16434 42030 16436 42082
rect 16380 42018 16436 42030
rect 16492 42420 16548 42430
rect 16492 42194 16548 42364
rect 16492 42142 16494 42194
rect 16546 42142 16548 42194
rect 16268 41682 16324 41692
rect 16380 41860 16436 41870
rect 16380 41188 16436 41804
rect 16380 41094 16436 41132
rect 16156 40114 16212 40124
rect 16268 41074 16324 41086
rect 16268 41022 16270 41074
rect 16322 41022 16324 41074
rect 16268 39844 16324 41022
rect 16492 41076 16548 42142
rect 16716 41970 16772 41982
rect 16716 41918 16718 41970
rect 16770 41918 16772 41970
rect 16716 41186 16772 41918
rect 16716 41134 16718 41186
rect 16770 41134 16772 41186
rect 16716 41122 16772 41134
rect 16492 41010 16548 41020
rect 16380 40628 16436 40638
rect 16380 40626 16772 40628
rect 16380 40574 16382 40626
rect 16434 40574 16772 40626
rect 16380 40572 16772 40574
rect 16380 40562 16436 40572
rect 16716 40514 16772 40572
rect 16716 40462 16718 40514
rect 16770 40462 16772 40514
rect 16604 40402 16660 40414
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 16268 39778 16324 39788
rect 16492 40292 16548 40302
rect 16380 39730 16436 39742
rect 16380 39678 16382 39730
rect 16434 39678 16436 39730
rect 15372 38612 16100 38668
rect 16268 38834 16324 38846
rect 16268 38782 16270 38834
rect 16322 38782 16324 38834
rect 16268 38724 16324 38782
rect 16268 38658 16324 38668
rect 16380 38668 16436 39678
rect 16492 39060 16548 40236
rect 16604 40180 16660 40350
rect 16604 40114 16660 40124
rect 16492 38966 16548 39004
rect 16380 38612 16660 38668
rect 15372 38162 15428 38612
rect 15372 38110 15374 38162
rect 15426 38110 15428 38162
rect 15372 38098 15428 38110
rect 14588 36978 14644 36988
rect 14924 37324 15092 37380
rect 16268 37380 16324 37390
rect 14364 34290 14420 34300
rect 14588 36484 14644 36494
rect 14924 36484 14980 37324
rect 15708 37266 15764 37278
rect 15708 37214 15710 37266
rect 15762 37214 15764 37266
rect 14588 36482 14980 36484
rect 14588 36430 14590 36482
rect 14642 36430 14980 36482
rect 14588 36428 14980 36430
rect 15036 37156 15092 37166
rect 13916 34244 13972 34254
rect 13916 34150 13972 34188
rect 14364 34132 14420 34142
rect 13580 34018 13636 34030
rect 13580 33966 13582 34018
rect 13634 33966 13636 34018
rect 13580 33236 13636 33966
rect 14140 33684 14196 33694
rect 13804 33572 13860 33582
rect 14028 33572 14084 33582
rect 13804 33570 14028 33572
rect 13804 33518 13806 33570
rect 13858 33518 14028 33570
rect 13804 33516 14028 33518
rect 13804 33506 13860 33516
rect 13636 33180 13748 33236
rect 13580 33142 13636 33180
rect 13692 32564 13748 33180
rect 13804 32564 13860 32574
rect 13692 32562 13860 32564
rect 13692 32510 13806 32562
rect 13858 32510 13860 32562
rect 13692 32508 13860 32510
rect 13804 32498 13860 32508
rect 14028 32562 14084 33516
rect 14140 33570 14196 33628
rect 14140 33518 14142 33570
rect 14194 33518 14196 33570
rect 14140 33506 14196 33518
rect 14364 32786 14420 34076
rect 14364 32734 14366 32786
rect 14418 32734 14420 32786
rect 14364 32722 14420 32734
rect 14476 33460 14532 33470
rect 14028 32510 14030 32562
rect 14082 32510 14084 32562
rect 14028 32498 14084 32510
rect 13468 31714 13524 31724
rect 14028 30996 14084 31006
rect 14028 30902 14084 30940
rect 14364 30994 14420 31006
rect 14364 30942 14366 30994
rect 14418 30942 14420 30994
rect 14028 30436 14084 30446
rect 14028 28196 14084 30380
rect 14140 30324 14196 30334
rect 14140 30230 14196 30268
rect 14364 30212 14420 30942
rect 14364 30146 14420 30156
rect 14476 30154 14532 33404
rect 14588 32116 14644 36428
rect 14700 34130 14756 34142
rect 14700 34078 14702 34130
rect 14754 34078 14756 34130
rect 14700 33572 14756 34078
rect 14700 33458 14756 33516
rect 14700 33406 14702 33458
rect 14754 33406 14756 33458
rect 14700 33394 14756 33406
rect 14924 33796 14980 33806
rect 14924 33346 14980 33740
rect 14924 33294 14926 33346
rect 14978 33294 14980 33346
rect 14812 33236 14868 33246
rect 14588 32050 14644 32060
rect 14700 33180 14812 33236
rect 14700 32004 14756 33180
rect 14812 33142 14868 33180
rect 14924 33012 14980 33294
rect 14700 31938 14756 31948
rect 14812 32956 14980 33012
rect 14588 31780 14644 31790
rect 14588 31778 14756 31780
rect 14588 31726 14590 31778
rect 14642 31726 14756 31778
rect 14588 31724 14756 31726
rect 14588 31714 14644 31724
rect 14700 31668 14756 31724
rect 14700 31602 14756 31612
rect 14812 31444 14868 32956
rect 14924 31780 14980 31790
rect 14924 31686 14980 31724
rect 14812 31378 14868 31388
rect 15036 31332 15092 37100
rect 15372 37156 15428 37166
rect 15708 37156 15764 37214
rect 16268 37266 16324 37324
rect 16268 37214 16270 37266
rect 16322 37214 16324 37266
rect 16268 37202 16324 37214
rect 15428 37100 15764 37156
rect 15372 37062 15428 37100
rect 16044 34916 16100 34926
rect 16044 34822 16100 34860
rect 15932 34804 15988 34814
rect 15484 34690 15540 34702
rect 15484 34638 15486 34690
rect 15538 34638 15540 34690
rect 15484 33460 15540 34638
rect 15932 34242 15988 34748
rect 16380 34692 16436 34702
rect 15932 34190 15934 34242
rect 15986 34190 15988 34242
rect 15932 34178 15988 34190
rect 16044 34690 16436 34692
rect 16044 34638 16382 34690
rect 16434 34638 16436 34690
rect 16044 34636 16436 34638
rect 15484 33394 15540 33404
rect 15820 34020 15876 34030
rect 15820 32676 15876 33964
rect 16044 33236 16100 34636
rect 16380 34626 16436 34636
rect 16492 34244 16548 34254
rect 16492 34150 16548 34188
rect 16268 34132 16324 34142
rect 16268 34038 16324 34076
rect 16380 34020 16436 34030
rect 16380 33926 16436 33964
rect 16044 33170 16100 33180
rect 16268 33234 16324 33246
rect 16268 33182 16270 33234
rect 16322 33182 16324 33234
rect 15708 32674 15876 32676
rect 15708 32622 15822 32674
rect 15874 32622 15876 32674
rect 15708 32620 15876 32622
rect 15708 31892 15764 32620
rect 15820 32610 15876 32620
rect 16044 32340 16100 32350
rect 16268 32340 16324 33182
rect 16044 32338 16324 32340
rect 16044 32286 16046 32338
rect 16098 32286 16324 32338
rect 16044 32284 16324 32286
rect 16044 32274 16100 32284
rect 15708 31798 15764 31836
rect 16156 31892 16212 31902
rect 15372 31780 15428 31790
rect 15036 31266 15092 31276
rect 15260 31332 15316 31342
rect 14924 30996 14980 31006
rect 14924 30994 15204 30996
rect 14924 30942 14926 30994
rect 14978 30942 15204 30994
rect 14924 30940 15204 30942
rect 14924 30930 14980 30940
rect 15148 30884 15204 30940
rect 15260 30884 15316 31276
rect 15148 30828 15316 30884
rect 15148 30324 15204 30334
rect 15036 30268 15148 30324
rect 14476 30102 14478 30154
rect 14530 30102 14532 30154
rect 14812 30212 14868 30222
rect 14812 30118 14868 30156
rect 14476 28644 14532 30102
rect 14588 29988 14644 29998
rect 14588 29894 14644 29932
rect 15036 29764 15092 30268
rect 15148 30230 15204 30268
rect 14588 29708 15092 29764
rect 14588 29316 14644 29708
rect 14812 29596 15092 29652
rect 14700 29540 14756 29550
rect 14700 29446 14756 29484
rect 14812 29538 14868 29596
rect 14812 29486 14814 29538
rect 14866 29486 14868 29538
rect 14812 29474 14868 29486
rect 15036 29316 15092 29596
rect 15260 29540 15316 30828
rect 15372 30884 15428 31724
rect 15372 30790 15428 30828
rect 16044 31666 16100 31678
rect 16044 31614 16046 31666
rect 16098 31614 16100 31666
rect 16044 31108 16100 31614
rect 16044 30322 16100 31052
rect 16156 30994 16212 31836
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 16156 30930 16212 30942
rect 16268 30884 16324 32284
rect 16380 32338 16436 32350
rect 16380 32286 16382 32338
rect 16434 32286 16436 32338
rect 16380 30996 16436 32286
rect 16380 30930 16436 30940
rect 16268 30772 16324 30828
rect 16380 30772 16436 30782
rect 16268 30770 16436 30772
rect 16268 30718 16382 30770
rect 16434 30718 16436 30770
rect 16268 30716 16436 30718
rect 16380 30706 16436 30716
rect 16604 30548 16660 38612
rect 16716 36932 16772 40462
rect 16828 38668 16884 43484
rect 18172 43428 18228 43438
rect 18508 43428 18564 43598
rect 20188 43650 20244 43662
rect 20188 43598 20190 43650
rect 20242 43598 20244 43650
rect 18172 43426 18564 43428
rect 18172 43374 18174 43426
rect 18226 43374 18564 43426
rect 18172 43372 18564 43374
rect 18172 43362 18228 43372
rect 18508 43092 18564 43372
rect 18620 43538 18676 43550
rect 18620 43486 18622 43538
rect 18674 43486 18676 43538
rect 18620 43316 18676 43486
rect 19852 43538 19908 43550
rect 19852 43486 19854 43538
rect 19906 43486 19908 43538
rect 18620 43250 18676 43260
rect 18956 43426 19012 43438
rect 18956 43374 18958 43426
rect 19010 43374 19012 43426
rect 18956 43092 19012 43374
rect 18508 43036 19012 43092
rect 18844 42532 18900 42542
rect 18956 42532 19012 43036
rect 18900 42476 19012 42532
rect 19180 43316 19236 43326
rect 17500 41858 17556 41870
rect 17500 41806 17502 41858
rect 17554 41806 17556 41858
rect 17500 41300 17556 41806
rect 17836 41300 17892 41310
rect 17500 41298 17892 41300
rect 17500 41246 17838 41298
rect 17890 41246 17892 41298
rect 17500 41244 17892 41246
rect 17052 41188 17108 41198
rect 16940 41186 17108 41188
rect 16940 41134 17054 41186
rect 17106 41134 17108 41186
rect 16940 41132 17108 41134
rect 16940 40626 16996 41132
rect 17052 41122 17108 41132
rect 17276 41188 17332 41198
rect 17500 41188 17556 41244
rect 17836 41234 17892 41244
rect 17332 41132 17556 41188
rect 17276 41094 17332 41132
rect 17052 40962 17108 40974
rect 17052 40910 17054 40962
rect 17106 40910 17108 40962
rect 17052 40852 17108 40910
rect 17052 40786 17108 40796
rect 18060 40852 18116 40862
rect 18116 40796 18228 40852
rect 18060 40786 18116 40796
rect 16940 40574 16942 40626
rect 16994 40574 16996 40626
rect 16940 40562 16996 40574
rect 17500 40628 17556 40638
rect 17500 40402 17556 40572
rect 18172 40514 18228 40796
rect 18172 40462 18174 40514
rect 18226 40462 18228 40514
rect 18172 40450 18228 40462
rect 17500 40350 17502 40402
rect 17554 40350 17556 40402
rect 17500 40292 17556 40350
rect 17500 40226 17556 40236
rect 17276 40180 17332 40190
rect 16940 39844 16996 39854
rect 16940 39618 16996 39788
rect 16940 39566 16942 39618
rect 16994 39566 16996 39618
rect 16940 39554 16996 39566
rect 17276 39618 17332 40124
rect 17276 39566 17278 39618
rect 17330 39566 17332 39618
rect 17276 39554 17332 39566
rect 17164 39394 17220 39406
rect 17164 39342 17166 39394
rect 17218 39342 17220 39394
rect 17164 39284 17220 39342
rect 17836 39394 17892 39406
rect 17836 39342 17838 39394
rect 17890 39342 17892 39394
rect 17836 39284 17892 39342
rect 17164 39228 17892 39284
rect 16828 38612 16996 38668
rect 16716 36866 16772 36876
rect 16716 35028 16772 35038
rect 16716 34802 16772 34972
rect 16716 34750 16718 34802
rect 16770 34750 16772 34802
rect 16716 34738 16772 34750
rect 16828 34130 16884 34142
rect 16828 34078 16830 34130
rect 16882 34078 16884 34130
rect 16828 33684 16884 34078
rect 16828 33618 16884 33628
rect 16940 32340 16996 38612
rect 17500 38162 17556 38174
rect 17500 38110 17502 38162
rect 17554 38110 17556 38162
rect 17164 36372 17220 36382
rect 17164 36370 17444 36372
rect 17164 36318 17166 36370
rect 17218 36318 17444 36370
rect 17164 36316 17444 36318
rect 17164 36306 17220 36316
rect 17388 36258 17444 36316
rect 17388 36206 17390 36258
rect 17442 36206 17444 36258
rect 17052 35364 17108 35374
rect 17052 32900 17108 35308
rect 17388 34692 17444 36206
rect 17500 35924 17556 38110
rect 17836 36820 17892 39228
rect 18844 38668 18900 42476
rect 18956 41972 19012 41982
rect 18956 41858 19012 41916
rect 18956 41806 18958 41858
rect 19010 41806 19012 41858
rect 18956 41410 19012 41806
rect 18956 41358 18958 41410
rect 19010 41358 19012 41410
rect 18956 41346 19012 41358
rect 19180 41858 19236 43260
rect 19852 43316 19908 43486
rect 19852 43250 19908 43260
rect 20076 42644 20132 42654
rect 19740 42532 19796 42570
rect 20076 42550 20132 42588
rect 19740 42466 19796 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19628 41972 19684 41982
rect 19628 41878 19684 41916
rect 19180 41806 19182 41858
rect 19234 41806 19236 41858
rect 18620 38612 18676 38622
rect 18508 38052 18564 38062
rect 18284 38050 18564 38052
rect 18284 37998 18510 38050
rect 18562 37998 18564 38050
rect 18284 37996 18564 37998
rect 18172 37938 18228 37950
rect 18172 37886 18174 37938
rect 18226 37886 18228 37938
rect 17836 36754 17892 36764
rect 18060 37492 18116 37502
rect 17948 36596 18004 36606
rect 18060 36596 18116 37436
rect 17500 35858 17556 35868
rect 17612 36594 18116 36596
rect 17612 36542 17950 36594
rect 18002 36542 18116 36594
rect 17612 36540 18116 36542
rect 17500 35700 17556 35710
rect 17612 35700 17668 36540
rect 17948 36530 18004 36540
rect 18172 36260 18228 37886
rect 18284 37490 18340 37996
rect 18508 37986 18564 37996
rect 18508 37492 18564 37502
rect 18620 37492 18676 38556
rect 18284 37438 18286 37490
rect 18338 37438 18340 37490
rect 18284 37426 18340 37438
rect 18396 37436 18508 37492
rect 18564 37436 18676 37492
rect 18732 38612 18900 38668
rect 18956 41188 19012 41198
rect 18396 36594 18452 37436
rect 18508 37398 18564 37436
rect 18620 37268 18676 37278
rect 18396 36542 18398 36594
rect 18450 36542 18452 36594
rect 18396 36530 18452 36542
rect 18508 37266 18676 37268
rect 18508 37214 18622 37266
rect 18674 37214 18676 37266
rect 18508 37212 18676 37214
rect 18284 36260 18340 36270
rect 18172 36204 18284 36260
rect 18284 36194 18340 36204
rect 18508 36036 18564 37212
rect 18620 37202 18676 37212
rect 17724 35980 18676 36036
rect 17724 35922 17780 35980
rect 17724 35870 17726 35922
rect 17778 35870 17780 35922
rect 17724 35858 17780 35870
rect 17948 35812 18004 35822
rect 17500 35698 17668 35700
rect 17500 35646 17502 35698
rect 17554 35646 17668 35698
rect 17500 35644 17668 35646
rect 17724 35700 17780 35710
rect 17500 35634 17556 35644
rect 17388 34598 17444 34636
rect 17724 34580 17780 35644
rect 17836 35588 17892 35598
rect 17836 35494 17892 35532
rect 17948 35364 18004 35756
rect 18172 35698 18228 35710
rect 18172 35646 18174 35698
rect 18226 35646 18228 35698
rect 18172 35476 18228 35646
rect 18396 35476 18452 35486
rect 18172 35420 18396 35476
rect 17836 35308 18004 35364
rect 17836 35028 17892 35308
rect 17836 34914 17892 34972
rect 17836 34862 17838 34914
rect 17890 34862 17892 34914
rect 17836 34850 17892 34862
rect 17948 34916 18004 34926
rect 17948 34802 18004 34860
rect 17948 34750 17950 34802
rect 18002 34750 18004 34802
rect 17724 34524 17892 34580
rect 17724 34356 17780 34366
rect 17724 34262 17780 34300
rect 17388 34130 17444 34142
rect 17388 34078 17390 34130
rect 17442 34078 17444 34130
rect 17388 33796 17444 34078
rect 17388 33730 17444 33740
rect 17164 33124 17220 33134
rect 17164 33122 17668 33124
rect 17164 33070 17166 33122
rect 17218 33070 17668 33122
rect 17164 33068 17668 33070
rect 17164 33058 17220 33068
rect 17052 32844 17220 32900
rect 17052 32340 17108 32350
rect 16940 32284 17052 32340
rect 17052 32274 17108 32284
rect 16716 30884 16772 30894
rect 16716 30790 16772 30828
rect 16492 30492 16660 30548
rect 16044 30270 16046 30322
rect 16098 30270 16100 30322
rect 16044 30258 16100 30270
rect 16380 30324 16436 30334
rect 16380 30230 16436 30268
rect 15596 30212 15652 30222
rect 15596 30118 15652 30156
rect 16492 30100 16548 30492
rect 16380 30044 16548 30100
rect 16604 30322 16660 30334
rect 16604 30270 16606 30322
rect 16658 30270 16660 30322
rect 15260 29484 15540 29540
rect 15372 29316 15428 29326
rect 14588 29260 14868 29316
rect 15036 29314 15428 29316
rect 15036 29262 15374 29314
rect 15426 29262 15428 29314
rect 15036 29260 15428 29262
rect 14812 29202 14868 29260
rect 14812 29150 14814 29202
rect 14866 29150 14868 29202
rect 14812 29138 14868 29150
rect 14588 28644 14644 28654
rect 14476 28642 14644 28644
rect 14476 28590 14590 28642
rect 14642 28590 14644 28642
rect 14476 28588 14644 28590
rect 14588 28578 14644 28588
rect 14028 28130 14084 28140
rect 14700 28532 14756 28542
rect 13580 27972 13636 27982
rect 13468 27916 13580 27972
rect 13468 26290 13524 27916
rect 13580 27906 13636 27916
rect 14476 27972 14532 27982
rect 14476 27878 14532 27916
rect 13804 27748 13860 27758
rect 13580 27076 13636 27114
rect 13580 27010 13636 27020
rect 13804 27074 13860 27692
rect 14700 27412 14756 28476
rect 14924 28420 14980 28430
rect 14924 28326 14980 28364
rect 15260 28420 15316 28430
rect 14588 27356 14756 27412
rect 14812 27858 14868 27870
rect 14812 27806 14814 27858
rect 14866 27806 14868 27858
rect 13804 27022 13806 27074
rect 13858 27022 13860 27074
rect 13804 27010 13860 27022
rect 13916 27076 13972 27086
rect 13468 26238 13470 26290
rect 13522 26238 13524 26290
rect 13468 26226 13524 26238
rect 13580 26852 13636 26862
rect 13580 24948 13636 26796
rect 13804 26516 13860 26526
rect 13916 26516 13972 27020
rect 14476 26964 14532 27002
rect 14476 26898 14532 26908
rect 13804 26514 13972 26516
rect 13804 26462 13806 26514
rect 13858 26462 13972 26514
rect 13804 26460 13972 26462
rect 14476 26516 14532 26526
rect 14588 26516 14644 27356
rect 14700 27188 14756 27198
rect 14812 27188 14868 27806
rect 14756 27132 14868 27188
rect 15260 27860 15316 28364
rect 14700 27122 14756 27132
rect 14476 26514 14644 26516
rect 14476 26462 14478 26514
rect 14530 26462 14644 26514
rect 14476 26460 14644 26462
rect 13804 26450 13860 26460
rect 14476 26450 14532 26460
rect 14140 26404 14196 26414
rect 14140 26402 14308 26404
rect 14140 26350 14142 26402
rect 14194 26350 14308 26402
rect 14140 26348 14308 26350
rect 14140 26338 14196 26348
rect 14252 25956 14308 26348
rect 15260 26290 15316 27804
rect 15260 26238 15262 26290
rect 15314 26238 15316 26290
rect 15260 26226 15316 26238
rect 15148 26178 15204 26190
rect 15148 26126 15150 26178
rect 15202 26126 15204 26178
rect 14252 25900 14868 25956
rect 14252 25732 14308 25742
rect 14252 25638 14308 25676
rect 14140 25508 14196 25518
rect 14364 25508 14420 25518
rect 14700 25508 14756 25518
rect 14140 25506 14364 25508
rect 14140 25454 14142 25506
rect 14194 25454 14364 25506
rect 14140 25452 14364 25454
rect 14420 25506 14756 25508
rect 14420 25454 14702 25506
rect 14754 25454 14756 25506
rect 14420 25452 14756 25454
rect 14140 25442 14196 25452
rect 14364 25414 14420 25452
rect 14700 25442 14756 25452
rect 14812 25394 14868 25900
rect 15148 25732 15204 26126
rect 15148 25666 15204 25676
rect 15036 25396 15092 25406
rect 14812 25342 14814 25394
rect 14866 25342 14868 25394
rect 14252 25284 14308 25294
rect 14252 25190 14308 25228
rect 14700 25284 14756 25294
rect 13356 23214 13358 23266
rect 13410 23214 13412 23266
rect 12908 22430 12910 22482
rect 12962 22430 12964 22482
rect 12908 22418 12964 22430
rect 13020 23042 13076 23054
rect 13020 22990 13022 23042
rect 13074 22990 13076 23042
rect 13020 21140 13076 22990
rect 13356 22372 13412 23214
rect 13356 22306 13412 22316
rect 13468 24892 14532 24948
rect 13468 21812 13524 24892
rect 14364 24724 14420 24734
rect 13916 24722 14420 24724
rect 13916 24670 14366 24722
rect 14418 24670 14420 24722
rect 13916 24668 14420 24670
rect 13804 24500 13860 24510
rect 13580 24498 13860 24500
rect 13580 24446 13806 24498
rect 13858 24446 13860 24498
rect 13580 24444 13860 24446
rect 13580 23938 13636 24444
rect 13804 24434 13860 24444
rect 13580 23886 13582 23938
rect 13634 23886 13636 23938
rect 13580 23874 13636 23886
rect 13804 23828 13860 23838
rect 13916 23828 13972 24668
rect 14364 24658 14420 24668
rect 14028 24388 14084 24398
rect 14084 24332 14196 24388
rect 14028 24322 14084 24332
rect 13804 23826 13972 23828
rect 13804 23774 13806 23826
rect 13858 23774 13972 23826
rect 13804 23772 13972 23774
rect 13804 23762 13860 23772
rect 13804 23604 13860 23614
rect 13692 23548 13804 23604
rect 13580 21812 13636 21822
rect 13468 21810 13636 21812
rect 13468 21758 13582 21810
rect 13634 21758 13636 21810
rect 13468 21756 13636 21758
rect 13580 21746 13636 21756
rect 12124 20514 12180 20524
rect 12236 21084 13076 21140
rect 12236 20188 12292 21084
rect 12684 20916 12740 20926
rect 11788 20132 12292 20188
rect 12572 20860 12684 20916
rect 11340 19404 11732 19460
rect 11228 19182 11230 19234
rect 11282 19182 11284 19234
rect 11004 19012 11060 19022
rect 11004 19010 11172 19012
rect 11004 18958 11006 19010
rect 11058 18958 11172 19010
rect 11004 18956 11172 18958
rect 11004 18946 11060 18956
rect 10668 18564 10724 18574
rect 11004 18564 11060 18574
rect 10668 18562 11004 18564
rect 10668 18510 10670 18562
rect 10722 18510 11004 18562
rect 10668 18508 11004 18510
rect 10668 18498 10724 18508
rect 11004 18470 11060 18508
rect 10556 18398 10558 18450
rect 10610 18398 10612 18450
rect 10556 18386 10612 18398
rect 11116 18452 11172 18956
rect 11116 18386 11172 18396
rect 11228 18674 11284 19182
rect 11564 19236 11620 19246
rect 11340 19124 11396 19134
rect 11340 19030 11396 19068
rect 11452 19012 11508 19022
rect 11452 18918 11508 18956
rect 11228 18622 11230 18674
rect 11282 18622 11284 18674
rect 11004 18340 11060 18350
rect 11004 17780 11060 18284
rect 11116 17780 11172 17790
rect 11004 17778 11172 17780
rect 11004 17726 11118 17778
rect 11170 17726 11172 17778
rect 11004 17724 11172 17726
rect 11116 17714 11172 17724
rect 9548 17490 9604 17500
rect 11116 17556 11172 17566
rect 11116 16994 11172 17500
rect 11228 17220 11284 18622
rect 11340 18228 11396 18238
rect 11340 18134 11396 18172
rect 11228 17164 11396 17220
rect 11116 16942 11118 16994
rect 11170 16942 11172 16994
rect 11116 16930 11172 16942
rect 11228 16994 11284 17006
rect 11228 16942 11230 16994
rect 11282 16942 11284 16994
rect 8988 16034 9044 16044
rect 10444 16100 10500 16110
rect 10668 16100 10724 16110
rect 10500 16098 10724 16100
rect 10500 16046 10670 16098
rect 10722 16046 10724 16098
rect 10500 16044 10724 16046
rect 10444 16006 10500 16044
rect 10668 16034 10724 16044
rect 11004 15876 11060 15886
rect 11228 15876 11284 16942
rect 11060 15820 11284 15876
rect 11004 15782 11060 15820
rect 11340 15652 11396 17164
rect 11340 15586 11396 15596
rect 11452 16882 11508 16894
rect 11452 16830 11454 16882
rect 11506 16830 11508 16882
rect 11452 16098 11508 16830
rect 11452 16046 11454 16098
rect 11506 16046 11508 16098
rect 11452 15428 11508 16046
rect 11564 16100 11620 19180
rect 11676 16884 11732 19404
rect 11676 16818 11732 16828
rect 11788 19234 11844 20132
rect 11788 19182 11790 19234
rect 11842 19182 11844 19234
rect 11788 16100 11844 19182
rect 11900 20018 11956 20030
rect 11900 19966 11902 20018
rect 11954 19966 11956 20018
rect 11900 18564 11956 19966
rect 12348 19908 12404 19918
rect 12124 19906 12404 19908
rect 12124 19854 12350 19906
rect 12402 19854 12404 19906
rect 12124 19852 12404 19854
rect 12012 19236 12068 19246
rect 12012 19142 12068 19180
rect 11900 18498 11956 18508
rect 12124 19012 12180 19852
rect 12348 19842 12404 19852
rect 12460 19236 12516 19246
rect 12572 19236 12628 20860
rect 12684 20850 12740 20860
rect 12796 20132 12852 20142
rect 12460 19234 12740 19236
rect 12460 19182 12462 19234
rect 12514 19182 12740 19234
rect 12460 19180 12740 19182
rect 12460 19170 12516 19180
rect 12124 18004 12180 18956
rect 12236 19012 12292 19022
rect 12572 19012 12628 19022
rect 12236 19010 12404 19012
rect 12236 18958 12238 19010
rect 12290 18958 12404 19010
rect 12236 18956 12404 18958
rect 12236 18946 12292 18956
rect 12236 18564 12292 18574
rect 12236 18470 12292 18508
rect 12012 17948 12180 18004
rect 12236 18340 12292 18350
rect 11900 16100 11956 16110
rect 11564 16098 11732 16100
rect 11564 16046 11566 16098
rect 11618 16046 11732 16098
rect 11564 16044 11732 16046
rect 11788 16098 11956 16100
rect 11788 16046 11902 16098
rect 11954 16046 11956 16098
rect 11788 16044 11956 16046
rect 11564 16034 11620 16044
rect 11452 15334 11508 15372
rect 11564 15540 11620 15550
rect 11564 15426 11620 15484
rect 11564 15374 11566 15426
rect 11618 15374 11620 15426
rect 11564 15362 11620 15374
rect 11676 15426 11732 16044
rect 11676 15374 11678 15426
rect 11730 15374 11732 15426
rect 11676 15362 11732 15374
rect 11788 15874 11844 15886
rect 11788 15822 11790 15874
rect 11842 15822 11844 15874
rect 11004 15092 11060 15102
rect 11788 15092 11844 15822
rect 11900 15540 11956 16044
rect 11900 15474 11956 15484
rect 11004 15090 11172 15092
rect 11004 15038 11006 15090
rect 11058 15038 11172 15090
rect 11004 15036 11172 15038
rect 11004 15026 11060 15036
rect 11116 14530 11172 15036
rect 11564 15036 11844 15092
rect 11564 14642 11620 15036
rect 12012 14980 12068 17948
rect 12236 16324 12292 18284
rect 12348 17108 12404 18956
rect 12572 18918 12628 18956
rect 12460 18450 12516 18462
rect 12460 18398 12462 18450
rect 12514 18398 12516 18450
rect 12460 18228 12516 18398
rect 12684 18228 12740 19180
rect 12796 18564 12852 20076
rect 13692 19572 13748 23548
rect 13804 23538 13860 23548
rect 13916 23268 13972 23278
rect 13916 23174 13972 23212
rect 13916 21924 13972 21934
rect 13916 21810 13972 21868
rect 13916 21758 13918 21810
rect 13970 21758 13972 21810
rect 13916 21746 13972 21758
rect 14028 20020 14084 20030
rect 13804 19796 13860 19806
rect 13804 19794 13972 19796
rect 13804 19742 13806 19794
rect 13858 19742 13972 19794
rect 13804 19740 13972 19742
rect 13804 19730 13860 19740
rect 13692 19516 13860 19572
rect 13468 19124 13524 19134
rect 13468 19030 13524 19068
rect 12908 19010 12964 19022
rect 12908 18958 12910 19010
rect 12962 18958 12964 19010
rect 12908 18676 12964 18958
rect 13692 19012 13748 19022
rect 13692 18918 13748 18956
rect 12908 18610 12964 18620
rect 12796 18498 12852 18508
rect 13244 18452 13300 18462
rect 13244 18358 13300 18396
rect 12684 18172 13300 18228
rect 12460 18162 12516 18172
rect 12348 17052 12964 17108
rect 12348 16884 12404 16894
rect 12404 16828 12516 16884
rect 12348 16818 12404 16828
rect 12348 16324 12404 16334
rect 12124 16322 12404 16324
rect 12124 16270 12350 16322
rect 12402 16270 12404 16322
rect 12124 16268 12404 16270
rect 12124 15538 12180 16268
rect 12348 16258 12404 16268
rect 12236 16100 12292 16110
rect 12460 16100 12516 16828
rect 12236 16098 12852 16100
rect 12236 16046 12238 16098
rect 12290 16046 12852 16098
rect 12236 16044 12852 16046
rect 12236 16034 12292 16044
rect 12348 15876 12404 15886
rect 12404 15820 12516 15876
rect 12348 15782 12404 15820
rect 12124 15486 12126 15538
rect 12178 15486 12180 15538
rect 12124 15474 12180 15486
rect 12348 15652 12404 15662
rect 12348 15538 12404 15596
rect 12348 15486 12350 15538
rect 12402 15486 12404 15538
rect 12348 15474 12404 15486
rect 11564 14590 11566 14642
rect 11618 14590 11620 14642
rect 11564 14578 11620 14590
rect 11788 14924 12068 14980
rect 12236 15202 12292 15214
rect 12236 15150 12238 15202
rect 12290 15150 12292 15202
rect 11116 14478 11118 14530
rect 11170 14478 11172 14530
rect 11116 14466 11172 14478
rect 11788 13746 11844 14924
rect 12236 14644 12292 15150
rect 12348 14644 12404 14654
rect 12236 14642 12404 14644
rect 12236 14590 12350 14642
rect 12402 14590 12404 14642
rect 12236 14588 12404 14590
rect 12348 14578 12404 14588
rect 11788 13694 11790 13746
rect 11842 13694 11844 13746
rect 11788 13412 11844 13694
rect 11900 14308 11956 14318
rect 11900 13634 11956 14252
rect 12012 13860 12068 13870
rect 12460 13860 12516 15820
rect 12572 15540 12628 15550
rect 12572 15446 12628 15484
rect 12572 14532 12628 14542
rect 12572 14438 12628 14476
rect 12684 13860 12740 13870
rect 12012 13858 12740 13860
rect 12012 13806 12014 13858
rect 12066 13806 12686 13858
rect 12738 13806 12740 13858
rect 12012 13804 12740 13806
rect 12012 13794 12068 13804
rect 12684 13794 12740 13804
rect 11900 13582 11902 13634
rect 11954 13582 11956 13634
rect 11900 13570 11956 13582
rect 12348 13636 12404 13646
rect 11788 13356 11956 13412
rect 11228 11732 11284 11742
rect 11228 11394 11284 11676
rect 11228 11342 11230 11394
rect 11282 11342 11284 11394
rect 11228 11330 11284 11342
rect 11564 11396 11620 11406
rect 11788 11396 11844 11406
rect 11564 11394 11844 11396
rect 11564 11342 11566 11394
rect 11618 11342 11790 11394
rect 11842 11342 11844 11394
rect 11564 11340 11844 11342
rect 11564 11330 11620 11340
rect 11788 11330 11844 11340
rect 11340 11284 11396 11294
rect 11340 11190 11396 11228
rect 11900 9828 11956 13356
rect 12236 12964 12292 12974
rect 12236 12870 12292 12908
rect 12348 12290 12404 13580
rect 12796 12964 12852 16044
rect 12796 12898 12852 12908
rect 12908 13972 12964 17052
rect 13132 15652 13188 15662
rect 13132 15538 13188 15596
rect 13132 15486 13134 15538
rect 13186 15486 13188 15538
rect 13132 15474 13188 15486
rect 13020 15428 13076 15438
rect 13020 15334 13076 15372
rect 13020 14530 13076 14542
rect 13020 14478 13022 14530
rect 13074 14478 13076 14530
rect 13020 14308 13076 14478
rect 13020 14242 13076 14252
rect 12572 12740 12628 12750
rect 12908 12740 12964 13916
rect 12572 12738 12964 12740
rect 12572 12686 12574 12738
rect 12626 12686 12964 12738
rect 12572 12684 12964 12686
rect 13244 13746 13300 18172
rect 13692 17668 13748 17678
rect 13692 17574 13748 17612
rect 13356 15314 13412 15326
rect 13356 15262 13358 15314
rect 13410 15262 13412 15314
rect 13356 13860 13412 15262
rect 13804 14756 13860 19516
rect 13916 19122 13972 19740
rect 14028 19458 14084 19964
rect 14028 19406 14030 19458
rect 14082 19406 14084 19458
rect 14028 19394 14084 19406
rect 13916 19070 13918 19122
rect 13970 19070 13972 19122
rect 13916 19058 13972 19070
rect 14140 18004 14196 24332
rect 14476 23268 14532 24892
rect 14700 24834 14756 25228
rect 14700 24782 14702 24834
rect 14754 24782 14756 24834
rect 14588 24610 14644 24622
rect 14588 24558 14590 24610
rect 14642 24558 14644 24610
rect 14588 23604 14644 24558
rect 14588 23538 14644 23548
rect 14700 23378 14756 24782
rect 14700 23326 14702 23378
rect 14754 23326 14756 23378
rect 14700 23314 14756 23326
rect 14588 23268 14644 23278
rect 14252 23212 14420 23268
rect 14476 23266 14644 23268
rect 14476 23214 14590 23266
rect 14642 23214 14644 23266
rect 14476 23212 14644 23214
rect 14252 23154 14308 23212
rect 14252 23102 14254 23154
rect 14306 23102 14308 23154
rect 14252 23090 14308 23102
rect 14364 23156 14420 23212
rect 14588 23202 14644 23212
rect 14364 23100 14532 23156
rect 14364 22932 14420 22942
rect 14364 18452 14420 22876
rect 14140 17948 14308 18004
rect 14140 17780 14196 17790
rect 13916 17108 13972 17118
rect 14140 17108 14196 17724
rect 14252 17220 14308 17948
rect 14364 17666 14420 18396
rect 14364 17614 14366 17666
rect 14418 17614 14420 17666
rect 14364 17602 14420 17614
rect 14476 20132 14532 23100
rect 14588 23044 14644 23054
rect 14588 22484 14644 22988
rect 14588 22370 14644 22428
rect 14700 22930 14756 22942
rect 14700 22878 14702 22930
rect 14754 22878 14756 22930
rect 14700 22596 14756 22878
rect 14812 22932 14868 25342
rect 14924 25394 15092 25396
rect 14924 25342 15038 25394
rect 15090 25342 15092 25394
rect 14924 25340 15092 25342
rect 14924 23044 14980 25340
rect 15036 25330 15092 25340
rect 14924 22978 14980 22988
rect 15036 25172 15092 25182
rect 14812 22866 14868 22876
rect 15036 22708 15092 25116
rect 15036 22642 15092 22652
rect 14700 22482 14756 22540
rect 14700 22430 14702 22482
rect 14754 22430 14756 22482
rect 14700 22418 14756 22430
rect 15036 22482 15092 22494
rect 15036 22430 15038 22482
rect 15090 22430 15092 22482
rect 14588 22318 14590 22370
rect 14642 22318 14644 22370
rect 14588 22306 14644 22318
rect 14924 21812 14980 21822
rect 14924 21718 14980 21756
rect 14812 21586 14868 21598
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14812 21252 14868 21534
rect 15036 21588 15092 22430
rect 15036 21522 15092 21532
rect 15148 21586 15204 21598
rect 15148 21534 15150 21586
rect 15202 21534 15204 21586
rect 14812 21186 14868 21196
rect 15148 21140 15204 21534
rect 15148 21074 15204 21084
rect 14588 20132 14644 20142
rect 14476 20130 14644 20132
rect 14476 20078 14590 20130
rect 14642 20078 14644 20130
rect 14476 20076 14644 20078
rect 14476 17668 14532 20076
rect 14588 20066 14644 20076
rect 15148 19906 15204 19918
rect 15148 19854 15150 19906
rect 15202 19854 15204 19906
rect 15148 19460 15204 19854
rect 15148 19394 15204 19404
rect 15036 19348 15092 19358
rect 14588 18564 14644 18574
rect 14588 18470 14644 18508
rect 14924 18452 14980 18462
rect 14588 17780 14644 17818
rect 14588 17714 14644 17724
rect 14476 17602 14532 17612
rect 14588 17554 14644 17566
rect 14588 17502 14590 17554
rect 14642 17502 14644 17554
rect 14252 17164 14420 17220
rect 13916 17106 14308 17108
rect 13916 17054 13918 17106
rect 13970 17054 14308 17106
rect 13916 17052 14308 17054
rect 13916 17042 13972 17052
rect 14252 16994 14308 17052
rect 14252 16942 14254 16994
rect 14306 16942 14308 16994
rect 14252 16930 14308 16942
rect 14140 16884 14196 16894
rect 14140 16790 14196 16828
rect 14252 16772 14308 16782
rect 13356 13794 13412 13804
rect 13468 14700 13860 14756
rect 14140 16660 14196 16670
rect 13468 14642 13524 14700
rect 13468 14590 13470 14642
rect 13522 14590 13524 14642
rect 13244 13694 13246 13746
rect 13298 13694 13300 13746
rect 12572 12674 12628 12684
rect 12348 12238 12350 12290
rect 12402 12238 12404 12290
rect 12236 11844 12292 11854
rect 12236 11282 12292 11788
rect 12348 11732 12404 12238
rect 12684 12404 12740 12414
rect 12684 12180 12740 12348
rect 12348 11666 12404 11676
rect 12460 12178 12740 12180
rect 12460 12126 12686 12178
rect 12738 12126 12740 12178
rect 12460 12124 12740 12126
rect 12236 11230 12238 11282
rect 12290 11230 12292 11282
rect 12124 10724 12180 10734
rect 12236 10724 12292 11230
rect 12124 10722 12292 10724
rect 12124 10670 12126 10722
rect 12178 10670 12292 10722
rect 12124 10668 12292 10670
rect 12460 11284 12516 12124
rect 12684 12114 12740 12124
rect 12684 11954 12740 11966
rect 12684 11902 12686 11954
rect 12738 11902 12740 11954
rect 12684 11394 12740 11902
rect 12684 11342 12686 11394
rect 12738 11342 12740 11394
rect 12684 11330 12740 11342
rect 13020 11732 13076 11742
rect 12124 10658 12180 10668
rect 12348 10612 12404 10622
rect 12460 10612 12516 11228
rect 12796 11172 12852 11182
rect 12796 11078 12852 11116
rect 12348 10610 12516 10612
rect 12348 10558 12350 10610
rect 12402 10558 12516 10610
rect 12348 10556 12516 10558
rect 13020 10610 13076 11676
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 12348 10546 12404 10556
rect 13020 10546 13076 10558
rect 13244 10052 13300 13694
rect 13468 13636 13524 14590
rect 13580 14420 13636 14430
rect 13580 14326 13636 14364
rect 13468 13570 13524 13580
rect 13804 14084 13860 14094
rect 13692 12964 13748 12974
rect 13692 12870 13748 12908
rect 13580 12852 13636 12862
rect 13580 12758 13636 12796
rect 13356 12738 13412 12750
rect 13356 12686 13358 12738
rect 13410 12686 13412 12738
rect 13356 12404 13412 12686
rect 13356 12338 13412 12348
rect 13692 12068 13748 12078
rect 13244 9986 13300 9996
rect 13468 12012 13692 12068
rect 12012 9828 12068 9838
rect 11900 9772 12012 9828
rect 12012 9762 12068 9772
rect 13468 6916 13524 12012
rect 13692 12002 13748 12012
rect 13804 10836 13860 14028
rect 14140 13748 14196 16604
rect 14252 15876 14308 16716
rect 14364 16436 14420 17164
rect 14476 16884 14532 16894
rect 14476 16790 14532 16828
rect 14588 16772 14644 17502
rect 14588 16706 14644 16716
rect 14700 17556 14756 17566
rect 14700 16994 14756 17500
rect 14812 17108 14868 17118
rect 14924 17108 14980 18396
rect 15036 17780 15092 19292
rect 15260 18676 15316 18686
rect 15372 18676 15428 29260
rect 15484 23604 15540 29484
rect 15484 23266 15540 23548
rect 15484 23214 15486 23266
rect 15538 23214 15540 23266
rect 15484 23202 15540 23214
rect 15596 28756 15652 28766
rect 15596 23268 15652 28700
rect 16380 28756 16436 30044
rect 16604 29876 16660 30270
rect 16716 30212 16772 30222
rect 16716 30118 16772 30156
rect 16604 29810 16660 29820
rect 16380 28532 16436 28700
rect 16604 29652 16660 29662
rect 16492 28532 16548 28542
rect 16380 28530 16548 28532
rect 16380 28478 16494 28530
rect 16546 28478 16548 28530
rect 16380 28476 16548 28478
rect 16492 28466 16548 28476
rect 16604 28532 16660 29596
rect 17052 28756 17108 28766
rect 17052 28662 17108 28700
rect 16604 28530 16884 28532
rect 16604 28478 16606 28530
rect 16658 28478 16884 28530
rect 16604 28476 16884 28478
rect 16604 28466 16660 28476
rect 16268 28418 16324 28430
rect 16268 28366 16270 28418
rect 16322 28366 16324 28418
rect 15820 27860 15876 27870
rect 15820 27766 15876 27804
rect 15708 27746 15764 27758
rect 15708 27694 15710 27746
rect 15762 27694 15764 27746
rect 15708 25732 15764 27694
rect 15932 27076 15988 27086
rect 15932 26982 15988 27020
rect 16156 26852 16212 26862
rect 16156 26758 16212 26796
rect 16268 26402 16324 28366
rect 16492 27858 16548 27870
rect 16492 27806 16494 27858
rect 16546 27806 16548 27858
rect 16268 26350 16270 26402
rect 16322 26350 16324 26402
rect 15708 25666 15764 25676
rect 15820 26068 15876 26078
rect 15820 25618 15876 26012
rect 15820 25566 15822 25618
rect 15874 25566 15876 25618
rect 15820 25554 15876 25566
rect 16156 25508 16212 25518
rect 16268 25508 16324 26350
rect 16380 27634 16436 27646
rect 16380 27582 16382 27634
rect 16434 27582 16436 27634
rect 16380 26180 16436 27582
rect 16492 26516 16548 27806
rect 16492 26450 16548 26460
rect 16604 27076 16660 27086
rect 16380 26114 16436 26124
rect 16492 26068 16548 26078
rect 16492 25974 16548 26012
rect 16604 25618 16660 27020
rect 16716 26516 16772 26526
rect 16716 26068 16772 26460
rect 16828 26292 16884 28476
rect 17052 27636 17108 27646
rect 16940 27076 16996 27086
rect 16940 26962 16996 27020
rect 17052 27074 17108 27580
rect 17052 27022 17054 27074
rect 17106 27022 17108 27074
rect 17052 27010 17108 27022
rect 16940 26910 16942 26962
rect 16994 26910 16996 26962
rect 16940 26898 16996 26910
rect 16828 26236 16996 26292
rect 16828 26068 16884 26078
rect 16716 26066 16884 26068
rect 16716 26014 16830 26066
rect 16882 26014 16884 26066
rect 16716 26012 16884 26014
rect 16828 26002 16884 26012
rect 16604 25566 16606 25618
rect 16658 25566 16660 25618
rect 16604 25554 16660 25566
rect 16156 25506 16324 25508
rect 16156 25454 16158 25506
rect 16210 25454 16324 25506
rect 16156 25452 16324 25454
rect 16940 25506 16996 26236
rect 16940 25454 16942 25506
rect 16994 25454 16996 25506
rect 16156 25442 16212 25452
rect 16940 25442 16996 25454
rect 16716 23604 16772 23614
rect 15596 23174 15652 23212
rect 16156 23268 16212 23278
rect 16156 23174 16212 23212
rect 15820 23156 15876 23166
rect 15820 23154 15988 23156
rect 15820 23102 15822 23154
rect 15874 23102 15988 23154
rect 15820 23100 15988 23102
rect 15820 23090 15876 23100
rect 15708 22596 15764 22606
rect 15708 22502 15764 22540
rect 15484 22484 15540 22494
rect 15484 22390 15540 22428
rect 15708 21586 15764 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15484 21364 15540 21374
rect 15484 20802 15540 21308
rect 15484 20750 15486 20802
rect 15538 20750 15540 20802
rect 15484 20738 15540 20750
rect 15708 21140 15764 21534
rect 15820 21588 15876 21598
rect 15820 21474 15876 21532
rect 15820 21422 15822 21474
rect 15874 21422 15876 21474
rect 15820 21410 15876 21422
rect 15708 20802 15764 21084
rect 15708 20750 15710 20802
rect 15762 20750 15764 20802
rect 15708 20738 15764 20750
rect 15596 20692 15652 20702
rect 15596 20598 15652 20636
rect 15260 18674 15428 18676
rect 15260 18622 15262 18674
rect 15314 18622 15428 18674
rect 15260 18620 15428 18622
rect 15260 18610 15316 18620
rect 15036 17714 15092 17724
rect 15260 17444 15316 17454
rect 14812 17106 14980 17108
rect 14812 17054 14814 17106
rect 14866 17054 14980 17106
rect 14812 17052 14980 17054
rect 15148 17388 15260 17444
rect 14812 17042 14868 17052
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16660 14756 16942
rect 15036 16996 15092 17006
rect 15148 16996 15204 17388
rect 15260 17378 15316 17388
rect 15036 16994 15204 16996
rect 15036 16942 15038 16994
rect 15090 16942 15204 16994
rect 15036 16940 15204 16942
rect 15036 16930 15092 16940
rect 15148 16884 15204 16940
rect 15260 16884 15316 16894
rect 15148 16882 15316 16884
rect 15148 16830 15262 16882
rect 15314 16830 15316 16882
rect 15148 16828 15316 16830
rect 15260 16818 15316 16828
rect 14700 16594 14756 16604
rect 14364 16380 14756 16436
rect 14364 16212 14420 16222
rect 14364 16098 14420 16156
rect 14364 16046 14366 16098
rect 14418 16046 14420 16098
rect 14364 16034 14420 16046
rect 14700 16210 14756 16380
rect 14700 16158 14702 16210
rect 14754 16158 14756 16210
rect 14252 15820 14420 15876
rect 14252 13748 14308 13758
rect 14140 13746 14308 13748
rect 14140 13694 14254 13746
rect 14306 13694 14308 13746
rect 14140 13692 14308 13694
rect 14252 13682 14308 13692
rect 13916 13522 13972 13534
rect 13916 13470 13918 13522
rect 13970 13470 13972 13522
rect 13916 11844 13972 13470
rect 14364 13412 14420 15820
rect 14700 15148 14756 16158
rect 15260 16212 15316 16222
rect 15372 16212 15428 18620
rect 15484 19460 15540 19470
rect 15484 17108 15540 19404
rect 15932 19124 15988 23100
rect 16716 22370 16772 23548
rect 16716 22318 16718 22370
rect 16770 22318 16772 22370
rect 16716 22306 16772 22318
rect 16044 22146 16100 22158
rect 16044 22094 16046 22146
rect 16098 22094 16100 22146
rect 16044 20802 16100 22094
rect 16828 22148 16884 22158
rect 16828 22054 16884 22092
rect 17052 22146 17108 22158
rect 17052 22094 17054 22146
rect 17106 22094 17108 22146
rect 16492 21588 16548 21598
rect 16492 21586 16996 21588
rect 16492 21534 16494 21586
rect 16546 21534 16996 21586
rect 16492 21532 16996 21534
rect 16492 21522 16548 21532
rect 16044 20750 16046 20802
rect 16098 20750 16100 20802
rect 16044 20738 16100 20750
rect 16940 20804 16996 21532
rect 16940 20710 16996 20748
rect 16716 20468 16772 20478
rect 15596 19068 16212 19124
rect 15596 17554 15652 19068
rect 15708 18340 15764 18350
rect 15708 18338 15876 18340
rect 15708 18286 15710 18338
rect 15762 18286 15876 18338
rect 15708 18284 15876 18286
rect 15708 18274 15764 18284
rect 15596 17502 15598 17554
rect 15650 17502 15652 17554
rect 15596 17490 15652 17502
rect 15820 17666 15876 18284
rect 15820 17614 15822 17666
rect 15874 17614 15876 17666
rect 15820 17444 15876 17614
rect 15820 17378 15876 17388
rect 15932 18226 15988 18238
rect 15932 18174 15934 18226
rect 15986 18174 15988 18226
rect 15932 17556 15988 18174
rect 15932 17220 15988 17500
rect 15708 17164 15988 17220
rect 15484 17052 15652 17108
rect 15484 16884 15540 16894
rect 15484 16790 15540 16828
rect 15316 16156 15428 16212
rect 14700 15092 14980 15148
rect 14700 14644 14756 14654
rect 14700 14550 14756 14588
rect 14588 14420 14644 14430
rect 14644 14364 14868 14420
rect 14588 14354 14644 14364
rect 14476 13860 14532 13870
rect 14532 13804 14644 13860
rect 14476 13794 14532 13804
rect 14476 13634 14532 13646
rect 14476 13582 14478 13634
rect 14530 13582 14532 13634
rect 14476 13524 14532 13582
rect 14476 13458 14532 13468
rect 14364 12962 14420 13356
rect 14364 12910 14366 12962
rect 14418 12910 14420 12962
rect 14364 12898 14420 12910
rect 14028 12852 14084 12862
rect 14028 12402 14084 12796
rect 14028 12350 14030 12402
rect 14082 12350 14084 12402
rect 14028 12338 14084 12350
rect 14252 12068 14308 12078
rect 14252 11974 14308 12012
rect 13916 11778 13972 11788
rect 13356 6860 13524 6916
rect 13580 10780 13860 10836
rect 13356 6468 13412 6860
rect 13468 6692 13524 6702
rect 13580 6692 13636 10780
rect 13692 10500 13748 10510
rect 13692 10498 14420 10500
rect 13692 10446 13694 10498
rect 13746 10446 14420 10498
rect 13692 10444 14420 10446
rect 13692 10434 13748 10444
rect 14364 9828 14420 10444
rect 14252 9826 14420 9828
rect 14252 9774 14366 9826
rect 14418 9774 14420 9826
rect 14252 9772 14420 9774
rect 13916 9156 13972 9166
rect 13916 9042 13972 9100
rect 13916 8990 13918 9042
rect 13970 8990 13972 9042
rect 13916 8978 13972 8990
rect 14252 9042 14308 9772
rect 14364 9762 14420 9772
rect 14588 9714 14644 13804
rect 14812 13858 14868 14364
rect 14812 13806 14814 13858
rect 14866 13806 14868 13858
rect 14700 13074 14756 13086
rect 14700 13022 14702 13074
rect 14754 13022 14756 13074
rect 14700 12178 14756 13022
rect 14812 12962 14868 13806
rect 14924 13970 14980 15092
rect 14924 13918 14926 13970
rect 14978 13918 14980 13970
rect 14924 13076 14980 13918
rect 15148 13860 15204 13870
rect 15148 13766 15204 13804
rect 14924 13010 14980 13020
rect 14812 12910 14814 12962
rect 14866 12910 14868 12962
rect 14812 12898 14868 12910
rect 15260 12852 15316 16156
rect 15596 15148 15652 17052
rect 15708 16884 15764 17164
rect 16156 17108 16212 19068
rect 16268 18228 16324 18238
rect 16268 18134 16324 18172
rect 16604 18228 16660 18238
rect 16380 17108 16436 17118
rect 16156 17106 16436 17108
rect 16156 17054 16382 17106
rect 16434 17054 16436 17106
rect 16156 17052 16436 17054
rect 16380 17042 16436 17052
rect 16604 17106 16660 18172
rect 16716 17892 16772 20412
rect 17052 20356 17108 22094
rect 17164 21364 17220 32844
rect 17388 32674 17444 32686
rect 17388 32622 17390 32674
rect 17442 32622 17444 32674
rect 17388 31778 17444 32622
rect 17612 32562 17668 33068
rect 17612 32510 17614 32562
rect 17666 32510 17668 32562
rect 17612 32498 17668 32510
rect 17388 31726 17390 31778
rect 17442 31726 17444 31778
rect 17388 31714 17444 31726
rect 17500 31108 17556 31118
rect 17500 31014 17556 31052
rect 17388 30996 17444 31006
rect 17388 30902 17444 30940
rect 17276 30098 17332 30110
rect 17276 30046 17278 30098
rect 17330 30046 17332 30098
rect 17276 29540 17332 30046
rect 17388 30100 17444 30110
rect 17388 30006 17444 30044
rect 17612 29988 17668 29998
rect 17612 29894 17668 29932
rect 17276 29474 17332 29484
rect 17724 27860 17780 27870
rect 17836 27860 17892 34524
rect 17948 33124 18004 34750
rect 18396 34468 18452 35420
rect 18508 34914 18564 34926
rect 18508 34862 18510 34914
rect 18562 34862 18564 34914
rect 18508 34692 18564 34862
rect 18508 34626 18564 34636
rect 18620 34916 18676 35980
rect 18396 34412 18564 34468
rect 18172 33572 18228 33582
rect 18172 33458 18228 33516
rect 18172 33406 18174 33458
rect 18226 33406 18228 33458
rect 18172 33394 18228 33406
rect 18508 33348 18564 34412
rect 18620 34356 18676 34860
rect 18620 34290 18676 34300
rect 18732 33684 18788 38612
rect 18844 38500 18900 38510
rect 18844 35924 18900 38444
rect 18844 35858 18900 35868
rect 18844 35698 18900 35710
rect 18844 35646 18846 35698
rect 18898 35646 18900 35698
rect 18844 35138 18900 35646
rect 18844 35086 18846 35138
rect 18898 35086 18900 35138
rect 18844 35074 18900 35086
rect 18956 35140 19012 41132
rect 19180 41188 19236 41806
rect 20076 41860 20132 41870
rect 20188 41860 20244 43598
rect 20412 42756 20468 42766
rect 20524 42756 20580 45164
rect 20748 45154 20804 45164
rect 20860 43650 20916 50316
rect 20972 50306 21028 50316
rect 20860 43598 20862 43650
rect 20914 43598 20916 43650
rect 20860 43586 20916 43598
rect 20972 47796 21028 47806
rect 20972 43540 21028 47740
rect 21084 43764 21140 52892
rect 21420 52836 21476 52846
rect 21756 52836 21812 53004
rect 21868 52994 21924 53004
rect 21980 52948 22036 52958
rect 22428 52948 22484 54460
rect 22988 54450 23044 54460
rect 23100 53730 23156 54796
rect 23324 54738 23380 55244
rect 23548 55298 23604 56924
rect 23548 55246 23550 55298
rect 23602 55246 23604 55298
rect 23548 55234 23604 55246
rect 23324 54686 23326 54738
rect 23378 54686 23380 54738
rect 23324 54674 23380 54686
rect 23100 53678 23102 53730
rect 23154 53678 23156 53730
rect 23100 53666 23156 53678
rect 22988 53620 23044 53630
rect 21980 52854 22036 52892
rect 22092 52946 22484 52948
rect 22092 52894 22430 52946
rect 22482 52894 22484 52946
rect 22092 52892 22484 52894
rect 21420 52834 21812 52836
rect 21420 52782 21422 52834
rect 21474 52782 21812 52834
rect 21420 52780 21812 52782
rect 21868 52836 21924 52846
rect 21420 52770 21476 52780
rect 21420 52162 21476 52174
rect 21420 52110 21422 52162
rect 21474 52110 21476 52162
rect 21420 52052 21476 52110
rect 21308 51996 21420 52052
rect 21196 51940 21252 51950
rect 21196 50708 21252 51884
rect 21308 50818 21364 51996
rect 21420 51986 21476 51996
rect 21308 50766 21310 50818
rect 21362 50766 21364 50818
rect 21308 50754 21364 50766
rect 21196 50642 21252 50652
rect 21420 50596 21476 50606
rect 21420 50482 21476 50540
rect 21420 50430 21422 50482
rect 21474 50430 21476 50482
rect 21420 50428 21476 50430
rect 21196 50372 21476 50428
rect 21196 49812 21252 50372
rect 21420 49924 21476 49934
rect 21196 49810 21364 49812
rect 21196 49758 21198 49810
rect 21250 49758 21364 49810
rect 21196 49756 21364 49758
rect 21196 49746 21252 49756
rect 21196 49364 21252 49374
rect 21196 47460 21252 49308
rect 21308 48804 21364 49756
rect 21308 48738 21364 48748
rect 21420 49026 21476 49868
rect 21420 48974 21422 49026
rect 21474 48974 21476 49026
rect 21308 47460 21364 47470
rect 21196 47458 21364 47460
rect 21196 47406 21310 47458
rect 21362 47406 21364 47458
rect 21196 47404 21364 47406
rect 21196 46676 21252 46686
rect 21196 46562 21252 46620
rect 21196 46510 21198 46562
rect 21250 46510 21252 46562
rect 21196 45106 21252 46510
rect 21308 45780 21364 47404
rect 21420 46452 21476 48974
rect 21532 47068 21588 52780
rect 21868 52722 21924 52780
rect 21868 52670 21870 52722
rect 21922 52670 21924 52722
rect 21868 52658 21924 52670
rect 21980 52388 22036 52398
rect 22092 52388 22148 52892
rect 22428 52882 22484 52892
rect 22652 53058 22708 53070
rect 22652 53006 22654 53058
rect 22706 53006 22708 53058
rect 22652 52948 22708 53006
rect 22652 52882 22708 52892
rect 22876 52724 22932 52734
rect 21980 52386 22148 52388
rect 21980 52334 21982 52386
rect 22034 52334 22148 52386
rect 21980 52332 22148 52334
rect 22540 52500 22596 52510
rect 21980 52322 22036 52332
rect 21644 52276 21700 52286
rect 21644 52274 21924 52276
rect 21644 52222 21646 52274
rect 21698 52222 21924 52274
rect 21644 52220 21924 52222
rect 21644 52210 21700 52220
rect 21868 51380 21924 52220
rect 22316 52164 22372 52174
rect 22316 52070 22372 52108
rect 22316 51828 22372 51838
rect 22540 51828 22596 52444
rect 22876 52274 22932 52668
rect 22988 52500 23044 53564
rect 23212 53060 23268 53070
rect 23212 52966 23268 53004
rect 23548 52946 23604 52958
rect 23548 52894 23550 52946
rect 23602 52894 23604 52946
rect 23548 52724 23604 52894
rect 23548 52658 23604 52668
rect 22988 52434 23044 52444
rect 23212 52612 23268 52622
rect 22876 52222 22878 52274
rect 22930 52222 22932 52274
rect 22764 51940 22820 51950
rect 22540 51772 22708 51828
rect 22316 51602 22372 51772
rect 22316 51550 22318 51602
rect 22370 51550 22372 51602
rect 22316 51538 22372 51550
rect 22540 51604 22596 51614
rect 22540 51510 22596 51548
rect 22204 51380 22260 51390
rect 21868 51378 22372 51380
rect 21868 51326 22206 51378
rect 22258 51326 22372 51378
rect 21868 51324 22372 51326
rect 22204 51314 22260 51324
rect 22204 50596 22260 50606
rect 22204 50502 22260 50540
rect 21644 50482 21700 50494
rect 21644 50430 21646 50482
rect 21698 50430 21700 50482
rect 21644 50036 21700 50430
rect 21644 49970 21700 49980
rect 21868 49924 21924 49934
rect 21868 49830 21924 49868
rect 22204 49810 22260 49822
rect 22204 49758 22206 49810
rect 22258 49758 22260 49810
rect 21756 49588 21812 49598
rect 21756 49138 21812 49532
rect 21756 49086 21758 49138
rect 21810 49086 21812 49138
rect 21532 47012 21700 47068
rect 21420 46386 21476 46396
rect 21308 45714 21364 45724
rect 21532 46004 21588 46014
rect 21532 45778 21588 45948
rect 21532 45726 21534 45778
rect 21586 45726 21588 45778
rect 21532 45714 21588 45726
rect 21644 45220 21700 47012
rect 21196 45054 21198 45106
rect 21250 45054 21252 45106
rect 21196 44884 21252 45054
rect 21532 45164 21700 45220
rect 21756 45220 21812 49086
rect 22204 49028 22260 49758
rect 22204 48934 22260 48972
rect 22204 47236 22260 47246
rect 22204 46564 22260 47180
rect 22092 46562 22260 46564
rect 22092 46510 22206 46562
rect 22258 46510 22260 46562
rect 22092 46508 22260 46510
rect 21868 45780 21924 45790
rect 21868 45686 21924 45724
rect 21980 45666 22036 45678
rect 21980 45614 21982 45666
rect 22034 45614 22036 45666
rect 21756 45164 21924 45220
rect 21420 44996 21476 45006
rect 21196 44818 21252 44828
rect 21308 44940 21420 44996
rect 21308 43876 21364 44940
rect 21420 44930 21476 44940
rect 21420 44772 21476 44782
rect 21420 44100 21476 44716
rect 21532 44660 21588 45164
rect 21868 45108 21924 45164
rect 21868 45042 21924 45052
rect 21532 44594 21588 44604
rect 21756 44994 21812 45006
rect 21756 44942 21758 44994
rect 21810 44942 21812 44994
rect 21756 44884 21812 44942
rect 21532 44436 21588 44446
rect 21588 44380 21700 44436
rect 21532 44370 21588 44380
rect 21420 44034 21476 44044
rect 21308 43820 21588 43876
rect 21084 43708 21476 43764
rect 20972 43474 21028 43484
rect 21308 43538 21364 43550
rect 21308 43486 21310 43538
rect 21362 43486 21364 43538
rect 20412 42754 20580 42756
rect 20412 42702 20414 42754
rect 20466 42702 20580 42754
rect 20412 42700 20580 42702
rect 20412 42690 20468 42700
rect 20300 42644 20356 42654
rect 20300 42196 20356 42588
rect 20524 42532 20580 42700
rect 20748 43428 20804 43438
rect 20524 42476 20692 42532
rect 20300 42140 20468 42196
rect 20300 41972 20356 41982
rect 20300 41878 20356 41916
rect 20132 41804 20244 41860
rect 20076 41766 20132 41804
rect 19180 41122 19236 41132
rect 19292 41410 19348 41422
rect 19292 41358 19294 41410
rect 19346 41358 19348 41410
rect 19292 40962 19348 41358
rect 19628 41188 19684 41198
rect 19628 41094 19684 41132
rect 19292 40910 19294 40962
rect 19346 40910 19348 40962
rect 19068 37380 19124 37390
rect 19068 36594 19124 37324
rect 19292 36708 19348 40910
rect 19516 41074 19572 41086
rect 19516 41022 19518 41074
rect 19570 41022 19572 41074
rect 19516 38500 19572 41022
rect 20188 41074 20244 41086
rect 20188 41022 20190 41074
rect 20242 41022 20244 41074
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20188 40404 20244 41022
rect 20412 41074 20468 42140
rect 20636 42194 20692 42476
rect 20636 42142 20638 42194
rect 20690 42142 20692 42194
rect 20636 42130 20692 42142
rect 20412 41022 20414 41074
rect 20466 41022 20468 41074
rect 20412 41010 20468 41022
rect 20636 41076 20692 41086
rect 20188 40338 20244 40348
rect 20300 40292 20356 40302
rect 20300 40290 20580 40292
rect 20300 40238 20302 40290
rect 20354 40238 20580 40290
rect 20300 40236 20580 40238
rect 20300 40226 20356 40236
rect 20412 39394 20468 39406
rect 20412 39342 20414 39394
rect 20466 39342 20468 39394
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20412 38668 20468 39342
rect 19516 38434 19572 38444
rect 20188 38612 20468 38668
rect 19628 38050 19684 38062
rect 19628 37998 19630 38050
rect 19682 37998 19684 38050
rect 19516 37380 19572 37390
rect 19516 37286 19572 37324
rect 19628 37156 19684 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19852 37268 19908 37278
rect 19852 37174 19908 37212
rect 19628 37100 19796 37156
rect 19292 36652 19684 36708
rect 19068 36542 19070 36594
rect 19122 36542 19124 36594
rect 19068 36530 19124 36542
rect 19292 36484 19348 36494
rect 19180 36260 19236 36270
rect 19180 35698 19236 36204
rect 19292 35812 19348 36428
rect 19292 35746 19348 35756
rect 19404 36372 19460 36382
rect 19180 35646 19182 35698
rect 19234 35646 19236 35698
rect 19068 35588 19124 35598
rect 19068 35494 19124 35532
rect 19180 35364 19236 35646
rect 19404 35476 19460 36316
rect 19628 36260 19684 36652
rect 19740 36706 19796 37100
rect 19964 37154 20020 37166
rect 19964 37102 19966 37154
rect 20018 37102 20020 37154
rect 19964 37044 20020 37102
rect 19964 36978 20020 36988
rect 19740 36654 19742 36706
rect 19794 36654 19796 36706
rect 19740 36642 19796 36654
rect 19740 36484 19796 36494
rect 19740 36370 19796 36428
rect 19740 36318 19742 36370
rect 19794 36318 19796 36370
rect 19740 36306 19796 36318
rect 19852 36372 19908 36382
rect 20188 36372 20244 38612
rect 19908 36316 20244 36372
rect 20300 38500 20356 38510
rect 20300 37268 20356 38444
rect 20300 36594 20356 37212
rect 20300 36542 20302 36594
rect 20354 36542 20356 36594
rect 19852 36278 19908 36316
rect 19404 35410 19460 35420
rect 19516 36204 19684 36260
rect 19180 35298 19236 35308
rect 18956 35084 19124 35140
rect 18956 34916 19012 34926
rect 18844 34132 18900 34142
rect 18956 34132 19012 34860
rect 18844 34130 19012 34132
rect 18844 34078 18846 34130
rect 18898 34078 19012 34130
rect 18844 34076 19012 34078
rect 18844 34066 18900 34076
rect 18732 33618 18788 33628
rect 19068 33572 19124 35084
rect 19292 34020 19348 34030
rect 19292 33926 19348 33964
rect 19068 33506 19124 33516
rect 18508 33282 18564 33292
rect 18732 33348 18788 33358
rect 18732 33234 18788 33292
rect 18732 33182 18734 33234
rect 18786 33182 18788 33234
rect 18732 33170 18788 33182
rect 17948 33058 18004 33068
rect 18396 33124 18452 33134
rect 18396 33030 18452 33068
rect 19404 33124 19460 33134
rect 18844 32564 18900 32574
rect 19404 32564 19460 33068
rect 18844 32562 19460 32564
rect 18844 32510 18846 32562
rect 18898 32510 19460 32562
rect 18844 32508 19460 32510
rect 18508 32452 18564 32462
rect 18844 32452 18900 32508
rect 18508 32450 18900 32452
rect 18508 32398 18510 32450
rect 18562 32398 18900 32450
rect 18508 32396 18900 32398
rect 18396 31666 18452 31678
rect 18396 31614 18398 31666
rect 18450 31614 18452 31666
rect 18284 30994 18340 31006
rect 18284 30942 18286 30994
rect 18338 30942 18340 30994
rect 18060 30882 18116 30894
rect 18060 30830 18062 30882
rect 18114 30830 18116 30882
rect 18060 30322 18116 30830
rect 18284 30884 18340 30942
rect 18396 30996 18452 31614
rect 18396 30930 18452 30940
rect 18284 30818 18340 30828
rect 18508 30660 18564 32396
rect 18956 32340 19012 32350
rect 18956 32246 19012 32284
rect 18060 30270 18062 30322
rect 18114 30270 18116 30322
rect 18060 30100 18116 30270
rect 18284 30604 18564 30660
rect 18060 30034 18116 30044
rect 18172 30098 18228 30110
rect 18172 30046 18174 30098
rect 18226 30046 18228 30098
rect 18172 29876 18228 30046
rect 18172 29810 18228 29820
rect 17836 27804 18228 27860
rect 17724 27186 17780 27804
rect 18060 27636 18116 27646
rect 18060 27542 18116 27580
rect 17724 27134 17726 27186
rect 17778 27134 17780 27186
rect 17612 27076 17668 27086
rect 17612 26982 17668 27020
rect 17724 26964 17780 27134
rect 17724 26898 17780 26908
rect 17836 27076 17892 27086
rect 17612 26740 17668 26750
rect 17276 25282 17332 25294
rect 17276 25230 17278 25282
rect 17330 25230 17332 25282
rect 17276 24724 17332 25230
rect 17276 24658 17332 24668
rect 17388 23492 17444 23502
rect 17164 21298 17220 21308
rect 17276 22146 17332 22158
rect 17276 22094 17278 22146
rect 17330 22094 17332 22146
rect 17276 21812 17332 22094
rect 17052 20290 17108 20300
rect 17164 20914 17220 20926
rect 17164 20862 17166 20914
rect 17218 20862 17220 20914
rect 17164 20132 17220 20862
rect 17276 20468 17332 21756
rect 17388 21026 17444 23436
rect 17612 22596 17668 26684
rect 17612 22258 17668 22540
rect 17612 22206 17614 22258
rect 17666 22206 17668 22258
rect 17612 22194 17668 22206
rect 17836 21812 17892 27020
rect 18172 24946 18228 27804
rect 18284 26740 18340 30604
rect 19404 30210 19460 30222
rect 19404 30158 19406 30210
rect 19458 30158 19460 30210
rect 18620 30100 18676 30110
rect 18508 29764 18564 29774
rect 18396 29540 18452 29550
rect 18396 27298 18452 29484
rect 18508 28756 18564 29708
rect 18620 29538 18676 30044
rect 19292 29988 19348 29998
rect 18956 29876 19012 29886
rect 18620 29486 18622 29538
rect 18674 29486 18676 29538
rect 18620 29474 18676 29486
rect 18844 29540 18900 29550
rect 18844 29446 18900 29484
rect 18508 28662 18564 28700
rect 18844 29314 18900 29326
rect 18844 29262 18846 29314
rect 18898 29262 18900 29314
rect 18844 28642 18900 29262
rect 18844 28590 18846 28642
rect 18898 28590 18900 28642
rect 18844 28578 18900 28590
rect 18956 28642 19012 29820
rect 18956 28590 18958 28642
rect 19010 28590 19012 28642
rect 18956 28578 19012 28590
rect 19180 28644 19236 28654
rect 19180 28550 19236 28588
rect 19292 28642 19348 29932
rect 19404 29540 19460 30158
rect 19404 29474 19460 29484
rect 19292 28590 19294 28642
rect 19346 28590 19348 28642
rect 19292 28578 19348 28590
rect 19068 27858 19124 27870
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 19068 27412 19124 27806
rect 19404 27860 19460 27870
rect 19404 27766 19460 27804
rect 19068 27356 19236 27412
rect 18396 27246 18398 27298
rect 18450 27246 18452 27298
rect 18396 27234 18452 27246
rect 19180 27298 19236 27356
rect 19180 27246 19182 27298
rect 19234 27246 19236 27298
rect 19180 27234 19236 27246
rect 19404 27300 19460 27310
rect 19404 27186 19460 27244
rect 19404 27134 19406 27186
rect 19458 27134 19460 27186
rect 19404 27122 19460 27134
rect 19516 26908 19572 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35812 19796 35822
rect 19740 35718 19796 35756
rect 20188 35026 20244 35038
rect 20188 34974 20190 35026
rect 20242 34974 20244 35026
rect 20188 34804 20244 34974
rect 20188 34738 20244 34748
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19964 34132 20020 34142
rect 19628 33572 19684 33582
rect 19628 33478 19684 33516
rect 19964 33570 20020 34076
rect 19964 33518 19966 33570
rect 20018 33518 20020 33570
rect 19964 33506 20020 33518
rect 19628 33236 19684 33246
rect 19628 32786 19684 33180
rect 19852 33124 19908 33162
rect 19852 33058 19908 33068
rect 20300 33124 20356 36542
rect 20412 37154 20468 37166
rect 20412 37102 20414 37154
rect 20466 37102 20468 37154
rect 20412 35812 20468 37102
rect 20412 35364 20468 35756
rect 20412 34914 20468 35308
rect 20412 34862 20414 34914
rect 20466 34862 20468 34914
rect 20412 34850 20468 34862
rect 20524 33236 20580 40236
rect 20636 39060 20692 41020
rect 20748 39506 20804 43372
rect 21308 42868 21364 43486
rect 20972 42812 21364 42868
rect 20972 42644 21028 42812
rect 21420 42756 21476 43708
rect 20972 42194 21028 42588
rect 20972 42142 20974 42194
rect 21026 42142 21028 42194
rect 20972 42130 21028 42142
rect 21084 42700 21476 42756
rect 20972 40404 21028 40414
rect 20972 39732 21028 40348
rect 20972 39666 21028 39676
rect 20748 39454 20750 39506
rect 20802 39454 20804 39506
rect 20748 39442 20804 39454
rect 20636 38994 20692 39004
rect 20748 38276 20804 38286
rect 20748 38182 20804 38220
rect 20860 37266 20916 37278
rect 20860 37214 20862 37266
rect 20914 37214 20916 37266
rect 20860 37044 20916 37214
rect 20860 36978 20916 36988
rect 20972 35924 21028 35934
rect 20972 35830 21028 35868
rect 21084 35700 21140 42700
rect 21420 42530 21476 42542
rect 21420 42478 21422 42530
rect 21474 42478 21476 42530
rect 21420 41860 21476 42478
rect 21532 41972 21588 43820
rect 21532 41878 21588 41916
rect 21308 41746 21364 41758
rect 21308 41694 21310 41746
rect 21362 41694 21364 41746
rect 21308 41410 21364 41694
rect 21308 41358 21310 41410
rect 21362 41358 21364 41410
rect 21308 41346 21364 41358
rect 21420 40964 21476 41804
rect 21644 41636 21700 44380
rect 21756 44324 21812 44828
rect 21756 44268 21924 44324
rect 21756 44100 21812 44110
rect 21756 44006 21812 44044
rect 21868 43876 21924 44268
rect 21196 40962 21476 40964
rect 21196 40910 21422 40962
rect 21474 40910 21476 40962
rect 21196 40908 21476 40910
rect 21196 35812 21252 40908
rect 21420 40898 21476 40908
rect 21532 41580 21700 41636
rect 21756 43820 21924 43876
rect 21980 43988 22036 45614
rect 22092 44772 22148 46508
rect 22204 46498 22260 46508
rect 22316 45892 22372 51324
rect 22652 50428 22708 51772
rect 22764 51602 22820 51884
rect 22876 51828 22932 52222
rect 22876 51762 22932 51772
rect 22764 51550 22766 51602
rect 22818 51550 22820 51602
rect 22764 51538 22820 51550
rect 22204 45890 22372 45892
rect 22204 45838 22318 45890
rect 22370 45838 22372 45890
rect 22204 45836 22372 45838
rect 22204 45220 22260 45836
rect 22316 45826 22372 45836
rect 22428 50372 22708 50428
rect 22764 51380 22820 51390
rect 22428 47346 22484 50372
rect 22428 47294 22430 47346
rect 22482 47294 22484 47346
rect 22204 45154 22260 45164
rect 22204 44996 22260 45006
rect 22204 44902 22260 44940
rect 22092 44716 22260 44772
rect 22092 44436 22148 44446
rect 22092 44322 22148 44380
rect 22092 44270 22094 44322
rect 22146 44270 22148 44322
rect 22092 44258 22148 44270
rect 22204 44100 22260 44716
rect 22428 44660 22484 47294
rect 22652 49138 22708 49150
rect 22652 49086 22654 49138
rect 22706 49086 22708 49138
rect 22652 47572 22708 49086
rect 22652 47068 22708 47516
rect 22540 47012 22708 47068
rect 22540 46004 22596 47012
rect 22652 46564 22708 46574
rect 22652 46470 22708 46508
rect 22764 46228 22820 51324
rect 23212 51266 23268 52556
rect 23436 52388 23492 52398
rect 23436 52276 23492 52332
rect 23436 52274 23716 52276
rect 23436 52222 23438 52274
rect 23490 52222 23716 52274
rect 23436 52220 23716 52222
rect 23436 52210 23492 52220
rect 23660 52162 23716 52220
rect 23660 52110 23662 52162
rect 23714 52110 23716 52162
rect 23660 52098 23716 52110
rect 23212 51214 23214 51266
rect 23266 51214 23268 51266
rect 23212 48914 23268 51214
rect 23436 51268 23492 51278
rect 23436 50708 23492 51212
rect 23436 50706 23716 50708
rect 23436 50654 23438 50706
rect 23490 50654 23716 50706
rect 23436 50652 23716 50654
rect 23436 50642 23492 50652
rect 23660 50594 23716 50652
rect 23660 50542 23662 50594
rect 23714 50542 23716 50594
rect 23660 50530 23716 50542
rect 23772 50428 23828 57036
rect 23884 56866 23940 57820
rect 24108 56980 24164 58380
rect 24220 58322 24276 58940
rect 24556 58436 24612 59164
rect 24668 58436 24724 58446
rect 24556 58434 24724 58436
rect 24556 58382 24670 58434
rect 24722 58382 24724 58434
rect 24556 58380 24724 58382
rect 24668 58370 24724 58380
rect 24220 58270 24222 58322
rect 24274 58270 24276 58322
rect 24220 58258 24276 58270
rect 24444 58324 24500 58334
rect 24444 58230 24500 58268
rect 24444 57876 24500 57886
rect 24444 57782 24500 57820
rect 24556 57650 24612 57662
rect 24556 57598 24558 57650
rect 24610 57598 24612 57650
rect 24108 56914 24164 56924
rect 24220 57092 24276 57102
rect 23884 56814 23886 56866
rect 23938 56814 23940 56866
rect 23884 56802 23940 56814
rect 24108 56754 24164 56766
rect 24108 56702 24110 56754
rect 24162 56702 24164 56754
rect 24108 55186 24164 56702
rect 24108 55134 24110 55186
rect 24162 55134 24164 55186
rect 23996 54516 24052 54526
rect 23884 54514 24052 54516
rect 23884 54462 23998 54514
rect 24050 54462 24052 54514
rect 23884 54460 24052 54462
rect 23884 51604 23940 54460
rect 23996 54450 24052 54460
rect 23884 51510 23940 51548
rect 23996 53732 24052 53742
rect 23996 52834 24052 53676
rect 23996 52782 23998 52834
rect 24050 52782 24052 52834
rect 23548 50372 23828 50428
rect 23436 49812 23492 49822
rect 23436 49718 23492 49756
rect 23324 49476 23380 49486
rect 23324 49026 23380 49420
rect 23324 48974 23326 49026
rect 23378 48974 23380 49026
rect 23324 48962 23380 48974
rect 23212 48862 23214 48914
rect 23266 48862 23268 48914
rect 22652 46004 22708 46014
rect 22540 45948 22652 46004
rect 22652 45938 22708 45948
rect 22764 45892 22820 46172
rect 22876 47404 23044 47460
rect 22876 47124 22932 47404
rect 22988 47402 23044 47404
rect 22988 47350 22990 47402
rect 23042 47350 23044 47402
rect 22988 47338 23044 47350
rect 23100 47346 23156 47358
rect 23100 47294 23102 47346
rect 23154 47294 23156 47346
rect 22988 47236 23044 47246
rect 23100 47236 23156 47294
rect 23044 47180 23156 47236
rect 22988 47170 23044 47180
rect 22876 46116 22932 47068
rect 22988 46788 23044 46798
rect 22988 46694 23044 46732
rect 23100 46786 23156 46798
rect 23100 46734 23102 46786
rect 23154 46734 23156 46786
rect 23100 46676 23156 46734
rect 23100 46610 23156 46620
rect 23212 46228 23268 48862
rect 23548 48132 23604 50372
rect 23772 49700 23828 49710
rect 23660 49698 23828 49700
rect 23660 49646 23774 49698
rect 23826 49646 23828 49698
rect 23660 49644 23828 49646
rect 23660 49476 23716 49644
rect 23772 49634 23828 49644
rect 23996 49700 24052 52782
rect 24108 52612 24164 55134
rect 24108 52546 24164 52556
rect 24220 52388 24276 57036
rect 24444 56308 24500 56318
rect 24444 56214 24500 56252
rect 24556 56082 24612 57598
rect 24668 56196 24724 56206
rect 24780 56196 24836 60844
rect 24892 60788 24948 61294
rect 25228 60900 25284 60910
rect 25284 60844 25396 60900
rect 25228 60806 25284 60844
rect 24892 60722 24948 60732
rect 24892 60004 24948 60014
rect 24892 59910 24948 59948
rect 25340 60002 25396 60844
rect 25340 59950 25342 60002
rect 25394 59950 25396 60002
rect 25340 59938 25396 59950
rect 25116 59892 25172 59902
rect 25116 59890 25284 59892
rect 25116 59838 25118 59890
rect 25170 59838 25284 59890
rect 25116 59836 25284 59838
rect 25116 59826 25172 59836
rect 25228 59444 25284 59836
rect 25452 59780 25508 62132
rect 25564 60788 25620 60798
rect 25564 60694 25620 60732
rect 25676 60002 25732 62860
rect 26460 62020 26516 65996
rect 26796 65986 26852 65996
rect 27132 64036 27188 68796
rect 27916 68516 27972 68526
rect 27356 68514 27972 68516
rect 27356 68462 27918 68514
rect 27970 68462 27972 68514
rect 27356 68460 27972 68462
rect 27356 67842 27412 68460
rect 27916 68450 27972 68460
rect 27356 67790 27358 67842
rect 27410 67790 27412 67842
rect 27244 67618 27300 67630
rect 27244 67566 27246 67618
rect 27298 67566 27300 67618
rect 27244 66836 27300 67566
rect 27356 67228 27412 67790
rect 27916 67618 27972 67630
rect 27916 67566 27918 67618
rect 27970 67566 27972 67618
rect 27356 67172 27860 67228
rect 27356 67060 27412 67172
rect 27356 66994 27412 67004
rect 27692 67058 27748 67070
rect 27692 67006 27694 67058
rect 27746 67006 27748 67058
rect 27692 66948 27748 67006
rect 27692 66882 27748 66892
rect 27356 66836 27412 66846
rect 27244 66780 27356 66836
rect 27356 66386 27412 66780
rect 27356 66334 27358 66386
rect 27410 66334 27412 66386
rect 27356 66322 27412 66334
rect 27804 66050 27860 67172
rect 27916 66948 27972 67566
rect 27916 66882 27972 66892
rect 27804 65998 27806 66050
rect 27858 65998 27860 66050
rect 27804 64820 27860 65998
rect 27804 64754 27860 64764
rect 27132 63980 27972 64036
rect 26684 63922 26740 63934
rect 26684 63870 26686 63922
rect 26738 63870 26740 63922
rect 26572 63810 26628 63822
rect 26572 63758 26574 63810
rect 26626 63758 26628 63810
rect 26572 63700 26628 63758
rect 26684 63812 26740 63870
rect 26740 63756 26964 63812
rect 26684 63746 26740 63756
rect 26572 63364 26628 63644
rect 26572 63308 26740 63364
rect 26572 63140 26628 63150
rect 26572 63046 26628 63084
rect 26460 61954 26516 61964
rect 26684 62242 26740 63308
rect 26908 62468 26964 63756
rect 27692 63810 27748 63822
rect 27692 63758 27694 63810
rect 27746 63758 27748 63810
rect 27692 63700 27748 63758
rect 27692 63634 27748 63644
rect 27020 63364 27076 63374
rect 27020 63270 27076 63308
rect 27356 63140 27412 63150
rect 27356 63046 27412 63084
rect 27580 63140 27636 63150
rect 27580 63138 27748 63140
rect 27580 63086 27582 63138
rect 27634 63086 27748 63138
rect 27580 63084 27748 63086
rect 27580 63074 27636 63084
rect 27020 62468 27076 62478
rect 26908 62466 27076 62468
rect 26908 62414 27022 62466
rect 27074 62414 27076 62466
rect 26908 62412 27076 62414
rect 27020 62402 27076 62412
rect 26684 62190 26686 62242
rect 26738 62190 26740 62242
rect 26684 62132 26740 62190
rect 27692 62188 27748 63084
rect 26684 61796 26740 62076
rect 27244 62132 27300 62142
rect 27244 62038 27300 62076
rect 27580 62130 27636 62142
rect 27692 62132 27860 62188
rect 27580 62078 27582 62130
rect 27634 62078 27636 62130
rect 25676 59950 25678 60002
rect 25730 59950 25732 60002
rect 25676 59938 25732 59950
rect 26348 61740 26740 61796
rect 26796 62020 26852 62030
rect 26348 59780 26404 61740
rect 26460 60004 26516 60014
rect 26460 59910 26516 59948
rect 25452 59724 25956 59780
rect 26348 59724 26628 59780
rect 25564 59556 25620 59566
rect 25340 59444 25396 59454
rect 25564 59444 25620 59500
rect 25228 59442 25396 59444
rect 25228 59390 25342 59442
rect 25394 59390 25396 59442
rect 25228 59388 25396 59390
rect 25340 59378 25396 59388
rect 25452 59442 25620 59444
rect 25452 59390 25566 59442
rect 25618 59390 25620 59442
rect 25452 59388 25620 59390
rect 25004 58212 25060 58222
rect 25004 58118 25060 58156
rect 25228 58100 25284 58110
rect 25228 57204 25284 58044
rect 25452 57876 25508 59388
rect 25564 59378 25620 59388
rect 25676 59218 25732 59230
rect 25676 59166 25678 59218
rect 25730 59166 25732 59218
rect 25564 58548 25620 58558
rect 25564 58210 25620 58492
rect 25676 58436 25732 59166
rect 25900 58548 25956 59724
rect 25900 58482 25956 58492
rect 26124 59108 26180 59118
rect 25676 58370 25732 58380
rect 25788 58434 25844 58446
rect 25788 58382 25790 58434
rect 25842 58382 25844 58434
rect 25788 58324 25844 58382
rect 25788 58258 25844 58268
rect 25564 58158 25566 58210
rect 25618 58158 25620 58210
rect 25564 58100 25620 58158
rect 26124 58210 26180 59052
rect 26236 59106 26292 59118
rect 26236 59054 26238 59106
rect 26290 59054 26292 59106
rect 26236 58884 26292 59054
rect 26236 58828 26516 58884
rect 26348 58660 26404 58670
rect 26236 58604 26348 58660
rect 26236 58434 26292 58604
rect 26348 58594 26404 58604
rect 26236 58382 26238 58434
rect 26290 58382 26292 58434
rect 26236 58370 26292 58382
rect 26348 58434 26404 58446
rect 26348 58382 26350 58434
rect 26402 58382 26404 58434
rect 26124 58158 26126 58210
rect 26178 58158 26180 58210
rect 26124 58146 26180 58158
rect 26348 58212 26404 58382
rect 25564 58034 25620 58044
rect 25564 57876 25620 57886
rect 25452 57874 25620 57876
rect 25452 57822 25566 57874
rect 25618 57822 25620 57874
rect 25452 57820 25620 57822
rect 25564 57810 25620 57820
rect 25788 57876 25844 57886
rect 25788 57874 26180 57876
rect 25788 57822 25790 57874
rect 25842 57822 26180 57874
rect 25788 57820 26180 57822
rect 25788 57810 25844 57820
rect 24668 56194 24836 56196
rect 24668 56142 24670 56194
rect 24722 56142 24836 56194
rect 24668 56140 24836 56142
rect 25116 57148 25284 57204
rect 25452 57650 25508 57662
rect 25452 57598 25454 57650
rect 25506 57598 25508 57650
rect 24668 56130 24724 56140
rect 24556 56030 24558 56082
rect 24610 56030 24612 56082
rect 24556 55748 24612 56030
rect 24556 55692 24948 55748
rect 24892 55412 24948 55692
rect 24668 55300 24724 55310
rect 24332 54628 24388 54638
rect 24332 54626 24500 54628
rect 24332 54574 24334 54626
rect 24386 54574 24500 54626
rect 24332 54572 24500 54574
rect 24332 54562 24388 54572
rect 24444 54180 24500 54572
rect 24444 53058 24500 54124
rect 24668 53618 24724 55244
rect 24668 53566 24670 53618
rect 24722 53566 24724 53618
rect 24668 53554 24724 53566
rect 24780 54068 24836 54078
rect 24780 53170 24836 54012
rect 24892 53730 24948 55356
rect 24892 53678 24894 53730
rect 24946 53678 24948 53730
rect 24892 53666 24948 53678
rect 24780 53118 24782 53170
rect 24834 53118 24836 53170
rect 24780 53106 24836 53118
rect 24444 53006 24446 53058
rect 24498 53006 24500 53058
rect 24444 52994 24500 53006
rect 24556 53060 24612 53070
rect 24612 53004 24724 53060
rect 24556 52966 24612 53004
rect 23996 49634 24052 49644
rect 24108 52332 24276 52388
rect 24444 52724 24500 52734
rect 23660 49410 23716 49420
rect 23660 48244 23716 48254
rect 23716 48188 23828 48244
rect 23660 48150 23716 48188
rect 23548 48066 23604 48076
rect 23772 47570 23828 48188
rect 23996 48242 24052 48254
rect 23996 48190 23998 48242
rect 24050 48190 24052 48242
rect 23772 47518 23774 47570
rect 23826 47518 23828 47570
rect 23772 47506 23828 47518
rect 23884 47572 23940 47582
rect 23436 47460 23492 47470
rect 23324 47236 23380 47246
rect 23324 47142 23380 47180
rect 23324 46900 23380 46910
rect 23436 46900 23492 47404
rect 23884 47012 23940 47516
rect 23996 47236 24052 48190
rect 23996 47170 24052 47180
rect 23324 46898 23492 46900
rect 23324 46846 23326 46898
rect 23378 46846 23492 46898
rect 23324 46844 23492 46846
rect 23660 46956 23940 47012
rect 23324 46834 23380 46844
rect 23100 46172 23268 46228
rect 23548 46674 23604 46686
rect 23548 46622 23550 46674
rect 23602 46622 23604 46674
rect 22876 46060 23044 46116
rect 22876 45892 22932 45902
rect 22764 45890 22932 45892
rect 22764 45838 22878 45890
rect 22930 45838 22932 45890
rect 22764 45836 22932 45838
rect 22876 45780 22932 45836
rect 22876 45714 22932 45724
rect 22428 44594 22484 44604
rect 22652 45108 22708 45118
rect 22428 44212 22484 44222
rect 22428 44118 22484 44156
rect 22204 44034 22260 44044
rect 21532 40516 21588 41580
rect 21756 41410 21812 43820
rect 21868 43540 21924 43550
rect 21980 43540 22036 43932
rect 21868 43538 22036 43540
rect 21868 43486 21870 43538
rect 21922 43486 22036 43538
rect 21868 43484 22036 43486
rect 22092 43650 22148 43662
rect 22092 43598 22094 43650
rect 22146 43598 22148 43650
rect 21868 43474 21924 43484
rect 22092 42980 22148 43598
rect 22092 42914 22148 42924
rect 22428 42754 22484 42766
rect 22428 42702 22430 42754
rect 22482 42702 22484 42754
rect 22092 42532 22148 42542
rect 22428 42532 22484 42702
rect 22092 42530 22484 42532
rect 22092 42478 22094 42530
rect 22146 42478 22484 42530
rect 22092 42476 22484 42478
rect 21980 41972 22036 41982
rect 21756 41358 21758 41410
rect 21810 41358 21812 41410
rect 21756 41346 21812 41358
rect 21868 41748 21924 41758
rect 21756 41188 21812 41198
rect 21644 41076 21700 41086
rect 21644 40626 21700 41020
rect 21644 40574 21646 40626
rect 21698 40574 21700 40626
rect 21644 40562 21700 40574
rect 21532 40422 21588 40460
rect 21420 40404 21476 40414
rect 21420 40292 21476 40348
rect 21420 40236 21588 40292
rect 21532 40180 21588 40236
rect 21644 40180 21700 40190
rect 21532 40178 21700 40180
rect 21532 40126 21646 40178
rect 21698 40126 21700 40178
rect 21532 40124 21700 40126
rect 21644 40114 21700 40124
rect 21532 39956 21588 39966
rect 21308 39396 21364 39406
rect 21308 39394 21476 39396
rect 21308 39342 21310 39394
rect 21362 39342 21476 39394
rect 21308 39340 21476 39342
rect 21308 39330 21364 39340
rect 21308 39060 21364 39070
rect 21308 38966 21364 39004
rect 21420 36484 21476 39340
rect 21420 36418 21476 36428
rect 21196 35756 21476 35812
rect 20972 35644 21140 35700
rect 20636 35588 20692 35598
rect 20636 35138 20692 35532
rect 20636 35086 20638 35138
rect 20690 35086 20692 35138
rect 20636 35074 20692 35086
rect 20972 34244 21028 35644
rect 21308 35588 21364 35598
rect 21308 35494 21364 35532
rect 21420 35476 21476 35756
rect 21420 35410 21476 35420
rect 21196 35364 21252 35374
rect 21252 35308 21364 35364
rect 21196 35298 21252 35308
rect 21308 35252 21364 35308
rect 21308 35196 21476 35252
rect 21308 34804 21364 34814
rect 21308 34710 21364 34748
rect 21420 34802 21476 35196
rect 21420 34750 21422 34802
rect 21474 34750 21476 34802
rect 21420 34738 21476 34750
rect 21420 34356 21476 34366
rect 21420 34262 21476 34300
rect 20972 34188 21252 34244
rect 20524 33170 20580 33180
rect 21084 34020 21140 34030
rect 20300 33058 20356 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 21084 32900 21140 33964
rect 19836 32890 20100 32900
rect 19628 32734 19630 32786
rect 19682 32734 19684 32786
rect 19628 32722 19684 32734
rect 20524 32844 21140 32900
rect 19964 32676 20020 32686
rect 19964 32582 20020 32620
rect 20412 32676 20468 32686
rect 20412 32582 20468 32620
rect 20524 32674 20580 32844
rect 21084 32786 21140 32844
rect 21084 32734 21086 32786
rect 21138 32734 21140 32786
rect 21084 32722 21140 32734
rect 20524 32622 20526 32674
rect 20578 32622 20580 32674
rect 20524 32610 20580 32622
rect 20972 32676 21028 32686
rect 20748 32564 20804 32574
rect 20412 32340 20468 32350
rect 20300 32338 20468 32340
rect 20300 32286 20414 32338
rect 20466 32286 20468 32338
rect 20300 32284 20468 32286
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 30996 20132 31006
rect 20076 30902 20132 30940
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20188 29652 20244 29662
rect 19852 28756 19908 28766
rect 19852 28642 19908 28700
rect 19852 28590 19854 28642
rect 19906 28590 19908 28642
rect 19852 28578 19908 28590
rect 20188 28754 20244 29596
rect 20188 28702 20190 28754
rect 20242 28702 20244 28754
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 28084 20244 28702
rect 19964 28028 20244 28084
rect 19852 27746 19908 27758
rect 19852 27694 19854 27746
rect 19906 27694 19908 27746
rect 19852 27298 19908 27694
rect 19852 27246 19854 27298
rect 19906 27246 19908 27298
rect 19852 27234 19908 27246
rect 19964 27186 20020 28028
rect 19964 27134 19966 27186
rect 20018 27134 20020 27186
rect 19964 27122 20020 27134
rect 18284 26674 18340 26684
rect 18508 26852 18564 26862
rect 18284 26180 18340 26190
rect 18284 25508 18340 26124
rect 18508 26178 18564 26796
rect 19404 26852 19572 26908
rect 20300 26908 20356 32284
rect 20412 32274 20468 32284
rect 20748 31106 20804 32508
rect 20748 31054 20750 31106
rect 20802 31054 20804 31106
rect 20748 31042 20804 31054
rect 20524 30884 20580 30894
rect 20524 30790 20580 30828
rect 20748 30322 20804 30334
rect 20748 30270 20750 30322
rect 20802 30270 20804 30322
rect 20748 30212 20804 30270
rect 20748 30146 20804 30156
rect 20636 29652 20692 29662
rect 20412 28644 20468 28654
rect 20412 28642 20580 28644
rect 20412 28590 20414 28642
rect 20466 28590 20580 28642
rect 20412 28588 20580 28590
rect 20412 28578 20468 28588
rect 20524 28084 20580 28588
rect 20524 28018 20580 28028
rect 20412 27970 20468 27982
rect 20412 27918 20414 27970
rect 20466 27918 20468 27970
rect 20412 27300 20468 27918
rect 20636 27970 20692 29596
rect 20636 27918 20638 27970
rect 20690 27918 20692 27970
rect 20636 27906 20692 27918
rect 20524 27748 20580 27758
rect 20524 27654 20580 27692
rect 20412 27234 20468 27244
rect 20636 27300 20692 27310
rect 20636 27186 20692 27244
rect 20636 27134 20638 27186
rect 20690 27134 20692 27186
rect 20636 27122 20692 27134
rect 20748 27076 20804 27086
rect 20748 26908 20804 27020
rect 20300 26852 20580 26908
rect 20748 26852 20916 26908
rect 19404 26628 19460 26852
rect 18508 26126 18510 26178
rect 18562 26126 18564 26178
rect 18284 25414 18340 25452
rect 18396 25618 18452 25630
rect 18396 25566 18398 25618
rect 18450 25566 18452 25618
rect 18172 24894 18174 24946
rect 18226 24894 18228 24946
rect 18060 24724 18116 24734
rect 17948 21812 18004 21822
rect 17836 21756 17948 21812
rect 17724 21700 17780 21710
rect 17724 21698 17892 21700
rect 17724 21646 17726 21698
rect 17778 21646 17892 21698
rect 17724 21644 17892 21646
rect 17724 21634 17780 21644
rect 17612 21588 17668 21598
rect 17612 21494 17668 21532
rect 17724 21364 17780 21374
rect 17724 21270 17780 21308
rect 17388 20974 17390 21026
rect 17442 20974 17444 21026
rect 17388 20962 17444 20974
rect 17836 20916 17892 21644
rect 17948 21252 18004 21756
rect 18060 21588 18116 24668
rect 18172 22372 18228 24894
rect 18396 24946 18452 25566
rect 18508 25284 18564 26126
rect 18844 26572 19460 26628
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18732 25844 18788 25854
rect 18508 25218 18564 25228
rect 18620 25788 18732 25844
rect 18396 24894 18398 24946
rect 18450 24894 18452 24946
rect 18396 24882 18452 24894
rect 18508 23828 18564 23838
rect 18172 22370 18452 22372
rect 18172 22318 18174 22370
rect 18226 22318 18452 22370
rect 18172 22316 18452 22318
rect 18172 22148 18228 22316
rect 18172 22082 18228 22092
rect 18284 21812 18340 21822
rect 18284 21698 18340 21756
rect 18396 21810 18452 22316
rect 18396 21758 18398 21810
rect 18450 21758 18452 21810
rect 18396 21746 18452 21758
rect 18508 22146 18564 23772
rect 18620 22260 18676 25788
rect 18732 25778 18788 25788
rect 18732 25620 18788 25630
rect 18732 24498 18788 25564
rect 18732 24446 18734 24498
rect 18786 24446 18788 24498
rect 18732 23492 18788 24446
rect 18732 23426 18788 23436
rect 18844 22372 18900 26572
rect 18956 26402 19012 26414
rect 18956 26350 18958 26402
rect 19010 26350 19012 26402
rect 18956 25396 19012 26350
rect 20188 26290 20244 26302
rect 20188 26238 20190 26290
rect 20242 26238 20244 26290
rect 19068 25396 19124 25406
rect 18956 25394 19124 25396
rect 18956 25342 19070 25394
rect 19122 25342 19124 25394
rect 18956 25340 19124 25342
rect 20188 25396 20244 26238
rect 20412 25396 20468 25406
rect 20188 25394 20468 25396
rect 20188 25342 20414 25394
rect 20466 25342 20468 25394
rect 20188 25340 20468 25342
rect 19068 25284 19124 25340
rect 20412 25330 20468 25340
rect 20076 25284 20132 25294
rect 19068 25228 19572 25284
rect 18956 25172 19012 25182
rect 18956 24946 19012 25116
rect 18956 24894 18958 24946
rect 19010 24894 19012 24946
rect 18956 24882 19012 24894
rect 19516 24836 19572 25228
rect 20132 25228 20244 25284
rect 20076 25218 20132 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 25228
rect 20076 24892 20244 24948
rect 19628 24836 19684 24846
rect 19516 24834 19684 24836
rect 19516 24782 19630 24834
rect 19682 24782 19684 24834
rect 19516 24780 19684 24782
rect 19628 24770 19684 24780
rect 19964 24836 20020 24846
rect 19404 24722 19460 24734
rect 19404 24670 19406 24722
rect 19458 24670 19460 24722
rect 19068 24612 19124 24622
rect 19404 24612 19460 24670
rect 19068 24610 19460 24612
rect 19068 24558 19070 24610
rect 19122 24558 19460 24610
rect 19068 24556 19460 24558
rect 19852 24610 19908 24622
rect 19852 24558 19854 24610
rect 19906 24558 19908 24610
rect 19068 24546 19124 24556
rect 19292 23716 19348 23726
rect 19292 23266 19348 23660
rect 19852 23716 19908 24558
rect 19964 23826 20020 24780
rect 20076 24722 20132 24892
rect 20076 24670 20078 24722
rect 20130 24670 20132 24722
rect 20076 24658 20132 24670
rect 20300 24724 20356 24734
rect 20300 24630 20356 24668
rect 19964 23774 19966 23826
rect 20018 23774 20020 23826
rect 19964 23762 20020 23774
rect 20188 23828 20244 23838
rect 20188 23734 20244 23772
rect 19852 23650 19908 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19292 23214 19294 23266
rect 19346 23214 19348 23266
rect 19292 23202 19348 23214
rect 20300 23042 20356 23054
rect 20300 22990 20302 23042
rect 20354 22990 20356 23042
rect 19404 22708 19460 22718
rect 19404 22482 19460 22652
rect 20188 22708 20244 22718
rect 19404 22430 19406 22482
rect 19458 22430 19460 22482
rect 19404 22418 19460 22430
rect 19740 22484 19796 22494
rect 19740 22390 19796 22428
rect 18844 22316 19124 22372
rect 18732 22260 18788 22270
rect 18620 22204 18732 22260
rect 18732 22194 18788 22204
rect 18508 22094 18510 22146
rect 18562 22094 18564 22146
rect 18284 21646 18286 21698
rect 18338 21646 18340 21698
rect 18284 21634 18340 21646
rect 18060 21522 18116 21532
rect 17948 21186 18004 21196
rect 17836 20850 17892 20860
rect 17276 20402 17332 20412
rect 17724 20804 17780 20814
rect 17724 20242 17780 20748
rect 17724 20190 17726 20242
rect 17778 20190 17780 20242
rect 17724 20178 17780 20190
rect 17164 18564 17220 20076
rect 17948 20132 18004 20142
rect 17948 20038 18004 20076
rect 17276 20020 17332 20030
rect 17276 19926 17332 19964
rect 17164 18498 17220 18508
rect 17836 19906 17892 19918
rect 17836 19854 17838 19906
rect 17890 19854 17892 19906
rect 17836 18452 17892 19854
rect 18508 19796 18564 22094
rect 18844 22146 18900 22158
rect 18844 22094 18846 22146
rect 18898 22094 18900 22146
rect 18844 21924 18900 22094
rect 18844 21858 18900 21868
rect 18620 21588 18676 21598
rect 18620 21586 19012 21588
rect 18620 21534 18622 21586
rect 18674 21534 19012 21586
rect 18620 21532 19012 21534
rect 18620 21522 18676 21532
rect 18956 20914 19012 21532
rect 18956 20862 18958 20914
rect 19010 20862 19012 20914
rect 18956 20850 19012 20862
rect 19068 20692 19124 22316
rect 20076 22370 20132 22382
rect 20076 22318 20078 22370
rect 20130 22318 20132 22370
rect 20076 22148 20132 22318
rect 20076 22082 20132 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21810 20244 22652
rect 20300 22482 20356 22990
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20300 22418 20356 22430
rect 20524 22372 20580 26852
rect 20860 26402 20916 26852
rect 20860 26350 20862 26402
rect 20914 26350 20916 26402
rect 20860 26338 20916 26350
rect 20748 25620 20804 25630
rect 20636 25508 20692 25518
rect 20636 23938 20692 25452
rect 20748 25506 20804 25564
rect 20748 25454 20750 25506
rect 20802 25454 20804 25506
rect 20748 25442 20804 25454
rect 20972 25060 21028 32620
rect 21196 32564 21252 34188
rect 21532 33460 21588 39900
rect 21756 39730 21812 41132
rect 21756 39678 21758 39730
rect 21810 39678 21812 39730
rect 21756 39666 21812 39678
rect 21868 40516 21924 41692
rect 21980 41298 22036 41916
rect 22092 41636 22148 42476
rect 22316 41972 22372 41982
rect 22316 41860 22372 41916
rect 22652 41972 22708 45052
rect 22988 44324 23044 46060
rect 23100 44996 23156 46172
rect 23548 45892 23604 46622
rect 23548 45826 23604 45836
rect 23212 45778 23268 45790
rect 23212 45726 23214 45778
rect 23266 45726 23268 45778
rect 23212 45108 23268 45726
rect 23436 45780 23492 45790
rect 23436 45686 23492 45724
rect 23324 45666 23380 45678
rect 23660 45668 23716 46956
rect 23884 46898 23940 46956
rect 23884 46846 23886 46898
rect 23938 46846 23940 46898
rect 23884 46834 23940 46846
rect 23324 45614 23326 45666
rect 23378 45614 23380 45666
rect 23324 45332 23380 45614
rect 23324 45266 23380 45276
rect 23548 45612 23716 45668
rect 23772 46788 23828 46798
rect 23324 45108 23380 45118
rect 23212 45106 23380 45108
rect 23212 45054 23326 45106
rect 23378 45054 23380 45106
rect 23212 45052 23380 45054
rect 23100 44940 23268 44996
rect 23100 44548 23156 44558
rect 23100 44454 23156 44492
rect 22988 44268 23156 44324
rect 22764 44210 22820 44222
rect 22764 44158 22766 44210
rect 22818 44158 22820 44210
rect 22764 43988 22820 44158
rect 22988 44100 23044 44110
rect 22988 44006 23044 44044
rect 22764 43922 22820 43932
rect 22652 41906 22708 41916
rect 22764 43652 22820 43662
rect 22092 41570 22148 41580
rect 22204 41858 22372 41860
rect 22204 41806 22318 41858
rect 22370 41806 22372 41858
rect 22204 41804 22372 41806
rect 21980 41246 21982 41298
rect 22034 41246 22036 41298
rect 21980 41188 22036 41246
rect 21980 41122 22036 41132
rect 22092 40516 22148 40526
rect 21868 40514 22148 40516
rect 21868 40462 22094 40514
rect 22146 40462 22148 40514
rect 21868 40460 22148 40462
rect 21868 39058 21924 40460
rect 22092 40450 22148 40460
rect 21868 39006 21870 39058
rect 21922 39006 21924 39058
rect 21868 38994 21924 39006
rect 21980 37266 22036 37278
rect 21980 37214 21982 37266
rect 22034 37214 22036 37266
rect 21868 37044 21924 37054
rect 21644 35700 21700 35710
rect 21644 34914 21700 35644
rect 21756 35700 21812 35710
rect 21868 35700 21924 36988
rect 21756 35698 21924 35700
rect 21756 35646 21758 35698
rect 21810 35646 21924 35698
rect 21756 35644 21924 35646
rect 21756 35634 21812 35644
rect 21644 34862 21646 34914
rect 21698 34862 21700 34914
rect 21644 34850 21700 34862
rect 21756 35476 21812 35486
rect 21532 33404 21700 33460
rect 21308 33348 21364 33358
rect 21308 33254 21364 33292
rect 21532 33236 21588 33246
rect 21532 33142 21588 33180
rect 21084 32508 21252 32564
rect 21308 33124 21364 33134
rect 21084 28756 21140 32508
rect 21196 30994 21252 31006
rect 21196 30942 21198 30994
rect 21250 30942 21252 30994
rect 21196 30212 21252 30942
rect 21196 30146 21252 30156
rect 21084 28690 21140 28700
rect 21196 25284 21252 25294
rect 21196 25190 21252 25228
rect 20636 23886 20638 23938
rect 20690 23886 20692 23938
rect 20636 23874 20692 23886
rect 20748 25004 21028 25060
rect 20748 23548 20804 25004
rect 21308 24948 21364 33068
rect 21420 31106 21476 31118
rect 21420 31054 21422 31106
rect 21474 31054 21476 31106
rect 21420 30210 21476 31054
rect 21420 30158 21422 30210
rect 21474 30158 21476 30210
rect 21420 30146 21476 30158
rect 21644 29652 21700 33404
rect 21756 31668 21812 35420
rect 21980 35252 22036 37214
rect 22204 36706 22260 41804
rect 22316 41794 22372 41804
rect 22764 41858 22820 43596
rect 23100 42196 23156 44268
rect 23212 42642 23268 44940
rect 23324 43988 23380 45052
rect 23548 44772 23604 45612
rect 23660 45218 23716 45230
rect 23660 45166 23662 45218
rect 23714 45166 23716 45218
rect 23660 44996 23716 45166
rect 23660 44930 23716 44940
rect 23548 44716 23716 44772
rect 23548 44436 23604 44446
rect 23548 44342 23604 44380
rect 23324 43922 23380 43932
rect 23548 44100 23604 44110
rect 23212 42590 23214 42642
rect 23266 42590 23268 42642
rect 23212 42578 23268 42590
rect 23548 42196 23604 44044
rect 23660 43204 23716 44716
rect 23772 44324 23828 46732
rect 23884 45892 23940 45902
rect 23884 45798 23940 45836
rect 23996 44436 24052 44446
rect 23884 44324 23940 44334
rect 23772 44322 23940 44324
rect 23772 44270 23886 44322
rect 23938 44270 23940 44322
rect 23772 44268 23940 44270
rect 23884 44212 23940 44268
rect 23772 43876 23828 43886
rect 23772 43650 23828 43820
rect 23772 43598 23774 43650
rect 23826 43598 23828 43650
rect 23772 43586 23828 43598
rect 23884 43652 23940 44156
rect 23996 44210 24052 44380
rect 23996 44158 23998 44210
rect 24050 44158 24052 44210
rect 23996 44146 24052 44158
rect 24108 44100 24164 52332
rect 24444 52052 24500 52668
rect 24668 52164 24724 53004
rect 25116 52948 25172 57148
rect 25452 57092 25508 57598
rect 26012 57650 26068 57662
rect 26012 57598 26014 57650
rect 26066 57598 26068 57650
rect 25452 57036 25732 57092
rect 25228 56980 25284 56990
rect 25228 56194 25284 56924
rect 25452 56866 25508 56878
rect 25452 56814 25454 56866
rect 25506 56814 25508 56866
rect 25340 56420 25396 56430
rect 25340 56306 25396 56364
rect 25340 56254 25342 56306
rect 25394 56254 25396 56306
rect 25340 56242 25396 56254
rect 25228 56142 25230 56194
rect 25282 56142 25284 56194
rect 25228 56130 25284 56142
rect 25452 55300 25508 56814
rect 25676 56868 25732 57036
rect 25452 55206 25508 55244
rect 25564 56082 25620 56094
rect 25564 56030 25566 56082
rect 25618 56030 25620 56082
rect 25564 55188 25620 56030
rect 25564 55122 25620 55132
rect 25340 55076 25396 55086
rect 25396 55020 25508 55076
rect 25340 55010 25396 55020
rect 25452 54516 25508 55020
rect 25564 54516 25620 54526
rect 25452 54514 25620 54516
rect 25452 54462 25566 54514
rect 25618 54462 25620 54514
rect 25452 54460 25620 54462
rect 25564 54450 25620 54460
rect 25340 54404 25396 54414
rect 25340 54402 25508 54404
rect 25340 54350 25342 54402
rect 25394 54350 25508 54402
rect 25340 54348 25508 54350
rect 25340 54338 25396 54348
rect 25452 53620 25508 54348
rect 25676 53732 25732 56812
rect 26012 55410 26068 57598
rect 26124 57652 26180 57820
rect 26236 57652 26292 57662
rect 26124 57650 26292 57652
rect 26124 57598 26238 57650
rect 26290 57598 26292 57650
rect 26124 57596 26292 57598
rect 26236 57586 26292 57596
rect 26124 56644 26180 56682
rect 26124 56578 26180 56588
rect 26124 56420 26180 56430
rect 26124 55972 26180 56364
rect 26348 55972 26404 58156
rect 26460 56868 26516 58828
rect 26460 56802 26516 56812
rect 26460 56644 26516 56654
rect 26460 56194 26516 56588
rect 26460 56142 26462 56194
rect 26514 56142 26516 56194
rect 26460 56130 26516 56142
rect 26124 55878 26180 55916
rect 26236 55916 26404 55972
rect 26012 55358 26014 55410
rect 26066 55358 26068 55410
rect 26012 55346 26068 55358
rect 26124 55188 26180 55198
rect 26124 54628 26180 55132
rect 26124 54562 26180 54572
rect 26236 54626 26292 55916
rect 26572 55860 26628 59724
rect 26236 54574 26238 54626
rect 26290 54574 26292 54626
rect 25788 54516 25844 54526
rect 25788 54422 25844 54460
rect 26012 54514 26068 54526
rect 26012 54462 26014 54514
rect 26066 54462 26068 54514
rect 26012 54292 26068 54462
rect 26236 54516 26292 54574
rect 26236 54450 26292 54460
rect 26348 55804 26628 55860
rect 26012 54226 26068 54236
rect 25676 53666 25732 53676
rect 25900 53730 25956 53742
rect 26236 53732 26292 53742
rect 25900 53678 25902 53730
rect 25954 53678 25956 53730
rect 25452 53554 25508 53564
rect 25340 53508 25396 53518
rect 25340 53414 25396 53452
rect 25676 53060 25732 53070
rect 24668 52098 24724 52108
rect 24780 52892 25172 52948
rect 25340 53058 25732 53060
rect 25340 53006 25678 53058
rect 25730 53006 25732 53058
rect 25340 53004 25732 53006
rect 24444 51986 24500 51996
rect 24220 51604 24276 51614
rect 24220 50428 24276 51548
rect 24220 50372 24500 50428
rect 24332 48916 24388 48926
rect 24332 48466 24388 48860
rect 24332 48414 24334 48466
rect 24386 48414 24388 48466
rect 24332 48402 24388 48414
rect 24444 48468 24500 50372
rect 24668 49700 24724 49710
rect 24668 49140 24724 49644
rect 24668 49074 24724 49084
rect 24444 48412 24724 48468
rect 24332 48242 24388 48254
rect 24332 48190 24334 48242
rect 24386 48190 24388 48242
rect 24332 47458 24388 48190
rect 24556 48242 24612 48254
rect 24556 48190 24558 48242
rect 24610 48190 24612 48242
rect 24556 48132 24612 48190
rect 24556 47572 24612 48076
rect 24556 47506 24612 47516
rect 24332 47406 24334 47458
rect 24386 47406 24388 47458
rect 24332 47394 24388 47406
rect 24668 47458 24724 48412
rect 24668 47406 24670 47458
rect 24722 47406 24724 47458
rect 24220 47236 24276 47246
rect 24556 47236 24612 47246
rect 24220 47234 24612 47236
rect 24220 47182 24222 47234
rect 24274 47182 24558 47234
rect 24610 47182 24612 47234
rect 24220 47180 24612 47182
rect 24220 47170 24276 47180
rect 24220 46788 24276 46798
rect 24220 46694 24276 46732
rect 24332 46786 24388 46798
rect 24332 46734 24334 46786
rect 24386 46734 24388 46786
rect 24332 46116 24388 46734
rect 24444 46452 24500 47180
rect 24556 47170 24612 47180
rect 24556 46676 24612 46686
rect 24556 46582 24612 46620
rect 24444 46396 24612 46452
rect 24332 46050 24388 46060
rect 24444 45892 24500 45902
rect 24444 45798 24500 45836
rect 24444 45220 24500 45230
rect 24444 44882 24500 45164
rect 24444 44830 24446 44882
rect 24498 44830 24500 44882
rect 24444 44818 24500 44830
rect 24108 44034 24164 44044
rect 24220 44098 24276 44110
rect 24220 44046 24222 44098
rect 24274 44046 24276 44098
rect 24108 43876 24164 43886
rect 23996 43652 24052 43662
rect 23884 43650 24052 43652
rect 23884 43598 23998 43650
rect 24050 43598 24052 43650
rect 23884 43596 24052 43598
rect 23996 43586 24052 43596
rect 24108 43650 24164 43820
rect 24108 43598 24110 43650
rect 24162 43598 24164 43650
rect 24108 43586 24164 43598
rect 24220 43652 24276 44046
rect 24220 43586 24276 43596
rect 24332 43538 24388 43550
rect 24332 43486 24334 43538
rect 24386 43486 24388 43538
rect 23660 43148 23940 43204
rect 23100 42140 23492 42196
rect 23548 42140 23828 42196
rect 22988 41972 23044 41982
rect 23212 41972 23268 41982
rect 23044 41970 23268 41972
rect 23044 41918 23214 41970
rect 23266 41918 23268 41970
rect 23044 41916 23268 41918
rect 23436 41972 23492 42140
rect 23436 41916 23604 41972
rect 22988 41906 23044 41916
rect 23212 41906 23268 41916
rect 22764 41806 22766 41858
rect 22818 41806 22820 41858
rect 22764 41748 22820 41806
rect 22764 41682 22820 41692
rect 22428 41410 22484 41422
rect 22428 41358 22430 41410
rect 22482 41358 22484 41410
rect 22428 41076 22484 41358
rect 22428 40982 22484 41020
rect 23436 41188 23492 41198
rect 22876 40964 22932 40974
rect 22932 40908 23156 40964
rect 22876 40870 22932 40908
rect 22428 40852 22484 40862
rect 22316 40796 22428 40852
rect 22316 39620 22372 40796
rect 22428 40786 22484 40796
rect 22428 40572 22932 40628
rect 22428 40402 22484 40572
rect 22428 40350 22430 40402
rect 22482 40350 22484 40402
rect 22428 40338 22484 40350
rect 22652 40404 22708 40414
rect 22652 40310 22708 40348
rect 22540 40290 22596 40302
rect 22540 40238 22542 40290
rect 22594 40238 22596 40290
rect 22428 39620 22484 39630
rect 22316 39618 22484 39620
rect 22316 39566 22430 39618
rect 22482 39566 22484 39618
rect 22316 39564 22484 39566
rect 22540 39620 22596 40238
rect 22876 39956 22932 40572
rect 23100 40626 23156 40908
rect 23100 40574 23102 40626
rect 23154 40574 23156 40626
rect 23100 40562 23156 40574
rect 22988 40516 23044 40526
rect 22988 40422 23044 40460
rect 23324 40516 23380 40526
rect 23324 40422 23380 40460
rect 23436 40180 23492 41132
rect 23548 40852 23604 41916
rect 23660 41970 23716 41982
rect 23660 41918 23662 41970
rect 23714 41918 23716 41970
rect 23660 41748 23716 41918
rect 23660 40964 23716 41692
rect 23772 41300 23828 42140
rect 23884 41636 23940 43148
rect 24108 42754 24164 42766
rect 24108 42702 24110 42754
rect 24162 42702 24164 42754
rect 24108 41858 24164 42702
rect 24108 41806 24110 41858
rect 24162 41806 24164 41858
rect 24108 41794 24164 41806
rect 24220 42082 24276 42094
rect 24220 42030 24222 42082
rect 24274 42030 24276 42082
rect 24220 41860 24276 42030
rect 24332 41972 24388 43486
rect 24332 41906 24388 41916
rect 24444 42980 24500 42990
rect 24220 41794 24276 41804
rect 23884 41580 24388 41636
rect 23772 41234 23828 41244
rect 23660 40898 23716 40908
rect 23884 41076 23940 41086
rect 23548 40514 23604 40796
rect 23660 40628 23716 40638
rect 23884 40628 23940 41020
rect 24220 40628 24276 40638
rect 23660 40626 24276 40628
rect 23660 40574 23662 40626
rect 23714 40574 24222 40626
rect 24274 40574 24276 40626
rect 23660 40572 24276 40574
rect 23660 40562 23716 40572
rect 24220 40562 24276 40572
rect 23548 40462 23550 40514
rect 23602 40462 23604 40514
rect 23548 40450 23604 40462
rect 23660 40180 23716 40190
rect 23996 40180 24052 40190
rect 23436 40124 23604 40180
rect 23548 39956 23604 40124
rect 23660 40086 23716 40124
rect 23772 40178 24052 40180
rect 23772 40126 23998 40178
rect 24050 40126 24052 40178
rect 23772 40124 24052 40126
rect 22876 39900 23156 39956
rect 23100 39842 23156 39900
rect 23100 39790 23102 39842
rect 23154 39790 23156 39842
rect 23100 39778 23156 39790
rect 23436 39900 23604 39956
rect 23212 39620 23268 39630
rect 22540 39564 23044 39620
rect 22428 39554 22484 39564
rect 22540 39394 22596 39406
rect 22540 39342 22542 39394
rect 22594 39342 22596 39394
rect 22316 39060 22372 39070
rect 22540 39060 22596 39342
rect 22372 39004 22596 39060
rect 22764 39394 22820 39406
rect 22764 39342 22766 39394
rect 22818 39342 22820 39394
rect 22316 38966 22372 39004
rect 22764 38836 22820 39342
rect 22764 38770 22820 38780
rect 22988 38668 23044 39564
rect 23212 39526 23268 39564
rect 23100 39394 23156 39406
rect 23100 39342 23102 39394
rect 23154 39342 23156 39394
rect 23100 39060 23156 39342
rect 23212 39060 23268 39070
rect 23100 39058 23268 39060
rect 23100 39006 23214 39058
rect 23266 39006 23268 39058
rect 23100 39004 23268 39006
rect 22204 36654 22206 36706
rect 22258 36654 22260 36706
rect 21868 35196 22036 35252
rect 22092 35364 22148 35374
rect 21868 34804 21924 35196
rect 21980 34916 22036 34926
rect 21980 34822 22036 34860
rect 21868 34738 21924 34748
rect 22092 34244 22148 35308
rect 22204 34916 22260 36654
rect 22428 38612 23044 38668
rect 22316 36596 22372 36606
rect 22316 36502 22372 36540
rect 22316 34916 22372 34926
rect 22204 34914 22372 34916
rect 22204 34862 22318 34914
rect 22370 34862 22372 34914
rect 22204 34860 22372 34862
rect 22204 34356 22260 34860
rect 22316 34850 22372 34860
rect 22204 34290 22260 34300
rect 21868 34242 22148 34244
rect 21868 34190 22094 34242
rect 22146 34190 22148 34242
rect 21868 34188 22148 34190
rect 21868 32788 21924 34188
rect 22092 34178 22148 34188
rect 22316 34018 22372 34030
rect 22316 33966 22318 34018
rect 22370 33966 22372 34018
rect 21980 33236 22036 33246
rect 21980 33142 22036 33180
rect 22092 32788 22148 32798
rect 21868 32786 22148 32788
rect 21868 32734 22094 32786
rect 22146 32734 22148 32786
rect 21868 32732 22148 32734
rect 22092 32722 22148 32732
rect 21868 32564 21924 32574
rect 21868 32470 21924 32508
rect 21980 32450 22036 32462
rect 21980 32398 21982 32450
rect 22034 32398 22036 32450
rect 21980 31780 22036 32398
rect 22092 31780 22148 31790
rect 21980 31778 22148 31780
rect 21980 31726 22094 31778
rect 22146 31726 22148 31778
rect 21980 31724 22148 31726
rect 22092 31714 22148 31724
rect 21756 31612 21924 31668
rect 21756 31444 21812 31454
rect 21756 30098 21812 31388
rect 21868 31332 21924 31612
rect 22316 31556 22372 33966
rect 22316 31490 22372 31500
rect 21868 31266 21924 31276
rect 21756 30046 21758 30098
rect 21810 30046 21812 30098
rect 21756 30034 21812 30046
rect 21644 29586 21700 29596
rect 21868 29988 21924 29998
rect 21756 29538 21812 29550
rect 21756 29486 21758 29538
rect 21810 29486 21812 29538
rect 21532 28644 21588 28654
rect 21532 28550 21588 28588
rect 21644 28532 21700 28542
rect 21532 27972 21588 27982
rect 21532 27878 21588 27916
rect 21644 27188 21700 28476
rect 21756 27860 21812 29486
rect 21868 28084 21924 29932
rect 22428 29540 22484 38612
rect 22652 37380 22708 37390
rect 23212 37380 23268 39004
rect 22652 37286 22708 37324
rect 22988 37324 23268 37380
rect 22652 36708 22708 36718
rect 22652 36594 22708 36652
rect 22652 36542 22654 36594
rect 22706 36542 22708 36594
rect 22652 36530 22708 36542
rect 22764 35924 22820 35934
rect 22764 34914 22820 35868
rect 22764 34862 22766 34914
rect 22818 34862 22820 34914
rect 22764 34850 22820 34862
rect 22988 34916 23044 37324
rect 23436 37268 23492 39900
rect 23548 39620 23604 39630
rect 23548 39526 23604 39564
rect 23660 39508 23716 39518
rect 23772 39508 23828 40124
rect 23996 40114 24052 40124
rect 23884 39676 24276 39732
rect 23884 39618 23940 39676
rect 23884 39566 23886 39618
rect 23938 39566 23940 39618
rect 23884 39554 23940 39566
rect 24220 39618 24276 39676
rect 24220 39566 24222 39618
rect 24274 39566 24276 39618
rect 24220 39554 24276 39566
rect 23660 39506 23828 39508
rect 23660 39454 23662 39506
rect 23714 39454 23828 39506
rect 23660 39452 23828 39454
rect 23548 38836 23604 38846
rect 23548 38742 23604 38780
rect 23212 37212 23492 37268
rect 23100 36706 23156 36718
rect 23100 36654 23102 36706
rect 23154 36654 23156 36706
rect 23100 36596 23156 36654
rect 23100 36502 23156 36540
rect 22988 34850 23044 34860
rect 23100 35364 23156 35374
rect 22540 32562 22596 32574
rect 22540 32510 22542 32562
rect 22594 32510 22596 32562
rect 22540 31780 22596 32510
rect 22764 32564 22820 32574
rect 22764 32470 22820 32508
rect 23100 32562 23156 35308
rect 23212 32900 23268 37212
rect 23436 36372 23492 36382
rect 23660 36372 23716 39452
rect 23996 38946 24052 38958
rect 23996 38894 23998 38946
rect 24050 38894 24052 38946
rect 23996 38388 24052 38894
rect 24332 38948 24388 41580
rect 24444 41186 24500 42924
rect 24556 42420 24612 46396
rect 24668 45444 24724 47406
rect 24668 45378 24724 45388
rect 24780 45332 24836 52892
rect 25340 52388 25396 53004
rect 25676 52994 25732 53004
rect 25788 53058 25844 53070
rect 25788 53006 25790 53058
rect 25842 53006 25844 53058
rect 25452 52834 25508 52846
rect 25452 52782 25454 52834
rect 25506 52782 25508 52834
rect 25452 52724 25508 52782
rect 25788 52724 25844 53006
rect 25900 52836 25956 53678
rect 26124 53730 26292 53732
rect 26124 53678 26238 53730
rect 26290 53678 26292 53730
rect 26124 53676 26292 53678
rect 26012 53060 26068 53070
rect 26124 53060 26180 53676
rect 26236 53666 26292 53676
rect 26236 53508 26292 53518
rect 26236 53414 26292 53452
rect 26012 53058 26180 53060
rect 26012 53006 26014 53058
rect 26066 53006 26180 53058
rect 26012 53004 26180 53006
rect 26012 52994 26068 53004
rect 25900 52770 25956 52780
rect 25452 52668 25844 52724
rect 25340 52332 25508 52388
rect 25004 52162 25060 52174
rect 25004 52110 25006 52162
rect 25058 52110 25060 52162
rect 25004 51940 25060 52110
rect 24892 51380 24948 51390
rect 24892 47012 24948 51324
rect 25004 50594 25060 51884
rect 25004 50542 25006 50594
rect 25058 50542 25060 50594
rect 25004 50530 25060 50542
rect 25340 52162 25396 52174
rect 25340 52110 25342 52162
rect 25394 52110 25396 52162
rect 25340 52052 25396 52110
rect 25340 50594 25396 51996
rect 25452 51604 25508 52332
rect 25788 52164 25844 52668
rect 26236 52724 26292 52734
rect 25788 52108 26068 52164
rect 25452 51538 25508 51548
rect 25788 51940 25844 51950
rect 25340 50542 25342 50594
rect 25394 50542 25396 50594
rect 25340 50530 25396 50542
rect 25788 51378 25844 51884
rect 25788 51326 25790 51378
rect 25842 51326 25844 51378
rect 25788 50260 25844 51326
rect 25788 50194 25844 50204
rect 25900 50484 25956 50494
rect 25340 50036 25396 50046
rect 25228 49924 25284 49934
rect 25340 49924 25396 49980
rect 25564 50036 25620 50046
rect 25900 50036 25956 50428
rect 26012 50428 26068 52108
rect 26236 51940 26292 52668
rect 26236 51874 26292 51884
rect 26236 50820 26292 50830
rect 26012 50372 26180 50428
rect 25564 50034 25956 50036
rect 25564 49982 25566 50034
rect 25618 49982 25956 50034
rect 25564 49980 25956 49982
rect 25564 49970 25620 49980
rect 25228 49922 25396 49924
rect 25228 49870 25230 49922
rect 25282 49870 25396 49922
rect 25228 49868 25396 49870
rect 25900 49922 25956 49980
rect 25900 49870 25902 49922
rect 25954 49870 25956 49922
rect 25228 49026 25284 49868
rect 25900 49858 25956 49870
rect 26012 49922 26068 49934
rect 26012 49870 26014 49922
rect 26066 49870 26068 49922
rect 25228 48974 25230 49026
rect 25282 48974 25284 49026
rect 25228 48962 25284 48974
rect 25340 49700 25396 49710
rect 25340 48466 25396 49644
rect 26012 49364 26068 49870
rect 26124 49924 26180 50372
rect 26236 50034 26292 50764
rect 26236 49982 26238 50034
rect 26290 49982 26292 50034
rect 26236 49970 26292 49982
rect 26124 49858 26180 49868
rect 26012 49028 26068 49308
rect 26012 48962 26068 48972
rect 26348 48916 26404 55804
rect 26796 55748 26852 61964
rect 27132 61684 27188 61694
rect 27188 61628 27524 61684
rect 27132 61590 27188 61628
rect 27468 61570 27524 61628
rect 27468 61518 27470 61570
rect 27522 61518 27524 61570
rect 27468 61506 27524 61518
rect 27132 59220 27188 59230
rect 27132 59218 27412 59220
rect 27132 59166 27134 59218
rect 27186 59166 27412 59218
rect 27132 59164 27412 59166
rect 27132 59154 27188 59164
rect 26908 58660 26964 58670
rect 26908 58566 26964 58604
rect 27020 58436 27076 58446
rect 27020 58322 27076 58380
rect 27020 58270 27022 58322
rect 27074 58270 27076 58322
rect 26908 58210 26964 58222
rect 26908 58158 26910 58210
rect 26962 58158 26964 58210
rect 26908 57428 26964 58158
rect 26908 57362 26964 57372
rect 26460 55692 26852 55748
rect 26460 50428 26516 55692
rect 27020 54964 27076 58270
rect 27356 57092 27412 59164
rect 27244 57036 27412 57092
rect 27244 55188 27300 57036
rect 27580 56980 27636 62078
rect 27804 61346 27860 62132
rect 27804 61294 27806 61346
rect 27858 61294 27860 61346
rect 27804 60676 27860 61294
rect 27804 60610 27860 60620
rect 27804 59108 27860 59118
rect 27804 59014 27860 59052
rect 27916 57092 27972 63980
rect 28028 63140 28084 63150
rect 28028 62914 28084 63084
rect 28028 62862 28030 62914
rect 28082 62862 28084 62914
rect 28028 62468 28084 62862
rect 28028 62374 28084 62412
rect 28140 62188 28196 71820
rect 28252 70532 28308 73950
rect 28588 74002 28644 74732
rect 28812 74786 28868 76414
rect 28812 74734 28814 74786
rect 28866 74734 28868 74786
rect 28812 74722 28868 74734
rect 29148 76468 29204 76478
rect 29148 74786 29204 76412
rect 29260 76354 29316 76636
rect 30380 76690 30436 77196
rect 30380 76638 30382 76690
rect 30434 76638 30436 76690
rect 30380 76626 30436 76638
rect 31164 76692 31220 79200
rect 31164 76626 31220 76636
rect 32620 76692 32676 76702
rect 32620 76598 32676 76636
rect 31164 76468 31220 76478
rect 31164 76374 31220 76412
rect 32396 76468 32452 76478
rect 29260 76302 29262 76354
rect 29314 76302 29316 76354
rect 29260 76290 29316 76302
rect 29260 75684 29316 75694
rect 29260 75590 29316 75628
rect 29596 75684 29652 75694
rect 29148 74734 29150 74786
rect 29202 74734 29204 74786
rect 29148 74722 29204 74734
rect 29596 74900 29652 75628
rect 31500 75684 31556 75694
rect 31500 75590 31556 75628
rect 31948 75684 32004 75694
rect 29596 74116 29652 74844
rect 31948 74898 32004 75628
rect 31948 74846 31950 74898
rect 32002 74846 32004 74898
rect 31948 74834 32004 74846
rect 31276 74788 31332 74798
rect 31276 74694 31332 74732
rect 32396 74226 32452 76412
rect 32956 76356 33012 79200
rect 34748 77364 34804 79200
rect 36540 77364 36596 79200
rect 34748 77308 35140 77364
rect 36540 77308 36932 77364
rect 35084 76580 35140 77308
rect 36876 76692 36932 77308
rect 38332 77028 38388 79200
rect 38332 76972 38836 77028
rect 33404 76468 33460 76478
rect 33404 76374 33460 76412
rect 34748 76468 34804 76478
rect 32956 76300 33348 76356
rect 32620 75572 32676 75582
rect 32620 75570 33124 75572
rect 32620 75518 32622 75570
rect 32674 75518 33124 75570
rect 32620 75516 33124 75518
rect 32620 75506 32676 75516
rect 32396 74174 32398 74226
rect 32450 74174 32452 74226
rect 32396 74162 32452 74174
rect 28588 73950 28590 74002
rect 28642 73950 28644 74002
rect 28588 73938 28644 73950
rect 29148 74114 29652 74116
rect 29148 74062 29598 74114
rect 29650 74062 29652 74114
rect 29148 74060 29652 74062
rect 29148 73554 29204 74060
rect 29596 74050 29652 74060
rect 30268 74004 30324 74014
rect 30268 74002 30660 74004
rect 30268 73950 30270 74002
rect 30322 73950 30660 74002
rect 30268 73948 30660 73950
rect 30268 73938 30324 73948
rect 29148 73502 29150 73554
rect 29202 73502 29204 73554
rect 29148 73490 29204 73502
rect 30604 73554 30660 73948
rect 33068 74002 33124 75516
rect 33292 75124 33348 76300
rect 34300 76242 34356 76254
rect 34300 76190 34302 76242
rect 34354 76190 34356 76242
rect 33516 75124 33572 75134
rect 33292 75122 33572 75124
rect 33292 75070 33294 75122
rect 33346 75070 33518 75122
rect 33570 75070 33572 75122
rect 33292 75068 33572 75070
rect 33292 75058 33348 75068
rect 33516 75058 33572 75068
rect 33964 74786 34020 74798
rect 33964 74734 33966 74786
rect 34018 74734 34020 74786
rect 33068 73950 33070 74002
rect 33122 73950 33124 74002
rect 33068 73938 33124 73950
rect 33292 74114 33348 74126
rect 33292 74062 33294 74114
rect 33346 74062 33348 74114
rect 30604 73502 30606 73554
rect 30658 73502 30660 73554
rect 30604 73490 30660 73502
rect 30828 73332 30884 73342
rect 30492 73330 30884 73332
rect 30492 73278 30830 73330
rect 30882 73278 30884 73330
rect 30492 73276 30884 73278
rect 28476 73218 28532 73230
rect 28476 73166 28478 73218
rect 28530 73166 28532 73218
rect 28364 72100 28420 72110
rect 28364 71652 28420 72044
rect 28476 71876 28532 73166
rect 30492 72658 30548 73276
rect 30828 73266 30884 73276
rect 30492 72606 30494 72658
rect 30546 72606 30548 72658
rect 30492 72594 30548 72606
rect 33180 72660 33236 72670
rect 33292 72660 33348 74062
rect 33964 73668 34020 74734
rect 33964 73602 34020 73612
rect 33180 72658 33348 72660
rect 33180 72606 33182 72658
rect 33234 72606 33348 72658
rect 33180 72604 33348 72606
rect 34300 72660 34356 76190
rect 34748 75794 34804 76412
rect 35084 76466 35140 76524
rect 36092 76580 36148 76590
rect 36092 76486 36148 76524
rect 35084 76414 35086 76466
rect 35138 76414 35140 76466
rect 35084 76402 35140 76414
rect 36876 76468 36932 76636
rect 37548 76692 37604 76702
rect 37548 76598 37604 76636
rect 36988 76468 37044 76478
rect 36876 76466 37044 76468
rect 36876 76414 36990 76466
rect 37042 76414 37044 76466
rect 36876 76412 37044 76414
rect 36988 76402 37044 76412
rect 38780 76468 38836 76972
rect 40124 76580 40180 79200
rect 41916 77252 41972 79200
rect 41916 77196 42420 77252
rect 42364 76692 42420 77196
rect 43708 77026 43764 79200
rect 43708 76974 43710 77026
rect 43762 76974 43764 77026
rect 43708 76962 43764 76974
rect 44268 77026 44324 77038
rect 44268 76974 44270 77026
rect 44322 76974 44324 77026
rect 40124 76514 40180 76524
rect 40796 76580 40852 76590
rect 38780 76466 39172 76468
rect 38780 76414 38782 76466
rect 38834 76414 39172 76466
rect 38780 76412 39172 76414
rect 38780 76402 38836 76412
rect 36540 76354 36596 76366
rect 36540 76302 36542 76354
rect 36594 76302 36596 76354
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 34748 75742 34750 75794
rect 34802 75742 34804 75794
rect 34748 75730 34804 75742
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 36540 73220 36596 76302
rect 38332 76354 38388 76366
rect 38332 76302 38334 76354
rect 38386 76302 38388 76354
rect 38332 75908 38388 76302
rect 38332 75842 38388 75852
rect 39116 75794 39172 76412
rect 40796 76466 40852 76524
rect 41468 76580 41524 76590
rect 41468 76486 41524 76524
rect 40796 76414 40798 76466
rect 40850 76414 40852 76466
rect 40796 76402 40852 76414
rect 42364 76466 42420 76636
rect 42924 76692 42980 76702
rect 42924 76598 42980 76636
rect 44268 76690 44324 76974
rect 44268 76638 44270 76690
rect 44322 76638 44324 76690
rect 44268 76626 44324 76638
rect 44716 77026 44772 77038
rect 44716 76974 44718 77026
rect 44770 76974 44772 77026
rect 44716 76690 44772 76974
rect 45500 77026 45556 79200
rect 45500 76974 45502 77026
rect 45554 76974 45556 77026
rect 45500 76962 45556 76974
rect 46060 77026 46116 77038
rect 46060 76974 46062 77026
rect 46114 76974 46116 77026
rect 44716 76638 44718 76690
rect 44770 76638 44772 76690
rect 44716 76626 44772 76638
rect 46060 76690 46116 76974
rect 46060 76638 46062 76690
rect 46114 76638 46116 76690
rect 46060 76626 46116 76638
rect 46508 77026 46564 77038
rect 46508 76974 46510 77026
rect 46562 76974 46564 77026
rect 46508 76690 46564 76974
rect 46508 76638 46510 76690
rect 46562 76638 46564 76690
rect 46508 76626 46564 76638
rect 42364 76414 42366 76466
rect 42418 76414 42420 76466
rect 42364 76402 42420 76414
rect 43708 76468 43764 76478
rect 43708 76374 43764 76412
rect 42028 76354 42084 76366
rect 42028 76302 42030 76354
rect 42082 76302 42084 76354
rect 39116 75742 39118 75794
rect 39170 75742 39172 75794
rect 39116 75730 39172 75742
rect 40012 76242 40068 76254
rect 40012 76190 40014 76242
rect 40066 76190 40068 76242
rect 40012 75796 40068 76190
rect 40012 75730 40068 75740
rect 36540 73154 36596 73164
rect 40348 74004 40404 74014
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 33180 72594 33236 72604
rect 34300 72594 34356 72604
rect 31164 72546 31220 72558
rect 31164 72494 31166 72546
rect 31218 72494 31220 72546
rect 31164 71988 31220 72494
rect 31164 71894 31220 71932
rect 31388 72546 31444 72558
rect 31388 72494 31390 72546
rect 31442 72494 31444 72546
rect 28476 71810 28532 71820
rect 29820 71876 29876 71886
rect 28364 71596 28532 71652
rect 28252 70466 28308 70476
rect 28476 70306 28532 71596
rect 29484 70866 29540 70878
rect 29484 70814 29486 70866
rect 29538 70814 29540 70866
rect 28700 70756 28756 70766
rect 29484 70756 29540 70814
rect 28700 70754 29540 70756
rect 28700 70702 28702 70754
rect 28754 70702 29540 70754
rect 28700 70700 29540 70702
rect 28700 70690 28756 70700
rect 29148 70532 29204 70542
rect 28476 70254 28478 70306
rect 28530 70254 28532 70306
rect 28476 70242 28532 70254
rect 29036 70420 29092 70430
rect 29036 70194 29092 70364
rect 29036 70142 29038 70194
rect 29090 70142 29092 70194
rect 29036 70130 29092 70142
rect 29148 67954 29204 70476
rect 29148 67902 29150 67954
rect 29202 67902 29204 67954
rect 29148 67890 29204 67902
rect 29372 70082 29428 70094
rect 29372 70030 29374 70082
rect 29426 70030 29428 70082
rect 29372 69634 29428 70030
rect 29372 69582 29374 69634
rect 29426 69582 29428 69634
rect 28364 67618 28420 67630
rect 28364 67566 28366 67618
rect 28418 67566 28420 67618
rect 28364 67228 28420 67566
rect 28364 67172 28644 67228
rect 28364 67060 28420 67070
rect 28364 66966 28420 67004
rect 28588 66836 28644 67172
rect 29260 67172 29316 67182
rect 28588 66770 28644 66780
rect 29148 67058 29204 67070
rect 29148 67006 29150 67058
rect 29202 67006 29204 67058
rect 29148 66052 29204 67006
rect 29148 65986 29204 65996
rect 29260 64036 29316 67116
rect 29372 66834 29428 69582
rect 29484 67228 29540 70700
rect 29596 70644 29652 70654
rect 29596 69298 29652 70588
rect 29820 69860 29876 71820
rect 30492 71876 30548 71886
rect 30492 71782 30548 71820
rect 31388 71874 31444 72494
rect 32508 72546 32564 72558
rect 32508 72494 32510 72546
rect 32562 72494 32564 72546
rect 32508 72324 32564 72494
rect 33068 72546 33124 72558
rect 33068 72494 33070 72546
rect 33122 72494 33124 72546
rect 33068 72436 33124 72494
rect 33852 72546 33908 72558
rect 34076 72548 34132 72558
rect 33852 72494 33854 72546
rect 33906 72494 33908 72546
rect 33516 72436 33572 72446
rect 32172 72268 32564 72324
rect 32620 72434 33572 72436
rect 32620 72382 33518 72434
rect 33570 72382 33572 72434
rect 32620 72380 33572 72382
rect 31948 71988 32004 71998
rect 31948 71894 32004 71932
rect 31388 71822 31390 71874
rect 31442 71822 31444 71874
rect 30044 71762 30100 71774
rect 30044 71710 30046 71762
rect 30098 71710 30100 71762
rect 29932 70980 29988 70990
rect 29932 70886 29988 70924
rect 30044 70306 30100 71710
rect 30716 71762 30772 71774
rect 30716 71710 30718 71762
rect 30770 71710 30772 71762
rect 30268 71650 30324 71662
rect 30268 71598 30270 71650
rect 30322 71598 30324 71650
rect 30268 70644 30324 71598
rect 30716 71652 30772 71710
rect 31052 71652 31108 71662
rect 30716 71650 31108 71652
rect 30716 71598 31054 71650
rect 31106 71598 31108 71650
rect 30716 71596 31108 71598
rect 31052 71586 31108 71596
rect 31388 71090 31444 71822
rect 31388 71038 31390 71090
rect 31442 71038 31444 71090
rect 31388 71026 31444 71038
rect 32172 71874 32228 72268
rect 32620 72212 32676 72380
rect 33516 72370 33572 72380
rect 33852 72324 33908 72494
rect 33852 72258 33908 72268
rect 33964 72546 34132 72548
rect 33964 72494 34078 72546
rect 34130 72494 34132 72546
rect 33964 72492 34132 72494
rect 32172 71822 32174 71874
rect 32226 71822 32228 71874
rect 30268 70578 30324 70588
rect 30492 70980 30548 70990
rect 30044 70254 30046 70306
rect 30098 70254 30100 70306
rect 30044 70242 30100 70254
rect 30492 70194 30548 70924
rect 30492 70142 30494 70194
rect 30546 70142 30548 70194
rect 30492 70130 30548 70142
rect 30940 70978 30996 70990
rect 30940 70926 30942 70978
rect 30994 70926 30996 70978
rect 30940 70868 30996 70926
rect 30940 70194 30996 70812
rect 30940 70142 30942 70194
rect 30994 70142 30996 70194
rect 30940 70130 30996 70142
rect 29820 69794 29876 69804
rect 29708 69524 29764 69534
rect 29708 69522 30212 69524
rect 29708 69470 29710 69522
rect 29762 69470 30212 69522
rect 29708 69468 30212 69470
rect 29708 69458 29764 69468
rect 29596 69246 29598 69298
rect 29650 69246 29652 69298
rect 29596 69234 29652 69246
rect 29820 67844 29876 67854
rect 29820 67750 29876 67788
rect 30044 67842 30100 67854
rect 30044 67790 30046 67842
rect 30098 67790 30100 67842
rect 29484 67172 29652 67228
rect 29596 67106 29652 67116
rect 29372 66782 29374 66834
rect 29426 66782 29428 66834
rect 29372 66770 29428 66782
rect 29484 67060 29540 67070
rect 29484 66276 29540 67004
rect 29484 66182 29540 66220
rect 29596 66836 29652 66846
rect 29596 66052 29652 66780
rect 29036 63980 29316 64036
rect 29484 65996 29652 66052
rect 29820 66276 29876 66286
rect 28924 63810 28980 63822
rect 28924 63758 28926 63810
rect 28978 63758 28980 63810
rect 28924 63028 28980 63758
rect 28924 62962 28980 62972
rect 28476 62916 28532 62926
rect 27916 57026 27972 57036
rect 28028 62132 28196 62188
rect 28364 62914 28532 62916
rect 28364 62862 28478 62914
rect 28530 62862 28532 62914
rect 28364 62860 28532 62862
rect 27468 56924 27636 56980
rect 27244 55122 27300 55132
rect 27356 56866 27412 56878
rect 27356 56814 27358 56866
rect 27410 56814 27412 56866
rect 27356 55298 27412 56814
rect 27468 55860 27524 56924
rect 27580 56754 27636 56766
rect 27580 56702 27582 56754
rect 27634 56702 27636 56754
rect 27580 56644 27636 56702
rect 27916 56644 27972 56654
rect 27580 56578 27636 56588
rect 27692 56642 27972 56644
rect 27692 56590 27918 56642
rect 27970 56590 27972 56642
rect 27692 56588 27972 56590
rect 27692 56082 27748 56588
rect 27916 56578 27972 56588
rect 28028 56420 28084 62132
rect 28364 60564 28420 62860
rect 28476 62850 28532 62860
rect 28924 60676 28980 60686
rect 28924 60564 28980 60620
rect 28364 60508 28980 60564
rect 28140 58548 28196 58558
rect 28140 57650 28196 58492
rect 28140 57598 28142 57650
rect 28194 57598 28196 57650
rect 28140 57586 28196 57598
rect 28364 57762 28420 57774
rect 28364 57710 28366 57762
rect 28418 57710 28420 57762
rect 28364 57652 28420 57710
rect 28364 57586 28420 57596
rect 28140 57428 28196 57438
rect 28140 56754 28196 57372
rect 28252 56868 28308 56878
rect 28252 56774 28308 56812
rect 28476 56756 28532 60508
rect 28588 60116 28644 60126
rect 28588 60114 28868 60116
rect 28588 60062 28590 60114
rect 28642 60062 28868 60114
rect 28588 60060 28868 60062
rect 28588 60050 28644 60060
rect 28140 56702 28142 56754
rect 28194 56702 28196 56754
rect 28140 56690 28196 56702
rect 28364 56700 28532 56756
rect 28588 58212 28644 58222
rect 27692 56030 27694 56082
rect 27746 56030 27748 56082
rect 27692 56018 27748 56030
rect 27804 56364 28084 56420
rect 27468 55804 27748 55860
rect 27356 55246 27358 55298
rect 27410 55246 27412 55298
rect 27020 54908 27300 54964
rect 27132 54628 27188 54638
rect 27132 54534 27188 54572
rect 26572 54516 26628 54526
rect 26572 53730 26628 54460
rect 26796 54516 26852 54526
rect 26796 54068 26852 54460
rect 26908 54516 26964 54526
rect 26908 54422 26964 54460
rect 27020 54404 27076 54414
rect 27020 54402 27188 54404
rect 27020 54350 27022 54402
rect 27074 54350 27188 54402
rect 27020 54348 27188 54350
rect 27020 54338 27076 54348
rect 26796 54002 26852 54012
rect 27020 53732 27076 53742
rect 26572 53678 26574 53730
rect 26626 53678 26628 53730
rect 26572 53666 26628 53678
rect 26796 53730 27076 53732
rect 26796 53678 27022 53730
rect 27074 53678 27076 53730
rect 26796 53676 27076 53678
rect 26796 53620 26852 53676
rect 27020 53666 27076 53676
rect 27132 53732 27188 54348
rect 27244 54180 27300 54908
rect 27244 54114 27300 54124
rect 27356 53956 27412 55246
rect 27580 55412 27636 55422
rect 27580 55186 27636 55356
rect 27580 55134 27582 55186
rect 27634 55134 27636 55186
rect 27580 55122 27636 55134
rect 27580 54738 27636 54750
rect 27580 54686 27582 54738
rect 27634 54686 27636 54738
rect 27468 54514 27524 54526
rect 27468 54462 27470 54514
rect 27522 54462 27524 54514
rect 27468 54180 27524 54462
rect 27580 54516 27636 54686
rect 27580 54450 27636 54460
rect 27580 54292 27636 54302
rect 27580 54198 27636 54236
rect 27468 54114 27524 54124
rect 27132 53666 27188 53676
rect 27244 53900 27412 53956
rect 26796 53554 26852 53564
rect 26908 52948 26964 52958
rect 26908 52946 27076 52948
rect 26908 52894 26910 52946
rect 26962 52894 27076 52946
rect 26908 52892 27076 52894
rect 26908 52882 26964 52892
rect 26684 52164 26740 52174
rect 26684 52070 26740 52108
rect 26908 51938 26964 51950
rect 26908 51886 26910 51938
rect 26962 51886 26964 51938
rect 26796 51828 26852 51838
rect 26796 51154 26852 51772
rect 26908 51378 26964 51886
rect 26908 51326 26910 51378
rect 26962 51326 26964 51378
rect 26908 51314 26964 51326
rect 27020 51716 27076 52892
rect 26796 51102 26798 51154
rect 26850 51102 26852 51154
rect 26796 51090 26852 51102
rect 26796 50932 26852 50942
rect 26684 50708 26740 50718
rect 26684 50594 26740 50652
rect 26684 50542 26686 50594
rect 26738 50542 26740 50594
rect 26684 50530 26740 50542
rect 26460 50372 26740 50428
rect 26572 49924 26628 49934
rect 26572 49830 26628 49868
rect 26460 49810 26516 49822
rect 26460 49758 26462 49810
rect 26514 49758 26516 49810
rect 26460 49140 26516 49758
rect 26460 49074 26516 49084
rect 26348 48860 26628 48916
rect 25788 48804 25844 48814
rect 25788 48802 26516 48804
rect 25788 48750 25790 48802
rect 25842 48750 26516 48802
rect 25788 48748 26516 48750
rect 25788 48738 25844 48748
rect 25340 48414 25342 48466
rect 25394 48414 25396 48466
rect 25340 48402 25396 48414
rect 26460 48354 26516 48748
rect 26460 48302 26462 48354
rect 26514 48302 26516 48354
rect 26460 48290 26516 48302
rect 25228 48242 25284 48254
rect 25228 48190 25230 48242
rect 25282 48190 25284 48242
rect 25116 47572 25172 47582
rect 24892 46946 24948 46956
rect 25004 47346 25060 47358
rect 25004 47294 25006 47346
rect 25058 47294 25060 47346
rect 25004 46900 25060 47294
rect 25116 47346 25172 47516
rect 25228 47460 25284 48190
rect 25452 48242 25508 48254
rect 25452 48190 25454 48242
rect 25506 48190 25508 48242
rect 25228 47394 25284 47404
rect 25340 47460 25396 47470
rect 25452 47460 25508 48190
rect 25788 48242 25844 48254
rect 25788 48190 25790 48242
rect 25842 48190 25844 48242
rect 25788 48132 25844 48190
rect 26572 48132 26628 48860
rect 25788 48066 25844 48076
rect 26348 48076 26628 48132
rect 25676 47572 25732 47582
rect 25676 47478 25732 47516
rect 26236 47572 26292 47582
rect 25340 47458 25508 47460
rect 25340 47406 25342 47458
rect 25394 47406 25508 47458
rect 25340 47404 25508 47406
rect 25340 47394 25396 47404
rect 25116 47294 25118 47346
rect 25170 47294 25172 47346
rect 25116 47282 25172 47294
rect 26124 47236 26180 47246
rect 26124 47142 26180 47180
rect 25004 46844 25844 46900
rect 25116 46676 25172 46686
rect 25116 46582 25172 46620
rect 25564 46674 25620 46686
rect 25564 46622 25566 46674
rect 25618 46622 25620 46674
rect 25340 46564 25396 46574
rect 25340 46470 25396 46508
rect 25564 46452 25620 46622
rect 25564 46386 25620 46396
rect 25676 46674 25732 46686
rect 25676 46622 25678 46674
rect 25730 46622 25732 46674
rect 24892 46116 24948 46126
rect 24892 46002 24948 46060
rect 24892 45950 24894 46002
rect 24946 45950 24948 46002
rect 24892 45938 24948 45950
rect 25676 45892 25732 46622
rect 25788 46676 25844 46844
rect 26236 46898 26292 47516
rect 26236 46846 26238 46898
rect 26290 46846 26292 46898
rect 26236 46834 26292 46846
rect 26124 46676 26180 46686
rect 25788 46674 26180 46676
rect 25788 46622 26126 46674
rect 26178 46622 26180 46674
rect 25788 46620 26180 46622
rect 25452 45332 25508 45342
rect 24780 45276 25060 45332
rect 24668 44994 24724 45006
rect 24668 44942 24670 44994
rect 24722 44942 24724 44994
rect 24668 44882 24724 44942
rect 24668 44830 24670 44882
rect 24722 44830 24724 44882
rect 24668 44434 24724 44830
rect 24668 44382 24670 44434
rect 24722 44382 24724 44434
rect 24668 44324 24724 44382
rect 24668 44258 24724 44268
rect 24892 44324 24948 44334
rect 24892 44230 24948 44268
rect 24556 42354 24612 42364
rect 24668 43764 24724 43774
rect 24444 41134 24446 41186
rect 24498 41134 24500 41186
rect 24444 39620 24500 41134
rect 24668 41860 24724 43708
rect 25004 42756 25060 45276
rect 25228 45220 25284 45230
rect 25228 45106 25284 45164
rect 25228 45054 25230 45106
rect 25282 45054 25284 45106
rect 25228 45042 25284 45054
rect 25452 44882 25508 45276
rect 25452 44830 25454 44882
rect 25506 44830 25508 44882
rect 25452 44818 25508 44830
rect 25564 44996 25620 45006
rect 25116 44548 25172 44558
rect 25116 44454 25172 44492
rect 25340 44322 25396 44334
rect 25340 44270 25342 44322
rect 25394 44270 25396 44322
rect 25340 43764 25396 44270
rect 25564 44324 25620 44940
rect 25676 44436 25732 45836
rect 25900 45220 25956 45230
rect 25900 45126 25956 45164
rect 25788 45108 25844 45118
rect 25788 45014 25844 45052
rect 26012 45106 26068 46620
rect 26124 46610 26180 46620
rect 26236 46452 26292 46462
rect 26236 46358 26292 46396
rect 26348 46004 26404 48076
rect 26572 47572 26628 47582
rect 26572 47478 26628 47516
rect 26684 46900 26740 50372
rect 26796 50036 26852 50876
rect 27020 50484 27076 51660
rect 27020 50418 27076 50428
rect 27132 52050 27188 52062
rect 27132 51998 27134 52050
rect 27186 51998 27188 52050
rect 27132 51492 27188 51998
rect 27132 50482 27188 51436
rect 27132 50430 27134 50482
rect 27186 50430 27188 50482
rect 27132 50418 27188 50430
rect 27244 50036 27300 53900
rect 27580 53620 27636 53630
rect 27468 53284 27524 53294
rect 27468 52946 27524 53228
rect 27468 52894 27470 52946
rect 27522 52894 27524 52946
rect 27468 52882 27524 52894
rect 26796 49980 27300 50036
rect 27468 50596 27524 50606
rect 26796 49810 26852 49822
rect 26796 49758 26798 49810
rect 26850 49758 26852 49810
rect 26796 48242 26852 49758
rect 26908 49026 26964 49980
rect 27132 49812 27188 49822
rect 27132 49364 27188 49756
rect 27132 49298 27188 49308
rect 27356 49140 27412 49150
rect 26908 48974 26910 49026
rect 26962 48974 26964 49026
rect 26908 48962 26964 48974
rect 27020 49028 27076 49038
rect 27020 48804 27076 48972
rect 27356 48916 27412 49084
rect 26796 48190 26798 48242
rect 26850 48190 26852 48242
rect 26796 48178 26852 48190
rect 26908 48748 27076 48804
rect 27132 48914 27412 48916
rect 27132 48862 27358 48914
rect 27410 48862 27412 48914
rect 27132 48860 27412 48862
rect 26908 48020 26964 48748
rect 26684 46834 26740 46844
rect 26796 47964 26964 48020
rect 26796 46676 26852 47964
rect 27132 47236 27188 48860
rect 27356 48850 27412 48860
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 44996 26068 45054
rect 26012 44930 26068 44940
rect 26124 45948 26404 46004
rect 26572 46674 26852 46676
rect 26572 46622 26798 46674
rect 26850 46622 26852 46674
rect 26572 46620 26852 46622
rect 25676 44380 25844 44436
rect 25564 44268 25732 44324
rect 25676 44210 25732 44268
rect 25676 44158 25678 44210
rect 25730 44158 25732 44210
rect 25676 44146 25732 44158
rect 25564 44098 25620 44110
rect 25564 44046 25566 44098
rect 25618 44046 25620 44098
rect 25564 43764 25620 44046
rect 25564 43708 25732 43764
rect 25340 43698 25396 43708
rect 25116 43652 25172 43662
rect 25116 43540 25172 43596
rect 25228 43540 25284 43550
rect 25116 43538 25284 43540
rect 25116 43486 25230 43538
rect 25282 43486 25284 43538
rect 25116 43484 25284 43486
rect 25228 43474 25284 43484
rect 25564 43540 25620 43550
rect 25564 43446 25620 43484
rect 25340 43428 25396 43438
rect 25340 43334 25396 43372
rect 25676 42868 25732 43708
rect 24892 42700 25060 42756
rect 25564 42812 25732 42868
rect 25788 43538 25844 44380
rect 25788 43486 25790 43538
rect 25842 43486 25844 43538
rect 24892 42532 24948 42700
rect 24892 42466 24948 42476
rect 25004 42532 25060 42542
rect 25004 42530 25284 42532
rect 25004 42478 25006 42530
rect 25058 42478 25284 42530
rect 25004 42476 25284 42478
rect 25004 42466 25060 42476
rect 25116 41972 25172 41982
rect 25116 41878 25172 41916
rect 24556 40964 24612 40974
rect 24556 40870 24612 40908
rect 24444 39554 24500 39564
rect 24556 40740 24612 40750
rect 24556 39396 24612 40684
rect 24668 39844 24724 41804
rect 24780 41412 24836 41422
rect 24780 41186 24836 41356
rect 24780 41134 24782 41186
rect 24834 41134 24836 41186
rect 24780 41122 24836 41134
rect 25228 40628 25284 42476
rect 25452 41970 25508 41982
rect 25452 41918 25454 41970
rect 25506 41918 25508 41970
rect 25340 41860 25396 41870
rect 25340 41766 25396 41804
rect 25452 41412 25508 41918
rect 25452 41346 25508 41356
rect 25228 40572 25508 40628
rect 25340 40404 25396 40414
rect 24780 40290 24836 40302
rect 24780 40238 24782 40290
rect 24834 40238 24836 40290
rect 24780 40178 24836 40238
rect 24780 40126 24782 40178
rect 24834 40126 24836 40178
rect 24780 40114 24836 40126
rect 25116 40180 25172 40190
rect 25172 40124 25284 40180
rect 25116 40114 25172 40124
rect 24668 39788 25172 39844
rect 24332 38882 24388 38892
rect 24444 39340 24612 39396
rect 23996 38322 24052 38332
rect 24220 38722 24276 38734
rect 24220 38670 24222 38722
rect 24274 38670 24276 38722
rect 23884 36820 23940 36830
rect 23772 36596 23828 36606
rect 23772 36482 23828 36540
rect 23772 36430 23774 36482
rect 23826 36430 23828 36482
rect 23772 36418 23828 36430
rect 23492 36316 23716 36372
rect 23436 36278 23492 36316
rect 23548 35700 23604 35710
rect 23548 35606 23604 35644
rect 23884 35700 23940 36764
rect 23996 36708 24052 36718
rect 23996 36260 24052 36652
rect 24220 36484 24276 38670
rect 24444 36708 24500 39340
rect 24780 39172 24836 39182
rect 24668 38948 24724 38958
rect 24668 38834 24724 38892
rect 24668 38782 24670 38834
rect 24722 38782 24724 38834
rect 24668 38770 24724 38782
rect 24556 38724 24612 38734
rect 24780 38668 24836 39116
rect 24556 38612 24836 38668
rect 24444 36652 24612 36708
rect 24220 36428 24500 36484
rect 24220 36260 24276 36270
rect 23996 36258 24276 36260
rect 23996 36206 24222 36258
rect 24274 36206 24276 36258
rect 23996 36204 24276 36206
rect 24220 36194 24276 36204
rect 23884 35634 23940 35644
rect 24220 36036 24276 36046
rect 23436 35586 23492 35598
rect 23436 35534 23438 35586
rect 23490 35534 23492 35586
rect 23436 35140 23492 35534
rect 24220 35588 24276 35980
rect 23436 35084 23604 35140
rect 23436 34914 23492 34926
rect 23436 34862 23438 34914
rect 23490 34862 23492 34914
rect 23324 32900 23380 32910
rect 23212 32844 23324 32900
rect 23324 32834 23380 32844
rect 23100 32510 23102 32562
rect 23154 32510 23156 32562
rect 23100 32498 23156 32510
rect 22876 32450 22932 32462
rect 22876 32398 22878 32450
rect 22930 32398 22932 32450
rect 22540 31714 22596 31724
rect 22652 31778 22708 31790
rect 22652 31726 22654 31778
rect 22706 31726 22708 31778
rect 22540 31556 22596 31566
rect 22540 30996 22596 31500
rect 22652 31220 22708 31726
rect 22876 31444 22932 32398
rect 23324 31892 23380 31902
rect 23324 31798 23380 31836
rect 22876 31378 22932 31388
rect 23324 31220 23380 31230
rect 22652 31218 23380 31220
rect 22652 31166 23326 31218
rect 23378 31166 23380 31218
rect 22652 31164 23380 31166
rect 23324 31154 23380 31164
rect 22540 30100 22596 30940
rect 23212 30884 23268 30894
rect 22652 30100 22708 30110
rect 22540 30098 22708 30100
rect 22540 30046 22654 30098
rect 22706 30046 22708 30098
rect 22540 30044 22708 30046
rect 22652 30034 22708 30044
rect 23212 30098 23268 30828
rect 23212 30046 23214 30098
rect 23266 30046 23268 30098
rect 23212 30034 23268 30046
rect 22764 29986 22820 29998
rect 22764 29934 22766 29986
rect 22818 29934 22820 29986
rect 22428 29484 22596 29540
rect 22092 29426 22148 29438
rect 22092 29374 22094 29426
rect 22146 29374 22148 29426
rect 22092 28868 22148 29374
rect 22092 28812 22484 28868
rect 22092 28532 22148 28542
rect 22092 28438 22148 28476
rect 22428 28530 22484 28812
rect 22428 28478 22430 28530
rect 22482 28478 22484 28530
rect 22428 28466 22484 28478
rect 21868 28028 22148 28084
rect 21868 27860 21924 27870
rect 21756 27858 21924 27860
rect 21756 27806 21870 27858
rect 21922 27806 21924 27858
rect 21756 27804 21924 27806
rect 21868 27794 21924 27804
rect 21980 27860 22036 27870
rect 21644 27074 21700 27132
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 21644 27010 21700 27022
rect 21868 27300 21924 27310
rect 21868 26964 21924 27244
rect 21868 26898 21924 26908
rect 21532 25620 21588 25630
rect 21532 25506 21588 25564
rect 21532 25454 21534 25506
rect 21586 25454 21588 25506
rect 21532 25442 21588 25454
rect 21420 25396 21476 25406
rect 21420 25302 21476 25340
rect 20860 24946 21364 24948
rect 20860 24894 21310 24946
rect 21362 24894 21364 24946
rect 20860 24892 21364 24894
rect 20860 24836 20916 24892
rect 21308 24882 21364 24892
rect 20860 24742 20916 24780
rect 21532 23938 21588 23950
rect 21532 23886 21534 23938
rect 21586 23886 21588 23938
rect 20524 22306 20580 22316
rect 20636 23492 20804 23548
rect 20860 23826 20916 23838
rect 20860 23774 20862 23826
rect 20914 23774 20916 23826
rect 20188 21758 20190 21810
rect 20242 21758 20244 21810
rect 20188 21588 20244 21758
rect 20524 21812 20580 21822
rect 20636 21812 20692 23492
rect 20860 23268 20916 23774
rect 21308 23828 21364 23838
rect 21308 23826 21476 23828
rect 21308 23774 21310 23826
rect 21362 23774 21476 23826
rect 21308 23772 21476 23774
rect 21308 23762 21364 23772
rect 21420 23716 21476 23772
rect 21308 23268 21364 23278
rect 20860 23266 21364 23268
rect 20860 23214 21310 23266
rect 21362 23214 21364 23266
rect 20860 23212 21364 23214
rect 21308 22372 21364 23212
rect 21420 23154 21476 23660
rect 21420 23102 21422 23154
rect 21474 23102 21476 23154
rect 21420 23090 21476 23102
rect 21308 22306 21364 22316
rect 21084 22260 21140 22270
rect 20972 21812 21028 21822
rect 20524 21810 20804 21812
rect 20524 21758 20526 21810
rect 20578 21758 20804 21810
rect 20524 21756 20804 21758
rect 20524 21746 20580 21756
rect 20188 21522 20244 21532
rect 20636 21588 20692 21598
rect 20636 21494 20692 21532
rect 19516 21364 19572 21374
rect 19292 20804 19348 20814
rect 19292 20710 19348 20748
rect 18956 20636 19124 20692
rect 18844 20356 18900 20366
rect 18732 19796 18788 19806
rect 18508 19740 18732 19796
rect 18732 19730 18788 19740
rect 17836 18386 17892 18396
rect 18508 18452 18564 18462
rect 16716 17836 16884 17892
rect 16716 17666 16772 17678
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 16716 17556 16772 17614
rect 16716 17490 16772 17500
rect 16828 17332 16884 17836
rect 18508 17666 18564 18396
rect 18732 18338 18788 18350
rect 18732 18286 18734 18338
rect 18786 18286 18788 18338
rect 18732 17892 18788 18286
rect 18508 17614 18510 17666
rect 18562 17614 18564 17666
rect 18508 17602 18564 17614
rect 18620 17890 18788 17892
rect 18620 17838 18734 17890
rect 18786 17838 18788 17890
rect 18620 17836 18788 17838
rect 16604 17054 16606 17106
rect 16658 17054 16660 17106
rect 16604 17042 16660 17054
rect 16716 17276 16884 17332
rect 17388 17554 17444 17566
rect 17388 17502 17390 17554
rect 17442 17502 17444 17554
rect 15708 16818 15764 16828
rect 15820 16884 15876 16894
rect 16156 16884 16212 16894
rect 15820 16882 16212 16884
rect 15820 16830 15822 16882
rect 15874 16830 16158 16882
rect 16210 16830 16212 16882
rect 15820 16828 16212 16830
rect 15820 16818 15876 16828
rect 16156 16818 16212 16828
rect 16268 16884 16324 16894
rect 16268 16770 16324 16828
rect 16268 16718 16270 16770
rect 16322 16718 16324 16770
rect 16268 16706 16324 16718
rect 15372 15092 15652 15148
rect 15708 15540 15764 15550
rect 15372 14420 15428 15092
rect 15708 14644 15764 15484
rect 16156 15540 16212 15550
rect 16212 15484 16324 15540
rect 16156 15474 16212 15484
rect 16268 15426 16324 15484
rect 16268 15374 16270 15426
rect 16322 15374 16324 15426
rect 16268 15362 16324 15374
rect 16716 15148 16772 17276
rect 15708 14530 15764 14588
rect 16492 15092 16772 15148
rect 17388 15148 17444 17502
rect 18620 17108 18676 17836
rect 18732 17826 18788 17836
rect 18396 17052 18676 17108
rect 18396 15426 18452 17052
rect 18732 16884 18788 16894
rect 18732 16790 18788 16828
rect 18844 16770 18900 20300
rect 18844 16718 18846 16770
rect 18898 16718 18900 16770
rect 18844 16706 18900 16718
rect 18732 16660 18788 16670
rect 18732 16548 18788 16604
rect 18732 16492 18900 16548
rect 18396 15374 18398 15426
rect 18450 15374 18452 15426
rect 18396 15362 18452 15374
rect 17724 15314 17780 15326
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17724 15148 17780 15262
rect 17948 15202 18004 15214
rect 17948 15150 17950 15202
rect 18002 15150 18004 15202
rect 17948 15148 18004 15150
rect 17388 15092 17780 15148
rect 17836 15092 18004 15148
rect 16492 14532 16548 15092
rect 15708 14478 15710 14530
rect 15762 14478 15764 14530
rect 15708 14466 15764 14478
rect 16044 14476 16548 14532
rect 15372 14326 15428 14364
rect 16044 14418 16100 14476
rect 16044 14366 16046 14418
rect 16098 14366 16100 14418
rect 16044 14354 16100 14366
rect 16492 14418 16548 14476
rect 16716 14644 16772 14654
rect 16492 14366 16494 14418
rect 16546 14366 16548 14418
rect 16268 14308 16324 14318
rect 16156 14306 16324 14308
rect 16156 14254 16270 14306
rect 16322 14254 16324 14306
rect 16156 14252 16324 14254
rect 16156 13972 16212 14252
rect 16268 14242 16324 14252
rect 15708 13916 16212 13972
rect 16492 13970 16548 14366
rect 16604 14420 16660 14430
rect 16604 14326 16660 14364
rect 16492 13918 16494 13970
rect 16546 13918 16548 13970
rect 15484 13860 15540 13870
rect 15484 13746 15540 13804
rect 15484 13694 15486 13746
rect 15538 13694 15540 13746
rect 15372 12852 15428 12862
rect 15260 12796 15372 12852
rect 15372 12404 15428 12796
rect 15372 12338 15428 12348
rect 14700 12126 14702 12178
rect 14754 12126 14756 12178
rect 14700 11394 14756 12126
rect 15148 12180 15204 12190
rect 15148 12086 15204 12124
rect 15484 12178 15540 13694
rect 15484 12126 15486 12178
rect 15538 12126 15540 12178
rect 15484 12114 15540 12126
rect 15596 13300 15652 13310
rect 15036 11844 15092 11854
rect 15036 11506 15092 11788
rect 15596 11844 15652 13244
rect 15708 12292 15764 13916
rect 16492 13906 16548 13918
rect 16716 13972 16772 14588
rect 17612 14530 17668 15092
rect 17612 14478 17614 14530
rect 17666 14478 17668 14530
rect 17612 14466 17668 14478
rect 17836 14532 17892 15092
rect 17836 14438 17892 14476
rect 16604 13860 16660 13870
rect 16716 13860 16772 13916
rect 16604 13858 16772 13860
rect 16604 13806 16606 13858
rect 16658 13806 16772 13858
rect 16604 13804 16772 13806
rect 17052 14420 17108 14430
rect 16604 13794 16660 13804
rect 15820 13746 15876 13758
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15820 13412 15876 13694
rect 16044 13748 16100 13758
rect 16268 13748 16324 13758
rect 16044 13746 16324 13748
rect 16044 13694 16046 13746
rect 16098 13694 16270 13746
rect 16322 13694 16324 13746
rect 16044 13692 16324 13694
rect 15932 13636 15988 13646
rect 15932 13542 15988 13580
rect 15820 12404 15876 13356
rect 15932 13300 15988 13310
rect 16044 13300 16100 13692
rect 16268 13682 16324 13692
rect 15988 13244 16100 13300
rect 15932 13234 15988 13244
rect 16044 13132 16436 13188
rect 15932 13076 15988 13086
rect 15932 12982 15988 13020
rect 15932 12404 15988 12414
rect 15820 12402 15988 12404
rect 15820 12350 15934 12402
rect 15986 12350 15988 12402
rect 15820 12348 15988 12350
rect 15932 12338 15988 12348
rect 16044 12402 16100 13132
rect 16380 12964 16436 13132
rect 17052 13074 17108 14364
rect 17388 14308 17444 14318
rect 17388 14214 17444 14252
rect 17724 14306 17780 14318
rect 17724 14254 17726 14306
rect 17778 14254 17780 14306
rect 17052 13022 17054 13074
rect 17106 13022 17108 13074
rect 17052 13010 17108 13022
rect 17612 13524 17668 13534
rect 16604 12964 16660 12974
rect 16380 12962 16660 12964
rect 16380 12910 16606 12962
rect 16658 12910 16660 12962
rect 16380 12908 16660 12910
rect 16604 12898 16660 12908
rect 16044 12350 16046 12402
rect 16098 12350 16100 12402
rect 16044 12338 16100 12350
rect 16156 12850 16212 12862
rect 16156 12798 16158 12850
rect 16210 12798 16212 12850
rect 16156 12404 16212 12798
rect 16604 12404 16660 12414
rect 16156 12348 16324 12404
rect 15708 12236 15876 12292
rect 15820 12180 15876 12236
rect 16156 12180 16212 12190
rect 15876 12178 16212 12180
rect 15876 12126 16158 12178
rect 16210 12126 16212 12178
rect 15876 12124 16212 12126
rect 15820 12086 15876 12124
rect 16156 12114 16212 12124
rect 16268 11844 16324 12348
rect 16604 12310 16660 12348
rect 15596 11778 15652 11788
rect 16156 11788 16324 11844
rect 15036 11454 15038 11506
rect 15090 11454 15092 11506
rect 15036 11442 15092 11454
rect 15148 11618 15204 11630
rect 15148 11566 15150 11618
rect 15202 11566 15204 11618
rect 14700 11342 14702 11394
rect 14754 11342 14756 11394
rect 14700 11330 14756 11342
rect 14588 9662 14590 9714
rect 14642 9662 14644 9714
rect 14364 9604 14420 9614
rect 14364 9154 14420 9548
rect 14364 9102 14366 9154
rect 14418 9102 14420 9154
rect 14364 9090 14420 9102
rect 14252 8990 14254 9042
rect 14306 8990 14308 9042
rect 14252 8978 14308 8990
rect 14588 8428 14644 9662
rect 14924 9156 14980 9166
rect 14924 8428 14980 9100
rect 15036 9044 15092 9054
rect 15148 9044 15204 11566
rect 15708 10052 15764 10062
rect 15596 9828 15652 9838
rect 15036 9042 15204 9044
rect 15036 8990 15038 9042
rect 15090 8990 15204 9042
rect 15036 8988 15204 8990
rect 15036 8978 15092 8988
rect 13468 6690 13636 6692
rect 13468 6638 13470 6690
rect 13522 6638 13636 6690
rect 13468 6636 13636 6638
rect 13692 8372 14644 8428
rect 14812 8372 14980 8428
rect 13692 6914 13748 8372
rect 14812 8258 14868 8372
rect 15148 8370 15204 8988
rect 15148 8318 15150 8370
rect 15202 8318 15204 8370
rect 15148 8306 15204 8318
rect 15484 9602 15540 9614
rect 15484 9550 15486 9602
rect 15538 9550 15540 9602
rect 15484 8372 15540 9550
rect 15596 9042 15652 9772
rect 15708 9154 15764 9996
rect 15820 9940 15876 9950
rect 15820 9714 15876 9884
rect 15820 9662 15822 9714
rect 15874 9662 15876 9714
rect 15820 9650 15876 9662
rect 15708 9102 15710 9154
rect 15762 9102 15764 9154
rect 15708 9090 15764 9102
rect 15596 8990 15598 9042
rect 15650 8990 15652 9042
rect 15596 8978 15652 8990
rect 15484 8306 15540 8316
rect 15932 8930 15988 8942
rect 15932 8878 15934 8930
rect 15986 8878 15988 8930
rect 14812 8206 14814 8258
rect 14866 8206 14868 8258
rect 14812 7364 14868 8206
rect 15708 8260 15764 8270
rect 15708 8166 15764 8204
rect 13692 6862 13694 6914
rect 13746 6862 13748 6914
rect 13692 6692 13748 6862
rect 14700 7308 14868 7364
rect 13692 6636 14308 6692
rect 13468 6626 13524 6636
rect 13356 6412 13524 6468
rect 13468 5908 13524 6412
rect 13580 6018 13636 6636
rect 13580 5966 13582 6018
rect 13634 5966 13636 6018
rect 13580 5954 13636 5966
rect 14028 6466 14084 6478
rect 14028 6414 14030 6466
rect 14082 6414 14084 6466
rect 13468 5814 13524 5852
rect 14028 5124 14084 6414
rect 14252 5906 14308 6636
rect 14252 5854 14254 5906
rect 14306 5854 14308 5906
rect 14252 5842 14308 5854
rect 14364 5908 14420 5918
rect 14420 5852 14532 5908
rect 14364 5842 14420 5852
rect 14476 5236 14532 5852
rect 14588 5684 14644 5694
rect 14588 5590 14644 5628
rect 14588 5236 14644 5246
rect 14476 5234 14644 5236
rect 14476 5182 14590 5234
rect 14642 5182 14644 5234
rect 14476 5180 14644 5182
rect 14588 5170 14644 5180
rect 14364 5124 14420 5134
rect 14028 5122 14532 5124
rect 14028 5070 14366 5122
rect 14418 5070 14532 5122
rect 14028 5068 14532 5070
rect 14364 5058 14420 5068
rect 14476 5012 14532 5068
rect 14700 5012 14756 7308
rect 15932 6692 15988 8878
rect 15596 6690 15988 6692
rect 15596 6638 15934 6690
rect 15986 6638 15988 6690
rect 15596 6636 15988 6638
rect 15596 5906 15652 6636
rect 15932 6626 15988 6636
rect 15596 5854 15598 5906
rect 15650 5854 15652 5906
rect 15596 5842 15652 5854
rect 15708 6466 15764 6478
rect 15708 6414 15710 6466
rect 15762 6414 15764 6466
rect 15036 5796 15092 5806
rect 15036 5234 15092 5740
rect 15708 5796 15764 6414
rect 15820 6466 15876 6478
rect 15820 6414 15822 6466
rect 15874 6414 15876 6466
rect 15820 6020 15876 6414
rect 15820 5964 15988 6020
rect 15820 5796 15876 5806
rect 15764 5794 15876 5796
rect 15764 5742 15822 5794
rect 15874 5742 15876 5794
rect 15764 5740 15876 5742
rect 15708 5702 15764 5740
rect 15820 5730 15876 5740
rect 15036 5182 15038 5234
rect 15090 5182 15092 5234
rect 15036 5170 15092 5182
rect 15932 5234 15988 5964
rect 15932 5182 15934 5234
rect 15986 5182 15988 5234
rect 15932 5170 15988 5182
rect 14476 4956 14756 5012
rect 16156 5010 16212 11788
rect 16604 10052 16660 10062
rect 16268 9940 16324 9950
rect 16268 9846 16324 9884
rect 16604 9826 16660 9996
rect 17164 9940 17220 9950
rect 17164 9846 17220 9884
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16604 9762 16660 9774
rect 16492 8372 16548 8382
rect 16492 8258 16548 8316
rect 16492 8206 16494 8258
rect 16546 8206 16548 8258
rect 16492 8194 16548 8206
rect 16604 8370 16660 8382
rect 16604 8318 16606 8370
rect 16658 8318 16660 8370
rect 16604 8260 16660 8318
rect 16604 8194 16660 8204
rect 17388 8148 17444 8158
rect 17388 8054 17444 8092
rect 16380 6692 16436 6702
rect 16380 6690 16548 6692
rect 16380 6638 16382 6690
rect 16434 6638 16548 6690
rect 16380 6636 16548 6638
rect 16380 6626 16436 6636
rect 16492 6130 16548 6636
rect 16492 6078 16494 6130
rect 16546 6078 16548 6130
rect 16492 6066 16548 6078
rect 16716 6018 16772 6030
rect 16716 5966 16718 6018
rect 16770 5966 16772 6018
rect 16268 5908 16324 5918
rect 16268 5814 16324 5852
rect 16716 5908 16772 5966
rect 16828 6020 16884 6030
rect 17612 6020 17668 13468
rect 17724 11620 17780 14254
rect 18732 13972 18788 13982
rect 18732 13878 18788 13916
rect 18844 13858 18900 16492
rect 18844 13806 18846 13858
rect 18898 13806 18900 13858
rect 18844 13794 18900 13806
rect 18732 13522 18788 13534
rect 18732 13470 18734 13522
rect 18786 13470 18788 13522
rect 18620 12740 18676 12750
rect 18508 12684 18620 12740
rect 18172 12178 18228 12190
rect 18172 12126 18174 12178
rect 18226 12126 18228 12178
rect 17724 11564 18004 11620
rect 17948 10612 18004 11564
rect 18172 11172 18228 12126
rect 18172 11106 18228 11116
rect 17948 10610 18228 10612
rect 17948 10558 17950 10610
rect 18002 10558 18228 10610
rect 17948 10556 18228 10558
rect 17948 10546 18004 10556
rect 17724 10498 17780 10510
rect 17724 10446 17726 10498
rect 17778 10446 17780 10498
rect 17724 9604 17780 10446
rect 18172 9938 18228 10556
rect 18172 9886 18174 9938
rect 18226 9886 18228 9938
rect 18172 9874 18228 9886
rect 17724 9538 17780 9548
rect 18396 9826 18452 9838
rect 18396 9774 18398 9826
rect 18450 9774 18452 9826
rect 18396 9604 18452 9774
rect 18396 9538 18452 9548
rect 18508 9380 18564 12684
rect 18620 12674 18676 12684
rect 18732 12066 18788 13470
rect 18956 13412 19012 20636
rect 19180 18340 19236 18350
rect 19180 18246 19236 18284
rect 19068 17556 19124 17566
rect 19068 17462 19124 17500
rect 19180 16770 19236 16782
rect 19180 16718 19182 16770
rect 19234 16718 19236 16770
rect 19180 16100 19236 16718
rect 19180 16034 19236 16044
rect 19292 15988 19348 15998
rect 19292 15894 19348 15932
rect 19516 13634 19572 21308
rect 20524 21364 20580 21374
rect 20524 21270 20580 21308
rect 20300 21252 20356 21262
rect 19628 20914 19684 20926
rect 19628 20862 19630 20914
rect 19682 20862 19684 20914
rect 19628 20020 19684 20862
rect 20300 20802 20356 21196
rect 20300 20750 20302 20802
rect 20354 20750 20356 20802
rect 20300 20738 20356 20750
rect 19964 20690 20020 20702
rect 19964 20638 19966 20690
rect 20018 20638 20020 20690
rect 19964 20580 20020 20638
rect 20188 20692 20244 20702
rect 20076 20580 20132 20590
rect 19964 20524 20076 20580
rect 20076 20514 20132 20524
rect 20188 20578 20244 20636
rect 20748 20692 20804 21756
rect 20748 20626 20804 20636
rect 20188 20526 20190 20578
rect 20242 20526 20244 20578
rect 20188 20514 20244 20526
rect 20412 20580 20468 20590
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19740 20020 19796 20030
rect 19628 19964 19740 20020
rect 19740 19926 19796 19964
rect 20412 20018 20468 20524
rect 20412 19966 20414 20018
rect 20466 19966 20468 20018
rect 20412 19954 20468 19966
rect 19628 19796 19684 19806
rect 19628 15092 19684 19740
rect 20300 19794 20356 19806
rect 20300 19742 20302 19794
rect 20354 19742 20356 19794
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20300 18450 20356 19742
rect 20972 18562 21028 21756
rect 20972 18510 20974 18562
rect 21026 18510 21028 18562
rect 20972 18498 21028 18510
rect 20300 18398 20302 18450
rect 20354 18398 20356 18450
rect 20076 18340 20132 18350
rect 20076 18246 20132 18284
rect 20300 17666 20356 18398
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 17602 20356 17614
rect 20524 18340 20580 18350
rect 21084 18340 21140 22204
rect 21532 22148 21588 23886
rect 21868 23716 21924 23726
rect 21756 23714 21924 23716
rect 21756 23662 21870 23714
rect 21922 23662 21924 23714
rect 21756 23660 21924 23662
rect 21756 22370 21812 23660
rect 21868 23650 21924 23660
rect 21756 22318 21758 22370
rect 21810 22318 21812 22370
rect 21756 22306 21812 22318
rect 21532 22082 21588 22092
rect 21420 20804 21476 20814
rect 21196 20692 21252 20702
rect 21196 20242 21252 20636
rect 21196 20190 21198 20242
rect 21250 20190 21252 20242
rect 21196 20178 21252 20190
rect 21420 19124 21476 20748
rect 21532 20132 21588 20142
rect 21532 20038 21588 20076
rect 21868 20020 21924 20030
rect 21868 19926 21924 19964
rect 21980 19796 22036 27804
rect 22092 26516 22148 28028
rect 22540 26908 22596 29484
rect 22652 28644 22708 28654
rect 22652 28550 22708 28588
rect 22764 27972 22820 29934
rect 22820 27916 23044 27972
rect 22764 27906 22820 27916
rect 22764 27188 22820 27198
rect 22820 27132 22932 27188
rect 22764 27094 22820 27132
rect 22764 26964 22820 26974
rect 22092 26422 22148 26460
rect 22204 26850 22260 26862
rect 22540 26852 22708 26908
rect 22204 26798 22206 26850
rect 22258 26798 22260 26850
rect 22204 26292 22260 26798
rect 22428 26292 22484 26302
rect 22204 26290 22484 26292
rect 22204 26238 22430 26290
rect 22482 26238 22484 26290
rect 22204 26236 22484 26238
rect 22428 26226 22484 26236
rect 22316 23154 22372 23166
rect 22316 23102 22318 23154
rect 22370 23102 22372 23154
rect 22092 22484 22148 22494
rect 22092 22390 22148 22428
rect 22204 22372 22260 22382
rect 22204 22278 22260 22316
rect 22204 22148 22260 22158
rect 22316 22148 22372 23102
rect 22260 22092 22372 22148
rect 22204 22082 22260 22092
rect 22652 21252 22708 26852
rect 22764 24724 22820 26908
rect 22876 25172 22932 27132
rect 22988 26962 23044 27916
rect 22988 26910 22990 26962
rect 23042 26910 23044 26962
rect 22988 26740 23044 26910
rect 23100 27970 23156 27982
rect 23100 27918 23102 27970
rect 23154 27918 23156 27970
rect 23100 27636 23156 27918
rect 23436 27972 23492 34862
rect 23548 34244 23604 35084
rect 24220 34914 24276 35532
rect 24220 34862 24222 34914
rect 24274 34862 24276 34914
rect 24220 34850 24276 34862
rect 23660 34244 23716 34254
rect 23548 34242 23716 34244
rect 23548 34190 23662 34242
rect 23714 34190 23716 34242
rect 23548 34188 23716 34190
rect 23660 34132 23716 34188
rect 23660 34076 23940 34132
rect 23548 31780 23604 31790
rect 23548 31686 23604 31724
rect 23884 31666 23940 34076
rect 23884 31614 23886 31666
rect 23938 31614 23940 31666
rect 23772 31556 23828 31566
rect 23772 31462 23828 31500
rect 23548 30994 23604 31006
rect 23548 30942 23550 30994
rect 23602 30942 23604 30994
rect 23548 30212 23604 30942
rect 23884 30884 23940 31614
rect 23884 30818 23940 30828
rect 23996 32340 24052 32350
rect 23548 30118 23604 30156
rect 23996 30212 24052 32284
rect 23996 30146 24052 30156
rect 24220 28756 24276 28766
rect 24220 28662 24276 28700
rect 23436 27906 23492 27916
rect 23100 26964 23156 27580
rect 23100 26898 23156 26908
rect 23436 27746 23492 27758
rect 23436 27694 23438 27746
rect 23490 27694 23492 27746
rect 23436 26908 23492 27694
rect 23772 27746 23828 27758
rect 23772 27694 23774 27746
rect 23826 27694 23828 27746
rect 23772 27188 23828 27694
rect 23996 27636 24052 27646
rect 23996 27542 24052 27580
rect 24332 27634 24388 27646
rect 24332 27582 24334 27634
rect 24386 27582 24388 27634
rect 23772 27122 23828 27132
rect 24220 27076 24276 27114
rect 24220 27010 24276 27020
rect 24332 26908 24388 27582
rect 23436 26852 24052 26908
rect 22988 26684 23380 26740
rect 23100 26290 23156 26302
rect 23100 26238 23102 26290
rect 23154 26238 23156 26290
rect 23100 25394 23156 26238
rect 23324 25506 23380 26684
rect 23324 25454 23326 25506
rect 23378 25454 23380 25506
rect 23324 25442 23380 25454
rect 23436 26290 23492 26302
rect 23436 26238 23438 26290
rect 23490 26238 23492 26290
rect 23100 25342 23102 25394
rect 23154 25342 23156 25394
rect 23100 25330 23156 25342
rect 22876 25116 23268 25172
rect 22988 24724 23044 24734
rect 22764 24722 23044 24724
rect 22764 24670 22990 24722
rect 23042 24670 23044 24722
rect 22764 24668 23044 24670
rect 22988 24658 23044 24668
rect 23212 24722 23268 25116
rect 23436 24948 23492 26238
rect 23772 26292 23828 26302
rect 23772 26198 23828 26236
rect 23996 26290 24052 26852
rect 23996 26238 23998 26290
rect 24050 26238 24052 26290
rect 23996 26226 24052 26238
rect 24220 26852 24388 26908
rect 24444 26908 24500 36428
rect 24556 36036 24612 36652
rect 24556 35970 24612 35980
rect 24556 35252 24612 35262
rect 24556 34354 24612 35196
rect 24556 34302 24558 34354
rect 24610 34302 24612 34354
rect 24556 34290 24612 34302
rect 24556 33348 24612 33358
rect 24780 33348 24836 38612
rect 24892 38388 24948 38398
rect 24892 38274 24948 38332
rect 24892 38222 24894 38274
rect 24946 38222 24948 38274
rect 24892 38210 24948 38222
rect 25004 38052 25060 38062
rect 25004 37958 25060 37996
rect 24892 37828 24948 37838
rect 24892 34914 24948 37772
rect 24892 34862 24894 34914
rect 24946 34862 24948 34914
rect 24892 34356 24948 34862
rect 24892 34290 24948 34300
rect 25004 36258 25060 36270
rect 25004 36206 25006 36258
rect 25058 36206 25060 36258
rect 24556 33346 24836 33348
rect 24556 33294 24558 33346
rect 24610 33294 24836 33346
rect 24556 33292 24836 33294
rect 24556 33282 24612 33292
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 24780 31332 24836 31342
rect 24668 29652 24724 29662
rect 24668 29558 24724 29596
rect 24444 26852 24612 26908
rect 24108 26066 24164 26078
rect 24108 26014 24110 26066
rect 24162 26014 24164 26066
rect 23548 24948 23604 24958
rect 23436 24946 23716 24948
rect 23436 24894 23550 24946
rect 23602 24894 23716 24946
rect 23436 24892 23716 24894
rect 23548 24882 23604 24892
rect 23212 24670 23214 24722
rect 23266 24670 23268 24722
rect 23212 24658 23268 24670
rect 23436 24612 23492 24622
rect 23212 23940 23268 23950
rect 23212 23846 23268 23884
rect 22876 23828 22932 23838
rect 22876 23266 22932 23772
rect 22988 23714 23044 23726
rect 22988 23662 22990 23714
rect 23042 23662 23044 23714
rect 22988 23604 23044 23662
rect 22988 23538 23044 23548
rect 22876 23214 22878 23266
rect 22930 23214 22932 23266
rect 22876 23202 22932 23214
rect 22876 22260 22932 22270
rect 22876 22258 23380 22260
rect 22876 22206 22878 22258
rect 22930 22206 23380 22258
rect 22876 22204 23380 22206
rect 22876 22194 22932 22204
rect 22204 21196 22708 21252
rect 22092 20244 22148 20254
rect 22092 20150 22148 20188
rect 21980 19740 22148 19796
rect 21980 19572 22036 19582
rect 21532 19348 21588 19358
rect 21980 19348 22036 19516
rect 21532 19346 22036 19348
rect 21532 19294 21534 19346
rect 21586 19294 22036 19346
rect 21532 19292 22036 19294
rect 21532 19282 21588 19292
rect 21980 19234 22036 19292
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21980 19170 22036 19182
rect 21756 19124 21812 19134
rect 21420 19122 21812 19124
rect 21420 19070 21758 19122
rect 21810 19070 21812 19122
rect 21420 19068 21812 19070
rect 21756 19058 21812 19068
rect 21868 19012 21924 19022
rect 21756 18450 21812 18462
rect 21756 18398 21758 18450
rect 21810 18398 21812 18450
rect 20524 17666 20580 18284
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 20972 18284 21140 18340
rect 21420 18340 21476 18350
rect 21756 18340 21812 18398
rect 21420 18338 21812 18340
rect 21420 18286 21422 18338
rect 21474 18286 21812 18338
rect 21420 18284 21812 18286
rect 19964 17556 20020 17566
rect 19964 17462 20020 17500
rect 20412 17442 20468 17454
rect 20412 17390 20414 17442
rect 20466 17390 20468 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 16212 20244 16222
rect 20188 16118 20244 16156
rect 19964 16100 20020 16110
rect 19964 16006 20020 16044
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20412 15148 20468 17390
rect 20860 16212 20916 16222
rect 20860 16118 20916 16156
rect 20412 15092 20692 15148
rect 19628 13972 19684 15036
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20636 13972 20692 15092
rect 20972 14532 21028 18284
rect 21420 18116 21476 18284
rect 21868 18228 21924 18956
rect 21420 18050 21476 18060
rect 21644 18172 21924 18228
rect 21644 17108 21700 18172
rect 21532 17106 21700 17108
rect 21532 17054 21646 17106
rect 21698 17054 21700 17106
rect 21532 17052 21700 17054
rect 21420 16996 21476 17006
rect 21420 16902 21476 16940
rect 21084 16884 21140 16894
rect 21084 16790 21140 16828
rect 21308 16658 21364 16670
rect 21308 16606 21310 16658
rect 21362 16606 21364 16658
rect 21308 16098 21364 16606
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 16034 21364 16046
rect 21532 15540 21588 17052
rect 21644 17042 21700 17052
rect 22092 16212 22148 19740
rect 22204 19572 22260 21196
rect 22540 20578 22596 20590
rect 22540 20526 22542 20578
rect 22594 20526 22596 20578
rect 22540 20244 22596 20526
rect 22540 20178 22596 20188
rect 22316 20132 22372 20142
rect 22316 20020 22372 20076
rect 23212 20132 23268 20142
rect 22764 20020 22820 20030
rect 22316 20018 23044 20020
rect 22316 19966 22766 20018
rect 22818 19966 23044 20018
rect 22316 19964 23044 19966
rect 22764 19954 22820 19964
rect 22428 19796 22484 19806
rect 22428 19794 22820 19796
rect 22428 19742 22430 19794
rect 22482 19742 22820 19794
rect 22428 19740 22820 19742
rect 22428 19730 22484 19740
rect 22204 19516 22708 19572
rect 22316 19236 22372 19246
rect 22540 19236 22596 19246
rect 22316 19234 22596 19236
rect 22316 19182 22318 19234
rect 22370 19182 22542 19234
rect 22594 19182 22596 19234
rect 22316 19180 22596 19182
rect 22316 19170 22372 19180
rect 22540 19170 22596 19180
rect 22204 19012 22260 19022
rect 22204 18918 22260 18956
rect 22540 18452 22596 18462
rect 22652 18452 22708 19516
rect 22764 19458 22820 19740
rect 22764 19406 22766 19458
rect 22818 19406 22820 19458
rect 22764 19394 22820 19406
rect 22540 18450 22708 18452
rect 22540 18398 22542 18450
rect 22594 18398 22708 18450
rect 22540 18396 22708 18398
rect 22540 18386 22596 18396
rect 22652 18340 22708 18396
rect 22652 18274 22708 18284
rect 22204 16996 22260 17006
rect 22204 16902 22260 16940
rect 22092 16118 22148 16156
rect 21980 16100 22036 16110
rect 21980 16006 22036 16044
rect 22652 15986 22708 15998
rect 22652 15934 22654 15986
rect 22706 15934 22708 15986
rect 21532 15446 21588 15484
rect 22316 15876 22372 15886
rect 22316 15540 22372 15820
rect 21196 15314 21252 15326
rect 21196 15262 21198 15314
rect 21250 15262 21252 15314
rect 21196 15092 21252 15262
rect 21252 15036 21476 15092
rect 21196 15026 21252 15036
rect 20972 14476 21364 14532
rect 21196 14306 21252 14318
rect 21196 14254 21198 14306
rect 21250 14254 21252 14306
rect 20636 13916 20916 13972
rect 19628 13906 19684 13916
rect 20076 13748 20132 13758
rect 20636 13748 20692 13758
rect 20076 13746 20636 13748
rect 20076 13694 20078 13746
rect 20130 13694 20636 13746
rect 20076 13692 20636 13694
rect 20076 13682 20132 13692
rect 20636 13654 20692 13692
rect 19516 13582 19518 13634
rect 19570 13582 19572 13634
rect 19516 13570 19572 13582
rect 19292 13524 19348 13534
rect 19292 13430 19348 13468
rect 18732 12014 18734 12066
rect 18786 12014 18788 12066
rect 18732 11394 18788 12014
rect 18732 11342 18734 11394
rect 18786 11342 18788 11394
rect 18732 11330 18788 11342
rect 18844 13356 19012 13412
rect 18844 11396 18900 13356
rect 18956 13186 19012 13198
rect 18956 13134 18958 13186
rect 19010 13134 19012 13186
rect 18956 13076 19012 13134
rect 19628 13076 19684 13086
rect 18956 13020 19236 13076
rect 19180 12964 19236 13020
rect 19404 12964 19460 12974
rect 19180 12962 19460 12964
rect 19180 12910 19406 12962
rect 19458 12910 19460 12962
rect 19180 12908 19460 12910
rect 19404 12898 19460 12908
rect 19068 12852 19124 12862
rect 19068 12758 19124 12796
rect 19628 12852 19684 13020
rect 20076 13076 20132 13086
rect 20076 12982 20132 13020
rect 20412 13076 20468 13086
rect 18956 12738 19012 12750
rect 18956 12686 18958 12738
rect 19010 12686 19012 12738
rect 18956 12292 19012 12686
rect 19516 12738 19572 12750
rect 19516 12686 19518 12738
rect 19570 12686 19572 12738
rect 19068 12292 19124 12302
rect 19404 12292 19460 12302
rect 18956 12290 19460 12292
rect 18956 12238 19070 12290
rect 19122 12238 19406 12290
rect 19458 12238 19460 12290
rect 18956 12236 19460 12238
rect 19068 12226 19124 12236
rect 19404 12226 19460 12236
rect 19068 11844 19124 11854
rect 19068 11732 19124 11788
rect 19068 11676 19236 11732
rect 18844 11340 19124 11396
rect 18844 11172 18900 11182
rect 18732 11170 18900 11172
rect 18732 11118 18846 11170
rect 18898 11118 18900 11170
rect 18732 11116 18900 11118
rect 18620 10612 18676 10622
rect 18620 10518 18676 10556
rect 18732 9940 18788 11116
rect 18844 11106 18900 11116
rect 18956 11172 19012 11182
rect 18956 11078 19012 11116
rect 18620 9884 18788 9940
rect 18620 9492 18676 9884
rect 18732 9716 18788 9726
rect 18732 9622 18788 9660
rect 18620 9436 19012 9492
rect 18508 9324 18788 9380
rect 17948 8372 18004 8382
rect 17724 8260 17780 8270
rect 17724 8166 17780 8204
rect 17948 8146 18004 8316
rect 18060 8372 18116 8382
rect 18060 8370 18340 8372
rect 18060 8318 18062 8370
rect 18114 8318 18340 8370
rect 18060 8316 18340 8318
rect 18060 8306 18116 8316
rect 17948 8094 17950 8146
rect 18002 8094 18004 8146
rect 17948 8082 18004 8094
rect 18172 6690 18228 6702
rect 18172 6638 18174 6690
rect 18226 6638 18228 6690
rect 18172 6132 18228 6638
rect 18284 6580 18340 8316
rect 18732 8370 18788 9324
rect 18732 8318 18734 8370
rect 18786 8318 18788 8370
rect 18620 8258 18676 8270
rect 18620 8206 18622 8258
rect 18674 8206 18676 8258
rect 18620 8148 18676 8206
rect 18396 8092 18620 8148
rect 18396 7698 18452 8092
rect 18620 8082 18676 8092
rect 18396 7646 18398 7698
rect 18450 7646 18452 7698
rect 18396 7634 18452 7646
rect 18620 7588 18676 7598
rect 18732 7588 18788 8318
rect 18620 7586 18788 7588
rect 18620 7534 18622 7586
rect 18674 7534 18788 7586
rect 18620 7532 18788 7534
rect 18620 7522 18676 7532
rect 18396 7362 18452 7374
rect 18396 7310 18398 7362
rect 18450 7310 18452 7362
rect 18396 6692 18452 7310
rect 18732 6692 18788 6702
rect 18396 6690 18788 6692
rect 18396 6638 18734 6690
rect 18786 6638 18788 6690
rect 18396 6636 18788 6638
rect 18956 6692 19012 9436
rect 19068 6804 19124 11340
rect 19180 10498 19236 11676
rect 19404 11396 19460 11406
rect 19516 11396 19572 12686
rect 19628 12178 19684 12796
rect 19740 12740 19796 12778
rect 19740 12674 19796 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20412 12402 20468 13020
rect 20412 12350 20414 12402
rect 20466 12350 20468 12402
rect 20412 12338 20468 12350
rect 19628 12126 19630 12178
rect 19682 12126 19684 12178
rect 19628 12114 19684 12126
rect 19964 11954 20020 11966
rect 19964 11902 19966 11954
rect 20018 11902 20020 11954
rect 19964 11396 20020 11902
rect 19404 11394 20020 11396
rect 19404 11342 19406 11394
rect 19458 11342 20020 11394
rect 19404 11340 20020 11342
rect 19404 11330 19460 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19628 10612 19684 10622
rect 20076 10612 20132 10622
rect 19684 10556 19796 10612
rect 19628 10518 19684 10556
rect 19180 10446 19182 10498
rect 19234 10446 19236 10498
rect 19180 9828 19236 10446
rect 19740 9828 19796 10556
rect 20076 10518 20132 10556
rect 20748 10612 20804 10622
rect 20748 10498 20804 10556
rect 20748 10446 20750 10498
rect 20802 10446 20804 10498
rect 20748 10434 20804 10446
rect 20860 10610 20916 13916
rect 21084 13746 21140 13758
rect 21084 13694 21086 13746
rect 21138 13694 21140 13746
rect 21084 13636 21140 13694
rect 21084 13570 21140 13580
rect 21196 13634 21252 14254
rect 21196 13582 21198 13634
rect 21250 13582 21252 13634
rect 21196 13570 21252 13582
rect 20860 10558 20862 10610
rect 20914 10558 20916 10610
rect 19852 9828 19908 9838
rect 19740 9826 19908 9828
rect 19740 9774 19854 9826
rect 19906 9774 19908 9826
rect 19740 9772 19908 9774
rect 19180 9762 19236 9772
rect 19852 9762 19908 9772
rect 20188 9828 20244 9838
rect 20188 9734 20244 9772
rect 19628 9716 19684 9726
rect 19628 9622 19684 9660
rect 20860 9716 20916 10558
rect 21308 10388 21364 14476
rect 21420 14418 21476 15036
rect 21532 14532 21588 14542
rect 21532 14438 21588 14476
rect 21756 14530 21812 14542
rect 21756 14478 21758 14530
rect 21810 14478 21812 14530
rect 21420 14366 21422 14418
rect 21474 14366 21476 14418
rect 21420 14354 21476 14366
rect 21756 13636 21812 14478
rect 22316 14418 22372 15484
rect 22540 15428 22596 15438
rect 22540 15148 22596 15372
rect 22428 15092 22596 15148
rect 22428 14754 22484 15092
rect 22428 14702 22430 14754
rect 22482 14702 22484 14754
rect 22428 14690 22484 14702
rect 22652 14644 22708 15934
rect 22876 15428 22932 15438
rect 22876 15334 22932 15372
rect 22316 14366 22318 14418
rect 22370 14366 22372 14418
rect 22316 14354 22372 14366
rect 22540 14588 22708 14644
rect 22764 15314 22820 15326
rect 22764 15262 22766 15314
rect 22818 15262 22820 15314
rect 22092 14308 22148 14318
rect 22092 14214 22148 14252
rect 22540 13972 22596 14588
rect 22652 14420 22708 14430
rect 22652 14326 22708 14364
rect 22764 14308 22820 15262
rect 22876 15090 22932 15102
rect 22876 15038 22878 15090
rect 22930 15038 22932 15090
rect 22876 14530 22932 15038
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22876 14466 22932 14478
rect 22764 14252 22932 14308
rect 22428 13916 22596 13972
rect 22876 13970 22932 14252
rect 22876 13918 22878 13970
rect 22930 13918 22932 13970
rect 22204 13748 22260 13758
rect 22204 13654 22260 13692
rect 21756 13570 21812 13580
rect 21532 10724 21588 10734
rect 21532 10630 21588 10668
rect 21868 10612 21924 10622
rect 21308 10332 21476 10388
rect 20860 9650 20916 9660
rect 20076 9604 20132 9614
rect 20076 9602 20244 9604
rect 20076 9550 20078 9602
rect 20130 9550 20244 9602
rect 20076 9548 20244 9550
rect 20076 9538 20132 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9548
rect 20076 9212 20244 9268
rect 19516 8148 19572 8158
rect 19516 8054 19572 8092
rect 20076 8036 20132 9212
rect 20748 8372 20804 8382
rect 20748 8370 21364 8372
rect 20748 8318 20750 8370
rect 20802 8318 21364 8370
rect 20748 8316 21364 8318
rect 20748 8306 20804 8316
rect 20412 8148 20468 8158
rect 20468 8092 20580 8148
rect 20412 8054 20468 8092
rect 20132 7980 20356 8036
rect 20076 7970 20132 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20300 7474 20356 7980
rect 20300 7422 20302 7474
rect 20354 7422 20356 7474
rect 20300 7410 20356 7422
rect 20524 7362 20580 8092
rect 20636 8036 20692 8046
rect 20636 7942 20692 7980
rect 20972 7588 21028 7598
rect 20972 7494 21028 7532
rect 21308 7586 21364 8316
rect 21308 7534 21310 7586
rect 21362 7534 21364 7586
rect 21308 7522 21364 7534
rect 20524 7310 20526 7362
rect 20578 7310 20580 7362
rect 20524 7298 20580 7310
rect 19068 6748 19684 6804
rect 18956 6636 19124 6692
rect 18732 6580 18788 6636
rect 18284 6524 18564 6580
rect 18732 6524 19012 6580
rect 18508 6466 18564 6524
rect 18508 6414 18510 6466
rect 18562 6414 18564 6466
rect 18172 6076 18452 6132
rect 16828 6018 17668 6020
rect 16828 5966 16830 6018
rect 16882 5966 17668 6018
rect 16828 5964 17668 5966
rect 16828 5954 16884 5964
rect 16716 5842 16772 5852
rect 17612 5794 17668 5964
rect 18396 6020 18452 6076
rect 18396 5926 18452 5964
rect 17724 5908 17780 5918
rect 18508 5908 18564 6414
rect 18620 6468 18676 6478
rect 18620 6466 18900 6468
rect 18620 6414 18622 6466
rect 18674 6414 18900 6466
rect 18620 6412 18900 6414
rect 18620 6402 18676 6412
rect 18844 6132 18900 6412
rect 18732 5908 18788 5918
rect 18508 5906 18788 5908
rect 18508 5854 18734 5906
rect 18786 5854 18788 5906
rect 18508 5852 18788 5854
rect 17724 5814 17780 5852
rect 18732 5842 18788 5852
rect 17612 5742 17614 5794
rect 17666 5742 17668 5794
rect 17612 5730 17668 5742
rect 17276 5684 17332 5694
rect 17276 5122 17332 5628
rect 17276 5070 17278 5122
rect 17330 5070 17332 5122
rect 17276 5058 17332 5070
rect 17948 5236 18004 5246
rect 16156 4958 16158 5010
rect 16210 4958 16212 5010
rect 16156 4946 16212 4958
rect 17948 5010 18004 5180
rect 18732 5236 18788 5246
rect 18844 5236 18900 6076
rect 18956 5906 19012 6524
rect 18956 5854 18958 5906
rect 19010 5854 19012 5906
rect 18956 5842 19012 5854
rect 19068 5908 19124 6636
rect 19628 6132 19684 6748
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20300 6132 20356 6142
rect 19628 6076 19796 6132
rect 19068 5842 19124 5852
rect 19180 6020 19236 6030
rect 19180 5906 19236 5964
rect 19180 5854 19182 5906
rect 19234 5854 19236 5906
rect 19180 5842 19236 5854
rect 19628 5684 19684 5694
rect 19292 5682 19684 5684
rect 19292 5630 19630 5682
rect 19682 5630 19684 5682
rect 19292 5628 19684 5630
rect 18956 5348 19012 5358
rect 19292 5348 19348 5628
rect 19628 5618 19684 5628
rect 18956 5346 19348 5348
rect 18956 5294 18958 5346
rect 19010 5294 19348 5346
rect 18956 5292 19348 5294
rect 19404 5348 19460 5358
rect 18956 5282 19012 5292
rect 18732 5234 18900 5236
rect 18732 5182 18734 5234
rect 18786 5182 18900 5234
rect 18732 5180 18900 5182
rect 18732 5170 18788 5180
rect 19292 5124 19348 5134
rect 19404 5124 19460 5292
rect 19292 5122 19460 5124
rect 19292 5070 19294 5122
rect 19346 5070 19460 5122
rect 19292 5068 19460 5070
rect 19292 5058 19348 5068
rect 17948 4958 17950 5010
rect 18002 4958 18004 5010
rect 17948 4946 18004 4958
rect 19740 4900 19796 6076
rect 20300 6038 20356 6076
rect 20860 6018 20916 6030
rect 20860 5966 20862 6018
rect 20914 5966 20916 6018
rect 19852 5908 19908 5918
rect 19852 5122 19908 5852
rect 20412 5908 20468 5918
rect 20636 5908 20692 5918
rect 20412 5906 20692 5908
rect 20412 5854 20414 5906
rect 20466 5854 20638 5906
rect 20690 5854 20692 5906
rect 20412 5852 20692 5854
rect 20412 5842 20468 5852
rect 20636 5842 20692 5852
rect 20860 5908 20916 5966
rect 20860 5842 20916 5852
rect 20972 5906 21028 5918
rect 20972 5854 20974 5906
rect 21026 5854 21028 5906
rect 20300 5684 20356 5694
rect 20300 5590 20356 5628
rect 20524 5348 20580 5358
rect 20972 5348 21028 5854
rect 20580 5292 21028 5348
rect 20524 5234 20580 5292
rect 20524 5182 20526 5234
rect 20578 5182 20580 5234
rect 20524 5170 20580 5182
rect 19852 5070 19854 5122
rect 19906 5070 19908 5122
rect 19852 5058 19908 5070
rect 20748 5124 20804 5134
rect 20748 5030 20804 5068
rect 19628 4844 19796 4900
rect 19628 4564 19684 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19740 4564 19796 4574
rect 19628 4562 19796 4564
rect 19628 4510 19742 4562
rect 19794 4510 19796 4562
rect 19628 4508 19796 4510
rect 19740 4498 19796 4508
rect 14700 4452 14756 4462
rect 14700 4358 14756 4396
rect 14028 4340 14084 4350
rect 14364 4340 14420 4350
rect 14028 4338 14420 4340
rect 14028 4286 14030 4338
rect 14082 4286 14366 4338
rect 14418 4286 14420 4338
rect 14028 4284 14420 4286
rect 14028 4274 14084 4284
rect 14364 4274 14420 4284
rect 11340 4228 11396 4238
rect 8764 3378 8820 3388
rect 10780 3444 10836 3454
rect 11004 3444 11060 3454
rect 10780 3442 11060 3444
rect 10780 3390 10782 3442
rect 10834 3390 11006 3442
rect 11058 3390 11060 3442
rect 10780 3388 11060 3390
rect 10780 800 10836 3388
rect 11004 3378 11060 3388
rect 11340 3442 11396 4172
rect 13468 4228 13524 4238
rect 13468 4134 13524 4172
rect 18956 4226 19012 4238
rect 18956 4174 18958 4226
rect 19010 4174 19012 4226
rect 13692 4116 13748 4126
rect 18956 4116 19012 4174
rect 19180 4228 19236 4238
rect 19180 4226 19348 4228
rect 19180 4174 19182 4226
rect 19234 4174 19348 4226
rect 19180 4172 19348 4174
rect 19180 4162 19236 4172
rect 13692 4114 15092 4116
rect 13692 4062 13694 4114
rect 13746 4062 15092 4114
rect 13692 4060 15092 4062
rect 13692 4050 13748 4060
rect 11340 3390 11342 3442
rect 11394 3390 11396 3442
rect 11340 3378 11396 3390
rect 14812 3444 14868 3454
rect 14812 800 14868 3388
rect 15036 3442 15092 4060
rect 18956 4050 19012 4060
rect 15036 3390 15038 3442
rect 15090 3390 15092 3442
rect 15036 3378 15092 3390
rect 15372 3444 15428 3482
rect 15372 3378 15428 3388
rect 18844 3444 18900 3482
rect 19068 3444 19124 3454
rect 18844 3442 19124 3444
rect 18844 3390 18846 3442
rect 18898 3390 19070 3442
rect 19122 3390 19124 3442
rect 18844 3388 19124 3390
rect 19292 3444 19348 4172
rect 19404 4116 19460 4126
rect 19404 4022 19460 4060
rect 19404 3444 19460 3454
rect 19292 3442 19460 3444
rect 19292 3390 19406 3442
rect 19458 3390 19460 3442
rect 19292 3388 19460 3390
rect 21420 3444 21476 10332
rect 21868 10050 21924 10556
rect 21868 9998 21870 10050
rect 21922 9998 21924 10050
rect 21868 9986 21924 9998
rect 22204 10610 22260 10622
rect 22204 10558 22206 10610
rect 22258 10558 22260 10610
rect 22204 10050 22260 10558
rect 22204 9998 22206 10050
rect 22258 9998 22260 10050
rect 22204 9986 22260 9998
rect 21644 9716 21700 9726
rect 21644 9622 21700 9660
rect 21756 8372 21812 8382
rect 21756 8260 21812 8316
rect 21644 8258 21812 8260
rect 21644 8206 21758 8258
rect 21810 8206 21812 8258
rect 21644 8204 21812 8206
rect 21644 7474 21700 8204
rect 21756 8194 21812 8204
rect 21868 8370 21924 8382
rect 21868 8318 21870 8370
rect 21922 8318 21924 8370
rect 21868 7588 21924 8318
rect 22428 8372 22484 13916
rect 22876 13906 22932 13918
rect 22764 13858 22820 13870
rect 22764 13806 22766 13858
rect 22818 13806 22820 13858
rect 22540 13746 22596 13758
rect 22540 13694 22542 13746
rect 22594 13694 22596 13746
rect 22540 12740 22596 13694
rect 22540 12674 22596 12684
rect 22764 13748 22820 13806
rect 22988 13748 23044 19964
rect 23212 20018 23268 20076
rect 23212 19966 23214 20018
rect 23266 19966 23268 20018
rect 23212 19954 23268 19966
rect 23100 19012 23156 19022
rect 23100 19010 23268 19012
rect 23100 18958 23102 19010
rect 23154 18958 23268 19010
rect 23100 18956 23268 18958
rect 23100 18946 23156 18956
rect 23100 16212 23156 16222
rect 23100 16118 23156 16156
rect 22764 13692 23044 13748
rect 22764 11732 22820 13692
rect 22764 11666 22820 11676
rect 22764 11394 22820 11406
rect 23212 11396 23268 18956
rect 23324 15652 23380 22204
rect 23436 18900 23492 24556
rect 23548 23938 23604 23950
rect 23548 23886 23550 23938
rect 23602 23886 23604 23938
rect 23548 23828 23604 23886
rect 23660 23940 23716 24892
rect 24108 24388 24164 26014
rect 24108 24322 24164 24332
rect 23884 23940 23940 23950
rect 23660 23938 23940 23940
rect 23660 23886 23886 23938
rect 23938 23886 23940 23938
rect 23660 23884 23940 23886
rect 23884 23874 23940 23884
rect 23604 23772 23828 23828
rect 23548 23762 23604 23772
rect 23772 23268 23828 23772
rect 23996 23716 24052 23726
rect 23996 23378 24052 23660
rect 23996 23326 23998 23378
rect 24050 23326 24052 23378
rect 23996 23314 24052 23326
rect 24220 23604 24276 26852
rect 23884 23268 23940 23278
rect 23772 23266 23940 23268
rect 23772 23214 23886 23266
rect 23938 23214 23940 23266
rect 23772 23212 23940 23214
rect 23884 23202 23940 23212
rect 24220 23154 24276 23548
rect 24220 23102 24222 23154
rect 24274 23102 24276 23154
rect 24220 23090 24276 23102
rect 24220 20132 24276 20142
rect 24220 20038 24276 20076
rect 23996 19348 24052 19358
rect 23996 19254 24052 19292
rect 23436 18834 23492 18844
rect 23548 19234 23604 19246
rect 23548 19182 23550 19234
rect 23602 19182 23604 19234
rect 23436 15876 23492 15886
rect 23436 15782 23492 15820
rect 23324 15596 23492 15652
rect 23324 15316 23380 15326
rect 23324 14530 23380 15260
rect 23324 14478 23326 14530
rect 23378 14478 23380 14530
rect 23324 14466 23380 14478
rect 23436 13970 23492 15596
rect 23548 14532 23604 19182
rect 24332 18452 24388 18462
rect 23772 15876 23828 15886
rect 24332 15876 24388 18396
rect 24444 17668 24500 17678
rect 24444 16210 24500 17612
rect 24556 16322 24612 26852
rect 24556 16270 24558 16322
rect 24610 16270 24612 16322
rect 24556 16258 24612 16270
rect 24668 18338 24724 18350
rect 24668 18286 24670 18338
rect 24722 18286 24724 18338
rect 24668 16324 24724 18286
rect 24668 16258 24724 16268
rect 24444 16158 24446 16210
rect 24498 16158 24500 16210
rect 24444 16146 24500 16158
rect 23772 15874 24388 15876
rect 23772 15822 23774 15874
rect 23826 15822 24388 15874
rect 23772 15820 24388 15822
rect 23772 15810 23828 15820
rect 24332 15538 24388 15820
rect 24332 15486 24334 15538
rect 24386 15486 24388 15538
rect 24332 15474 24388 15486
rect 24444 15540 24500 15550
rect 24444 15426 24500 15484
rect 24444 15374 24446 15426
rect 24498 15374 24500 15426
rect 24444 15362 24500 15374
rect 24108 15316 24164 15326
rect 24108 15222 24164 15260
rect 23548 14466 23604 14476
rect 24668 14308 24724 14318
rect 23436 13918 23438 13970
rect 23490 13918 23492 13970
rect 23436 13748 23492 13918
rect 23996 13970 24052 13982
rect 23996 13918 23998 13970
rect 24050 13918 24052 13970
rect 23996 13860 24052 13918
rect 23996 13794 24052 13804
rect 23436 13682 23492 13692
rect 23548 13746 23604 13758
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 23436 13524 23492 13534
rect 23548 13524 23604 13694
rect 24108 13748 24164 13758
rect 24108 13654 24164 13692
rect 24556 13748 24612 13758
rect 24444 13634 24500 13646
rect 24444 13582 24446 13634
rect 24498 13582 24500 13634
rect 24444 13524 24500 13582
rect 23548 13468 24500 13524
rect 23436 13430 23492 13468
rect 24444 13074 24500 13468
rect 24444 13022 24446 13074
rect 24498 13022 24500 13074
rect 23772 11844 23828 11854
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 10724 22820 11342
rect 22764 10498 22820 10668
rect 22876 11394 23268 11396
rect 22876 11342 23214 11394
rect 23266 11342 23268 11394
rect 22876 11340 23268 11342
rect 22876 10610 22932 11340
rect 23212 11330 23268 11340
rect 23660 11732 23716 11742
rect 23660 10834 23716 11676
rect 23660 10782 23662 10834
rect 23714 10782 23716 10834
rect 23660 10770 23716 10782
rect 23212 10724 23268 10734
rect 23212 10722 23492 10724
rect 23212 10670 23214 10722
rect 23266 10670 23492 10722
rect 23212 10668 23492 10670
rect 23212 10658 23268 10668
rect 22876 10558 22878 10610
rect 22930 10558 22932 10610
rect 22876 10546 22932 10558
rect 22764 10446 22766 10498
rect 22818 10446 22820 10498
rect 22764 10434 22820 10446
rect 23436 8428 23492 10668
rect 23772 10722 23828 11788
rect 24332 11508 24388 11518
rect 24444 11508 24500 13022
rect 24556 12962 24612 13692
rect 24556 12910 24558 12962
rect 24610 12910 24612 12962
rect 24556 12898 24612 12910
rect 24332 11506 24500 11508
rect 24332 11454 24334 11506
rect 24386 11454 24500 11506
rect 24332 11452 24500 11454
rect 24332 11442 24388 11452
rect 24668 11396 24724 14252
rect 23772 10670 23774 10722
rect 23826 10670 23828 10722
rect 23772 10658 23828 10670
rect 24444 11394 24724 11396
rect 24444 11342 24670 11394
rect 24722 11342 24724 11394
rect 24444 11340 24724 11342
rect 24444 10722 24500 11340
rect 24668 11330 24724 11340
rect 24556 11172 24612 11182
rect 24556 10834 24612 11116
rect 24780 11060 24836 31276
rect 24892 29652 24948 29662
rect 24892 20132 24948 29596
rect 25004 26180 25060 36206
rect 25004 26114 25060 26124
rect 25116 24052 25172 39788
rect 25228 38946 25284 40124
rect 25340 39618 25396 40348
rect 25340 39566 25342 39618
rect 25394 39566 25396 39618
rect 25340 39554 25396 39566
rect 25228 38894 25230 38946
rect 25282 38894 25284 38946
rect 25228 38882 25284 38894
rect 25340 38722 25396 38734
rect 25340 38670 25342 38722
rect 25394 38670 25396 38722
rect 25340 33458 25396 38670
rect 25452 36372 25508 40572
rect 25564 40516 25620 42812
rect 25676 42642 25732 42654
rect 25676 42590 25678 42642
rect 25730 42590 25732 42642
rect 25676 42420 25732 42590
rect 25676 42354 25732 42364
rect 25788 41972 25844 43486
rect 26124 42308 26180 45948
rect 26236 45780 26292 45790
rect 26572 45780 26628 46620
rect 26796 46610 26852 46620
rect 26908 47180 27188 47236
rect 26236 45686 26292 45724
rect 26348 45778 26628 45780
rect 26348 45726 26574 45778
rect 26626 45726 26628 45778
rect 26348 45724 26628 45726
rect 26348 45106 26404 45724
rect 26572 45714 26628 45724
rect 26684 46452 26740 46462
rect 26908 46452 26964 47180
rect 27468 46788 27524 50540
rect 27580 47348 27636 53564
rect 27580 47282 27636 47292
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 26348 45042 26404 45054
rect 26236 44098 26292 44110
rect 26236 44046 26238 44098
rect 26290 44046 26292 44098
rect 26236 43764 26292 44046
rect 26236 43698 26292 43708
rect 26460 43538 26516 43550
rect 26460 43486 26462 43538
rect 26514 43486 26516 43538
rect 26236 42756 26292 42766
rect 26236 42662 26292 42700
rect 26124 42252 26404 42308
rect 25788 41970 25956 41972
rect 25788 41918 25790 41970
rect 25842 41918 25956 41970
rect 25788 41916 25956 41918
rect 25788 41906 25844 41916
rect 25564 40450 25620 40460
rect 25788 40402 25844 40414
rect 25788 40350 25790 40402
rect 25842 40350 25844 40402
rect 25788 39172 25844 40350
rect 25900 39618 25956 41916
rect 25900 39566 25902 39618
rect 25954 39566 25956 39618
rect 25900 39554 25956 39566
rect 25788 39106 25844 39116
rect 26012 39506 26068 39518
rect 26012 39454 26014 39506
rect 26066 39454 26068 39506
rect 25564 38946 25620 38958
rect 25564 38894 25566 38946
rect 25618 38894 25620 38946
rect 25564 38836 25620 38894
rect 25788 38948 25844 38958
rect 25788 38854 25844 38892
rect 25676 38836 25732 38846
rect 25564 38780 25676 38836
rect 25676 38770 25732 38780
rect 25564 37828 25620 37838
rect 25564 37734 25620 37772
rect 25676 36484 25732 36494
rect 25676 36390 25732 36428
rect 25452 36316 25620 36372
rect 25452 34132 25508 34142
rect 25452 34038 25508 34076
rect 25564 34018 25620 36316
rect 25900 35586 25956 35598
rect 25900 35534 25902 35586
rect 25954 35534 25956 35586
rect 25788 35474 25844 35486
rect 25788 35422 25790 35474
rect 25842 35422 25844 35474
rect 25788 34914 25844 35422
rect 25788 34862 25790 34914
rect 25842 34862 25844 34914
rect 25788 34850 25844 34862
rect 25900 34916 25956 35534
rect 25900 34132 25956 34860
rect 25564 33966 25566 34018
rect 25618 33966 25620 34018
rect 25564 33954 25620 33966
rect 25676 34076 25956 34132
rect 25340 33406 25342 33458
rect 25394 33406 25396 33458
rect 25340 33394 25396 33406
rect 25228 32562 25284 32574
rect 25228 32510 25230 32562
rect 25282 32510 25284 32562
rect 25228 32452 25284 32510
rect 25228 32386 25284 32396
rect 25564 30994 25620 31006
rect 25564 30942 25566 30994
rect 25618 30942 25620 30994
rect 25452 29652 25508 29662
rect 25452 29426 25508 29596
rect 25564 29540 25620 30942
rect 25676 30996 25732 34076
rect 25900 33908 25956 33918
rect 25900 33814 25956 33852
rect 26012 32788 26068 39454
rect 26236 38948 26292 38958
rect 26124 38834 26180 38846
rect 26124 38782 26126 38834
rect 26178 38782 26180 38834
rect 26124 38052 26180 38782
rect 26124 37986 26180 37996
rect 26124 37156 26180 37166
rect 26124 37062 26180 37100
rect 26236 36482 26292 38892
rect 26348 38668 26404 42252
rect 26460 41972 26516 43486
rect 26684 42756 26740 46396
rect 26684 42690 26740 42700
rect 26796 46396 26964 46452
rect 27356 46732 27524 46788
rect 26796 42196 26852 46396
rect 26908 46004 26964 46014
rect 26908 45890 26964 45948
rect 26908 45838 26910 45890
rect 26962 45838 26964 45890
rect 26908 45826 26964 45838
rect 27132 45220 27188 45230
rect 27132 45126 27188 45164
rect 27020 43540 27076 43550
rect 26908 42980 26964 42990
rect 26908 42754 26964 42924
rect 27020 42978 27076 43484
rect 27244 43428 27300 43438
rect 27244 43334 27300 43372
rect 27020 42926 27022 42978
rect 27074 42926 27076 42978
rect 27020 42914 27076 42926
rect 27356 42756 27412 46732
rect 27468 46564 27524 46574
rect 27468 46470 27524 46508
rect 27692 43764 27748 55804
rect 27804 50428 27860 56364
rect 28028 55412 28084 55422
rect 28028 55318 28084 55356
rect 27916 55188 27972 55198
rect 27916 53844 27972 55132
rect 28364 54852 28420 56700
rect 28476 56308 28532 56318
rect 28476 56214 28532 56252
rect 27916 53618 27972 53788
rect 27916 53566 27918 53618
rect 27970 53566 27972 53618
rect 27916 53284 27972 53566
rect 27916 53218 27972 53228
rect 28028 54796 28420 54852
rect 28476 55188 28532 55198
rect 28028 52836 28084 54796
rect 28140 54516 28196 54526
rect 28140 54402 28196 54460
rect 28476 54514 28532 55132
rect 28476 54462 28478 54514
rect 28530 54462 28532 54514
rect 28476 54450 28532 54462
rect 28140 54350 28142 54402
rect 28194 54350 28196 54402
rect 28140 54068 28196 54350
rect 28140 54002 28196 54012
rect 28252 53620 28308 53630
rect 28308 53564 28420 53620
rect 28252 53554 28308 53564
rect 28140 53508 28196 53518
rect 28140 53058 28196 53452
rect 28364 53506 28420 53564
rect 28364 53454 28366 53506
rect 28418 53454 28420 53506
rect 28364 53442 28420 53454
rect 28140 53006 28142 53058
rect 28194 53006 28196 53058
rect 28140 52994 28196 53006
rect 28028 52780 28196 52836
rect 28028 51378 28084 51390
rect 28028 51326 28030 51378
rect 28082 51326 28084 51378
rect 28028 50484 28084 51326
rect 27804 50372 27972 50428
rect 28028 50418 28084 50428
rect 28140 50428 28196 52780
rect 28476 52276 28532 52286
rect 28476 52162 28532 52220
rect 28476 52110 28478 52162
rect 28530 52110 28532 52162
rect 28476 52098 28532 52110
rect 28252 51378 28308 51390
rect 28252 51326 28254 51378
rect 28306 51326 28308 51378
rect 28252 50820 28308 51326
rect 28476 51268 28532 51278
rect 28252 50754 28308 50764
rect 28364 51212 28476 51268
rect 28364 50596 28420 51212
rect 28476 51202 28532 51212
rect 28588 50932 28644 58156
rect 28700 57652 28756 57662
rect 28700 56194 28756 57596
rect 28700 56142 28702 56194
rect 28754 56142 28756 56194
rect 28700 52724 28756 56142
rect 28700 52658 28756 52668
rect 28812 51492 28868 60060
rect 28924 57540 28980 57550
rect 28924 57446 28980 57484
rect 29036 56420 29092 63980
rect 29260 63812 29316 63822
rect 29260 63718 29316 63756
rect 29372 63810 29428 63822
rect 29372 63758 29374 63810
rect 29426 63758 29428 63810
rect 29372 63252 29428 63758
rect 29484 63700 29540 65996
rect 29820 64820 29876 66220
rect 29596 64818 29876 64820
rect 29596 64766 29822 64818
rect 29874 64766 29876 64818
rect 29596 64764 29876 64766
rect 29596 63922 29652 64764
rect 29820 64754 29876 64764
rect 29932 66274 29988 66286
rect 29932 66222 29934 66274
rect 29986 66222 29988 66274
rect 29932 66052 29988 66222
rect 29596 63870 29598 63922
rect 29650 63870 29652 63922
rect 29596 63858 29652 63870
rect 29932 63812 29988 65996
rect 30044 65604 30100 67790
rect 30156 67228 30212 69468
rect 30940 67844 30996 67854
rect 30716 67618 30772 67630
rect 30716 67566 30718 67618
rect 30770 67566 30772 67618
rect 30716 67228 30772 67566
rect 30156 67172 30324 67228
rect 30268 67058 30324 67172
rect 30268 67006 30270 67058
rect 30322 67006 30324 67058
rect 30268 66994 30324 67006
rect 30604 67172 30884 67228
rect 30604 66836 30660 67172
rect 30828 67170 30884 67172
rect 30828 67118 30830 67170
rect 30882 67118 30884 67170
rect 30828 67106 30884 67118
rect 30604 66770 30660 66780
rect 30716 67058 30772 67070
rect 30716 67006 30718 67058
rect 30770 67006 30772 67058
rect 30716 66612 30772 67006
rect 30156 66556 30772 66612
rect 30828 66948 30884 66958
rect 30940 66948 30996 67788
rect 30828 66946 30996 66948
rect 30828 66894 30830 66946
rect 30882 66894 30996 66946
rect 30828 66892 30996 66894
rect 31052 67618 31108 67630
rect 31052 67566 31054 67618
rect 31106 67566 31108 67618
rect 31052 67508 31108 67566
rect 31724 67620 31780 67630
rect 31724 67526 31780 67564
rect 30156 66386 30212 66556
rect 30156 66334 30158 66386
rect 30210 66334 30212 66386
rect 30156 66322 30212 66334
rect 30604 66276 30660 66286
rect 30604 66182 30660 66220
rect 30044 65548 30324 65604
rect 30268 65380 30324 65548
rect 30604 65492 30660 65502
rect 30828 65492 30884 66892
rect 31052 66052 31108 67452
rect 32172 67228 32228 71822
rect 32284 72156 32676 72212
rect 32732 72212 32788 72222
rect 32284 71874 32340 72156
rect 32284 71822 32286 71874
rect 32338 71822 32340 71874
rect 32284 71810 32340 71822
rect 32508 71204 32564 71214
rect 32732 71204 32788 72156
rect 33852 71762 33908 71774
rect 33852 71710 33854 71762
rect 33906 71710 33908 71762
rect 33180 71652 33236 71662
rect 32508 71202 32788 71204
rect 32508 71150 32510 71202
rect 32562 71150 32788 71202
rect 32508 71148 32788 71150
rect 33068 71650 33236 71652
rect 33068 71598 33182 71650
rect 33234 71598 33236 71650
rect 33068 71596 33236 71598
rect 32508 71138 32564 71148
rect 32956 70980 33012 70990
rect 33068 70980 33124 71596
rect 33180 71586 33236 71596
rect 32956 70978 33124 70980
rect 32956 70926 32958 70978
rect 33010 70926 33124 70978
rect 32956 70924 33124 70926
rect 33180 70980 33236 70990
rect 33180 70978 33348 70980
rect 33180 70926 33182 70978
rect 33234 70926 33348 70978
rect 33180 70924 33348 70926
rect 32956 70194 33012 70924
rect 33180 70914 33236 70924
rect 33292 70308 33348 70924
rect 33404 70978 33460 70990
rect 33404 70926 33406 70978
rect 33458 70926 33460 70978
rect 33404 70420 33460 70926
rect 33852 70644 33908 71710
rect 33852 70578 33908 70588
rect 33964 70978 34020 72492
rect 34076 72482 34132 72492
rect 35084 71762 35140 71774
rect 35084 71710 35086 71762
rect 35138 71710 35140 71762
rect 34076 71650 34132 71662
rect 34076 71598 34078 71650
rect 34130 71598 34132 71650
rect 34076 71092 34132 71598
rect 34972 71652 35028 71662
rect 34076 71026 34132 71036
rect 34860 71092 34916 71102
rect 33964 70926 33966 70978
rect 34018 70926 34020 70978
rect 33404 70364 33796 70420
rect 33292 70252 33684 70308
rect 32956 70142 32958 70194
rect 33010 70142 33012 70194
rect 32956 70130 33012 70142
rect 33404 69634 33460 70252
rect 33628 70082 33684 70252
rect 33628 70030 33630 70082
rect 33682 70030 33684 70082
rect 33628 70018 33684 70030
rect 33740 70194 33796 70364
rect 33964 70306 34020 70926
rect 34860 70978 34916 71036
rect 34860 70926 34862 70978
rect 34914 70926 34916 70978
rect 34860 70914 34916 70926
rect 33964 70254 33966 70306
rect 34018 70254 34020 70306
rect 33964 70242 34020 70254
rect 34076 70644 34132 70654
rect 33740 70142 33742 70194
rect 33794 70142 33796 70194
rect 33404 69582 33406 69634
rect 33458 69582 33460 69634
rect 33404 69570 33460 69582
rect 33404 69410 33460 69422
rect 33404 69358 33406 69410
rect 33458 69358 33460 69410
rect 33068 69298 33124 69310
rect 33068 69246 33070 69298
rect 33122 69246 33124 69298
rect 33068 68628 33124 69246
rect 33404 68740 33460 69358
rect 33740 68850 33796 70142
rect 33740 68798 33742 68850
rect 33794 68798 33796 68850
rect 33740 68786 33796 68798
rect 33404 68674 33460 68684
rect 32396 68516 32452 68526
rect 32396 67842 32452 68460
rect 32396 67790 32398 67842
rect 32450 67790 32452 67842
rect 32396 67620 32452 67790
rect 32956 67842 33012 67854
rect 32956 67790 32958 67842
rect 33010 67790 33012 67842
rect 32956 67732 33012 67790
rect 32956 67666 33012 67676
rect 33068 67730 33124 68572
rect 33628 68626 33684 68638
rect 33628 68574 33630 68626
rect 33682 68574 33684 68626
rect 33068 67678 33070 67730
rect 33122 67678 33124 67730
rect 33068 67666 33124 67678
rect 33404 67732 33460 67742
rect 33404 67638 33460 67676
rect 32396 67554 32452 67564
rect 33628 67228 33684 68574
rect 34076 67954 34132 70588
rect 34972 70418 35028 71596
rect 34972 70366 34974 70418
rect 35026 70366 35028 70418
rect 34972 70354 35028 70366
rect 35084 70418 35140 71710
rect 35644 71762 35700 71774
rect 35644 71710 35646 71762
rect 35698 71710 35700 71762
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35084 70366 35086 70418
rect 35138 70366 35140 70418
rect 35084 70354 35140 70366
rect 35532 71092 35588 71102
rect 35532 70306 35588 71036
rect 35644 70868 35700 71710
rect 35868 71762 35924 71774
rect 35868 71710 35870 71762
rect 35922 71710 35924 71762
rect 35644 70802 35700 70812
rect 35756 71650 35812 71662
rect 35756 71598 35758 71650
rect 35810 71598 35812 71650
rect 35532 70254 35534 70306
rect 35586 70254 35588 70306
rect 35532 70242 35588 70254
rect 35196 69972 35252 69982
rect 35196 69970 35588 69972
rect 35196 69918 35198 69970
rect 35250 69918 35588 69970
rect 35196 69916 35588 69918
rect 35196 69906 35252 69916
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35532 69524 35588 69916
rect 35644 69524 35700 69534
rect 35532 69468 35644 69524
rect 35644 69430 35700 69468
rect 35196 69188 35252 69198
rect 35196 69094 35252 69132
rect 34300 68740 34356 68750
rect 35756 68740 35812 71598
rect 35868 71204 35924 71710
rect 35868 71110 35924 71148
rect 37100 71762 37156 71774
rect 37100 71710 37102 71762
rect 37154 71710 37156 71762
rect 35980 70978 36036 70990
rect 35980 70926 35982 70978
rect 36034 70926 36036 70978
rect 35980 70644 36036 70926
rect 36988 70868 37044 70878
rect 36988 70774 37044 70812
rect 35980 70578 36036 70588
rect 36876 70196 36932 70206
rect 37100 70196 37156 71710
rect 37548 71764 37604 71774
rect 37548 71762 37716 71764
rect 37548 71710 37550 71762
rect 37602 71710 37716 71762
rect 37548 71708 37716 71710
rect 37548 71698 37604 71708
rect 37324 71652 37380 71662
rect 37324 71558 37380 71596
rect 36876 70194 37156 70196
rect 36876 70142 36878 70194
rect 36930 70142 37156 70194
rect 36876 70140 37156 70142
rect 37660 70194 37716 71708
rect 37772 71762 37828 71774
rect 37772 71710 37774 71762
rect 37826 71710 37828 71762
rect 37772 70532 37828 71710
rect 37996 71652 38052 71662
rect 37996 70978 38052 71596
rect 37996 70926 37998 70978
rect 38050 70926 38052 70978
rect 37996 70914 38052 70926
rect 38556 70978 38612 70990
rect 38556 70926 38558 70978
rect 38610 70926 38612 70978
rect 38556 70756 38612 70926
rect 39116 70756 39172 70766
rect 38556 70754 39172 70756
rect 38556 70702 39118 70754
rect 39170 70702 39172 70754
rect 38556 70700 39172 70702
rect 37772 70466 37828 70476
rect 38892 70532 38948 70542
rect 38892 70418 38948 70476
rect 38892 70366 38894 70418
rect 38946 70366 38948 70418
rect 38892 70354 38948 70366
rect 37660 70142 37662 70194
rect 37714 70142 37716 70194
rect 36428 70084 36484 70094
rect 36428 69634 36484 70028
rect 36428 69582 36430 69634
rect 36482 69582 36484 69634
rect 36428 69570 36484 69582
rect 34188 68628 34244 68638
rect 34188 68534 34244 68572
rect 34076 67902 34078 67954
rect 34130 67902 34132 67954
rect 34076 67890 34132 67902
rect 32172 67172 32340 67228
rect 31836 66946 31892 66958
rect 31836 66894 31838 66946
rect 31890 66894 31892 66946
rect 31836 66388 31892 66894
rect 31052 65958 31108 65996
rect 31276 66276 31332 66286
rect 30604 65490 30884 65492
rect 30604 65438 30606 65490
rect 30658 65438 30884 65490
rect 30604 65436 30884 65438
rect 30604 65426 30660 65436
rect 30492 65380 30548 65390
rect 30268 65378 30548 65380
rect 30268 65326 30494 65378
rect 30546 65326 30548 65378
rect 30268 65324 30548 65326
rect 30156 65266 30212 65278
rect 30156 65214 30158 65266
rect 30210 65214 30212 65266
rect 29932 63746 29988 63756
rect 30044 63810 30100 63822
rect 30044 63758 30046 63810
rect 30098 63758 30100 63810
rect 29484 63644 29764 63700
rect 29372 63250 29652 63252
rect 29372 63198 29374 63250
rect 29426 63198 29652 63250
rect 29372 63196 29652 63198
rect 29372 63186 29428 63196
rect 29484 63028 29540 63038
rect 29484 62934 29540 62972
rect 29372 62916 29428 62926
rect 29148 62860 29372 62916
rect 29148 62354 29204 62860
rect 29372 62850 29428 62860
rect 29148 62302 29150 62354
rect 29202 62302 29204 62354
rect 29148 62290 29204 62302
rect 29372 62132 29428 62142
rect 29260 60676 29316 60686
rect 29260 60582 29316 60620
rect 29260 58322 29316 58334
rect 29260 58270 29262 58322
rect 29314 58270 29316 58322
rect 29148 58212 29204 58222
rect 29260 58212 29316 58270
rect 29204 58156 29316 58212
rect 29148 58146 29204 58156
rect 29260 56868 29316 56878
rect 29260 56774 29316 56812
rect 29036 56082 29092 56364
rect 29036 56030 29038 56082
rect 29090 56030 29092 56082
rect 29036 56018 29092 56030
rect 29260 54404 29316 54414
rect 29260 54310 29316 54348
rect 29148 53844 29204 53854
rect 29148 53730 29204 53788
rect 29148 53678 29150 53730
rect 29202 53678 29204 53730
rect 29148 53666 29204 53678
rect 29372 53508 29428 62076
rect 29484 61794 29540 61806
rect 29484 61742 29486 61794
rect 29538 61742 29540 61794
rect 29484 60786 29540 61742
rect 29596 61570 29652 63196
rect 29596 61518 29598 61570
rect 29650 61518 29652 61570
rect 29596 61506 29652 61518
rect 29484 60734 29486 60786
rect 29538 60734 29540 60786
rect 29484 60722 29540 60734
rect 29708 58772 29764 63644
rect 30044 62916 30100 63758
rect 30156 63812 30212 65214
rect 30492 65156 30548 65324
rect 30492 65100 30660 65156
rect 30268 64484 30324 64494
rect 30268 64482 30436 64484
rect 30268 64430 30270 64482
rect 30322 64430 30436 64482
rect 30268 64428 30436 64430
rect 30268 64418 30324 64428
rect 30268 63812 30324 63822
rect 30156 63810 30324 63812
rect 30156 63758 30270 63810
rect 30322 63758 30324 63810
rect 30156 63756 30324 63758
rect 29820 62860 30044 62916
rect 29820 61010 29876 62860
rect 30044 62850 30100 62860
rect 30268 62354 30324 63756
rect 30268 62302 30270 62354
rect 30322 62302 30324 62354
rect 30268 62290 30324 62302
rect 30380 63812 30436 64428
rect 29932 61684 29988 61694
rect 29932 61590 29988 61628
rect 29820 60958 29822 61010
rect 29874 60958 29876 61010
rect 29820 60946 29876 60958
rect 29932 59108 29988 59118
rect 29932 59106 30100 59108
rect 29932 59054 29934 59106
rect 29986 59054 30100 59106
rect 29932 59052 30100 59054
rect 29932 59042 29988 59052
rect 29708 58716 29988 58772
rect 29820 58548 29876 58558
rect 29708 58546 29876 58548
rect 29708 58494 29822 58546
rect 29874 58494 29876 58546
rect 29708 58492 29876 58494
rect 29596 58212 29652 58222
rect 29708 58212 29764 58492
rect 29820 58482 29876 58492
rect 29652 58156 29764 58212
rect 29596 58146 29652 58156
rect 29708 57650 29764 58156
rect 29708 57598 29710 57650
rect 29762 57598 29764 57650
rect 29708 57586 29764 57598
rect 29148 53452 29428 53508
rect 29596 57538 29652 57550
rect 29932 57540 29988 58716
rect 29596 57486 29598 57538
rect 29650 57486 29652 57538
rect 28812 51426 28868 51436
rect 29036 51716 29092 51726
rect 29036 51378 29092 51660
rect 29036 51326 29038 51378
rect 29090 51326 29092 51378
rect 29036 51314 29092 51326
rect 28924 51266 28980 51278
rect 28924 51214 28926 51266
rect 28978 51214 28980 51266
rect 28812 51156 28868 51166
rect 28812 51062 28868 51100
rect 28588 50876 28868 50932
rect 28364 50530 28420 50540
rect 28140 50372 28420 50428
rect 27804 49810 27860 49822
rect 27804 49758 27806 49810
rect 27858 49758 27860 49810
rect 27804 49028 27860 49758
rect 27804 48962 27860 48972
rect 27804 48804 27860 48814
rect 27804 48710 27860 48748
rect 26908 42702 26910 42754
rect 26962 42702 26964 42754
rect 26908 42690 26964 42702
rect 27020 42700 27412 42756
rect 27020 42642 27076 42700
rect 27020 42590 27022 42642
rect 27074 42590 27076 42642
rect 27020 42578 27076 42590
rect 26796 42140 26964 42196
rect 26460 40740 26516 41916
rect 26684 41972 26740 41982
rect 26684 41878 26740 41916
rect 26908 41076 26964 42140
rect 27356 41972 27412 42700
rect 27356 41906 27412 41916
rect 27580 43708 27748 43764
rect 27468 41860 27524 41870
rect 27468 41766 27524 41804
rect 26908 41010 26964 41020
rect 26460 40674 26516 40684
rect 26460 40516 26516 40526
rect 26516 40460 26628 40516
rect 26460 40450 26516 40460
rect 26572 40402 26628 40460
rect 26572 40350 26574 40402
rect 26626 40350 26628 40402
rect 26572 40338 26628 40350
rect 26796 38948 26852 38958
rect 26460 38836 26516 38874
rect 26796 38854 26852 38892
rect 26460 38770 26516 38780
rect 26348 38612 26516 38668
rect 26236 36430 26238 36482
rect 26290 36430 26292 36482
rect 26236 35476 26292 36430
rect 26236 35410 26292 35420
rect 26348 36932 26404 36942
rect 26348 35922 26404 36876
rect 26348 35870 26350 35922
rect 26402 35870 26404 35922
rect 26348 35474 26404 35870
rect 26348 35422 26350 35474
rect 26402 35422 26404 35474
rect 26348 35252 26404 35422
rect 26236 35196 26404 35252
rect 26012 32732 26180 32788
rect 26012 32452 26068 32462
rect 25788 32450 26068 32452
rect 25788 32398 26014 32450
rect 26066 32398 26068 32450
rect 25788 32396 26068 32398
rect 25788 31218 25844 32396
rect 26012 32386 26068 32396
rect 25788 31166 25790 31218
rect 25842 31166 25844 31218
rect 25788 31154 25844 31166
rect 25676 30940 26068 30996
rect 25564 29474 25620 29484
rect 25452 29374 25454 29426
rect 25506 29374 25508 29426
rect 25452 29362 25508 29374
rect 25900 29314 25956 29326
rect 25900 29262 25902 29314
rect 25954 29262 25956 29314
rect 25452 28868 25508 28878
rect 25452 28642 25508 28812
rect 25788 28644 25844 28654
rect 25452 28590 25454 28642
rect 25506 28590 25508 28642
rect 25452 28578 25508 28590
rect 25676 28642 25844 28644
rect 25676 28590 25790 28642
rect 25842 28590 25844 28642
rect 25676 28588 25844 28590
rect 25676 27970 25732 28588
rect 25788 28578 25844 28588
rect 25900 28082 25956 29262
rect 26012 29092 26068 30940
rect 26124 29204 26180 32732
rect 26236 29652 26292 35196
rect 26348 35028 26404 35038
rect 26460 35028 26516 38612
rect 27020 38050 27076 38062
rect 27468 38052 27524 38062
rect 27020 37998 27022 38050
rect 27074 37998 27076 38050
rect 26572 37492 26628 37502
rect 26572 37398 26628 37436
rect 26684 37380 26740 37390
rect 26684 37286 26740 37324
rect 27020 37380 27076 37998
rect 27244 37996 27468 38052
rect 27244 37492 27300 37996
rect 27468 37958 27524 37996
rect 27244 37398 27300 37436
rect 27020 37314 27076 37324
rect 27356 37156 27412 37166
rect 26572 37042 26628 37054
rect 26572 36990 26574 37042
rect 26626 36990 26628 37042
rect 26572 35364 26628 36990
rect 26572 35298 26628 35308
rect 26684 37044 26740 37054
rect 26348 35026 26516 35028
rect 26348 34974 26350 35026
rect 26402 34974 26516 35026
rect 26348 34972 26516 34974
rect 26348 34962 26404 34972
rect 26236 29586 26292 29596
rect 26460 34356 26516 34366
rect 26460 34020 26516 34300
rect 26572 34020 26628 34030
rect 26460 34018 26628 34020
rect 26460 33966 26574 34018
rect 26626 33966 26628 34018
rect 26460 33964 26628 33966
rect 26348 29204 26404 29214
rect 26124 29148 26348 29204
rect 26348 29138 26404 29148
rect 26012 29036 26292 29092
rect 25900 28030 25902 28082
rect 25954 28030 25956 28082
rect 25900 28018 25956 28030
rect 26012 28868 26068 28878
rect 25676 27918 25678 27970
rect 25730 27918 25732 27970
rect 25564 27188 25620 27198
rect 25564 27094 25620 27132
rect 25676 26908 25732 27918
rect 26012 27970 26068 28812
rect 26012 27918 26014 27970
rect 26066 27918 26068 27970
rect 26012 27906 26068 27918
rect 26124 27858 26180 27870
rect 26124 27806 26126 27858
rect 26178 27806 26180 27858
rect 26124 26908 26180 27806
rect 25340 26852 25732 26908
rect 25788 26852 26180 26908
rect 25228 25506 25284 25518
rect 25228 25454 25230 25506
rect 25282 25454 25284 25506
rect 25228 25060 25284 25454
rect 25228 24994 25284 25004
rect 25228 24836 25284 24846
rect 25340 24836 25396 26852
rect 25788 25730 25844 26852
rect 25788 25678 25790 25730
rect 25842 25678 25844 25730
rect 25788 25666 25844 25678
rect 25228 24834 25396 24836
rect 25228 24782 25230 24834
rect 25282 24782 25396 24834
rect 25228 24780 25396 24782
rect 25452 25506 25508 25518
rect 25452 25454 25454 25506
rect 25506 25454 25508 25506
rect 25228 24770 25284 24780
rect 25452 24724 25508 25454
rect 25452 24630 25508 24668
rect 25900 25060 25956 25070
rect 25900 24722 25956 25004
rect 25900 24670 25902 24722
rect 25954 24670 25956 24722
rect 24892 19234 24948 20076
rect 24892 19182 24894 19234
rect 24946 19182 24948 19234
rect 24892 19170 24948 19182
rect 25004 23996 25172 24052
rect 25676 24388 25732 24398
rect 25004 17780 25060 23996
rect 25452 23940 25508 23950
rect 25452 23846 25508 23884
rect 25116 23828 25172 23838
rect 25116 23734 25172 23772
rect 25676 23826 25732 24332
rect 25676 23774 25678 23826
rect 25730 23774 25732 23826
rect 25340 23156 25396 23166
rect 25676 23156 25732 23774
rect 25340 23154 25732 23156
rect 25340 23102 25342 23154
rect 25394 23102 25732 23154
rect 25340 23100 25732 23102
rect 25340 23090 25396 23100
rect 25788 23044 25844 23054
rect 25788 22950 25844 22988
rect 25900 22820 25956 24670
rect 25676 22764 25956 22820
rect 26124 24052 26180 24062
rect 26124 23266 26180 23996
rect 26124 23214 26126 23266
rect 26178 23214 26180 23266
rect 25340 21588 25396 21598
rect 25676 21588 25732 22764
rect 25900 22596 25956 22606
rect 25900 22482 25956 22540
rect 26124 22596 26180 23214
rect 26236 23268 26292 29036
rect 26460 26908 26516 33964
rect 26572 33954 26628 33964
rect 26684 26908 26740 36988
rect 27132 36482 27188 36494
rect 27132 36430 27134 36482
rect 27186 36430 27188 36482
rect 26908 35700 26964 35710
rect 27132 35700 27188 36430
rect 26964 35644 27188 35700
rect 27356 36484 27412 37100
rect 26796 35588 26852 35598
rect 26796 35494 26852 35532
rect 26796 29428 26852 29438
rect 26796 29334 26852 29372
rect 26348 26852 26516 26908
rect 26572 26852 26740 26908
rect 26796 29092 26852 29102
rect 26348 24948 26404 26852
rect 26348 24882 26404 24892
rect 26460 25282 26516 25294
rect 26460 25230 26462 25282
rect 26514 25230 26516 25282
rect 26460 24836 26516 25230
rect 26460 24052 26516 24780
rect 26460 23986 26516 23996
rect 26348 23938 26404 23950
rect 26348 23886 26350 23938
rect 26402 23886 26404 23938
rect 26348 23716 26404 23886
rect 26348 23650 26404 23660
rect 26460 23714 26516 23726
rect 26460 23662 26462 23714
rect 26514 23662 26516 23714
rect 26236 23212 26404 23268
rect 26124 22530 26180 22540
rect 26236 23042 26292 23054
rect 26236 22990 26238 23042
rect 26290 22990 26292 23042
rect 25900 22430 25902 22482
rect 25954 22430 25956 22482
rect 25900 22418 25956 22430
rect 26236 22372 26292 22990
rect 26236 22036 26292 22316
rect 25340 21586 25732 21588
rect 25340 21534 25342 21586
rect 25394 21534 25732 21586
rect 25340 21532 25732 21534
rect 26012 21980 26292 22036
rect 25228 20916 25284 20926
rect 25228 20822 25284 20860
rect 25228 19908 25284 19918
rect 25228 19814 25284 19852
rect 25340 19684 25396 21532
rect 25788 21474 25844 21486
rect 25788 21422 25790 21474
rect 25842 21422 25844 21474
rect 25788 20916 25844 21422
rect 25788 20850 25844 20860
rect 25900 20804 25956 20814
rect 26012 20804 26068 21980
rect 26124 21700 26180 21710
rect 26124 21606 26180 21644
rect 26236 21028 26292 21038
rect 25900 20802 26068 20804
rect 25900 20750 25902 20802
rect 25954 20750 26068 20802
rect 25900 20748 26068 20750
rect 26124 20804 26180 20814
rect 25900 20738 25956 20748
rect 26124 20710 26180 20748
rect 25676 20580 25732 20590
rect 25676 20486 25732 20524
rect 26012 20578 26068 20590
rect 26012 20526 26014 20578
rect 26066 20526 26068 20578
rect 25228 19628 25396 19684
rect 25564 20132 25620 20142
rect 25228 18452 25284 19628
rect 25564 19346 25620 20076
rect 26012 20130 26068 20526
rect 26012 20078 26014 20130
rect 26066 20078 26068 20130
rect 26012 20066 26068 20078
rect 25564 19294 25566 19346
rect 25618 19294 25620 19346
rect 25564 19282 25620 19294
rect 26236 19348 26292 20972
rect 26348 19460 26404 23212
rect 26460 19796 26516 23662
rect 26572 21028 26628 26852
rect 26684 23156 26740 23166
rect 26684 23062 26740 23100
rect 26572 20962 26628 20972
rect 26460 19740 26740 19796
rect 26348 19404 26628 19460
rect 26236 19292 26516 19348
rect 25452 19236 25508 19246
rect 25452 19142 25508 19180
rect 26124 19236 26180 19246
rect 26124 19142 26180 19180
rect 25228 18386 25284 18396
rect 26236 18452 26292 18462
rect 25340 18340 25396 18350
rect 25340 18246 25396 18284
rect 25004 17714 25060 17724
rect 26236 17778 26292 18396
rect 26236 17726 26238 17778
rect 26290 17726 26292 17778
rect 25116 17668 25172 17678
rect 24892 16322 24948 16334
rect 24892 16270 24894 16322
rect 24946 16270 24948 16322
rect 24892 16212 24948 16270
rect 24892 16118 24948 16156
rect 25116 16098 25172 17612
rect 25564 17668 25620 17678
rect 25564 17574 25620 17612
rect 26236 17108 26292 17726
rect 26236 17042 26292 17052
rect 25116 16046 25118 16098
rect 25170 16046 25172 16098
rect 25116 16034 25172 16046
rect 25788 16324 25844 16334
rect 25340 15540 25396 15550
rect 25340 15446 25396 15484
rect 25788 15538 25844 16268
rect 25900 16212 25956 16222
rect 25900 16118 25956 16156
rect 25788 15486 25790 15538
rect 25842 15486 25844 15538
rect 25788 15316 25844 15486
rect 25788 15250 25844 15260
rect 26348 15202 26404 15214
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 25900 15092 25956 15102
rect 25788 15036 25900 15092
rect 25564 14532 25620 14542
rect 25228 13860 25284 13870
rect 25228 13746 25284 13804
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25228 13682 25284 13694
rect 25564 13074 25620 14476
rect 25676 14420 25732 14430
rect 25676 13746 25732 14364
rect 25676 13694 25678 13746
rect 25730 13694 25732 13746
rect 25676 13682 25732 13694
rect 25564 13022 25566 13074
rect 25618 13022 25620 13074
rect 25564 13010 25620 13022
rect 25340 12740 25396 12750
rect 25340 12290 25396 12684
rect 25452 12404 25508 12414
rect 25788 12404 25844 15036
rect 25900 15026 25956 15036
rect 26348 14980 26404 15150
rect 26460 15148 26516 19292
rect 26460 15082 26516 15092
rect 26572 14980 26628 19404
rect 26012 14924 26628 14980
rect 25452 12310 25508 12348
rect 25564 12348 25844 12404
rect 25900 13522 25956 13534
rect 25900 13470 25902 13522
rect 25954 13470 25956 13522
rect 25340 12238 25342 12290
rect 25394 12238 25396 12290
rect 25340 12226 25396 12238
rect 25004 11844 25060 11854
rect 25004 11282 25060 11788
rect 25004 11230 25006 11282
rect 25058 11230 25060 11282
rect 25004 11218 25060 11230
rect 25116 11172 25172 11182
rect 24780 11004 24948 11060
rect 24556 10782 24558 10834
rect 24610 10782 24612 10834
rect 24556 10770 24612 10782
rect 24780 10836 24836 10846
rect 24780 10742 24836 10780
rect 24444 10670 24446 10722
rect 24498 10670 24500 10722
rect 24444 10658 24500 10670
rect 23660 10386 23716 10398
rect 23660 10334 23662 10386
rect 23714 10334 23716 10386
rect 23436 8372 23604 8428
rect 22428 8306 22484 8316
rect 23548 8370 23604 8372
rect 23548 8318 23550 8370
rect 23602 8318 23604 8370
rect 22316 8260 22372 8270
rect 22316 8166 22372 8204
rect 21868 7494 21924 7532
rect 22876 8036 22932 8046
rect 21644 7422 21646 7474
rect 21698 7422 21700 7474
rect 21644 7410 21700 7422
rect 21756 7362 21812 7374
rect 21756 7310 21758 7362
rect 21810 7310 21812 7362
rect 21532 5234 21588 5246
rect 21532 5182 21534 5234
rect 21586 5182 21588 5234
rect 21532 5124 21588 5182
rect 21532 5058 21588 5068
rect 21756 5122 21812 7310
rect 22316 5906 22372 5918
rect 22316 5854 22318 5906
rect 22370 5854 22372 5906
rect 22316 5684 22372 5854
rect 22876 5906 22932 7980
rect 23548 7476 23604 8318
rect 23660 8036 23716 10334
rect 23772 8260 23828 8270
rect 23828 8204 23940 8260
rect 23772 8166 23828 8204
rect 23660 7970 23716 7980
rect 23772 7476 23828 7486
rect 23548 7474 23828 7476
rect 23548 7422 23774 7474
rect 23826 7422 23828 7474
rect 23548 7420 23828 7422
rect 23772 6802 23828 7420
rect 23884 7364 23940 8204
rect 24108 8034 24164 8046
rect 24108 7982 24110 8034
rect 24162 7982 24164 8034
rect 24108 7476 24164 7982
rect 24108 7410 24164 7420
rect 23884 7362 24052 7364
rect 23884 7310 23886 7362
rect 23938 7310 24052 7362
rect 23884 7308 24052 7310
rect 23884 7298 23940 7308
rect 23996 6914 24052 7308
rect 24556 7250 24612 7262
rect 24556 7198 24558 7250
rect 24610 7198 24612 7250
rect 23996 6862 23998 6914
rect 24050 6862 24052 6914
rect 23996 6850 24052 6862
rect 24332 6916 24388 6926
rect 23772 6750 23774 6802
rect 23826 6750 23828 6802
rect 23772 6738 23828 6750
rect 24332 6690 24388 6860
rect 24332 6638 24334 6690
rect 24386 6638 24388 6690
rect 24332 6626 24388 6638
rect 22876 5854 22878 5906
rect 22930 5854 22932 5906
rect 22876 5842 22932 5854
rect 24556 5908 24612 7198
rect 24556 5842 24612 5852
rect 22988 5796 23044 5806
rect 22988 5794 23156 5796
rect 22988 5742 22990 5794
rect 23042 5742 23156 5794
rect 22988 5740 23156 5742
rect 22988 5730 23044 5740
rect 22316 5618 22372 5628
rect 23100 5234 23156 5740
rect 23100 5182 23102 5234
rect 23154 5182 23156 5234
rect 23100 5170 23156 5182
rect 24332 5236 24388 5246
rect 21756 5070 21758 5122
rect 21810 5070 21812 5122
rect 21756 5012 21812 5070
rect 22316 5124 22372 5134
rect 21756 4956 22148 5012
rect 22092 4450 22148 4956
rect 22092 4398 22094 4450
rect 22146 4398 22148 4450
rect 22092 4386 22148 4398
rect 22316 4338 22372 5068
rect 22428 5124 22484 5134
rect 22652 5124 22708 5134
rect 22428 5122 22652 5124
rect 22428 5070 22430 5122
rect 22482 5070 22652 5122
rect 22428 5068 22652 5070
rect 22428 5058 22484 5068
rect 22652 5058 22708 5068
rect 23324 5124 23380 5134
rect 23324 5122 23492 5124
rect 23324 5070 23326 5122
rect 23378 5070 23492 5122
rect 23324 5068 23492 5070
rect 23324 5058 23380 5068
rect 23436 4564 23492 5068
rect 24332 5122 24388 5180
rect 24332 5070 24334 5122
rect 24386 5070 24388 5122
rect 24332 5058 24388 5070
rect 23772 5012 23828 5022
rect 23660 4564 23716 4574
rect 23436 4562 23716 4564
rect 23436 4510 23662 4562
rect 23714 4510 23716 4562
rect 23436 4508 23716 4510
rect 23660 4498 23716 4508
rect 23772 4562 23828 4956
rect 23772 4510 23774 4562
rect 23826 4510 23828 4562
rect 23772 4498 23828 4510
rect 23100 4340 23156 4350
rect 22316 4286 22318 4338
rect 22370 4286 22372 4338
rect 22316 4274 22372 4286
rect 22652 4338 23156 4340
rect 22652 4286 23102 4338
rect 23154 4286 23156 4338
rect 22652 4284 23156 4286
rect 22652 4226 22708 4284
rect 23100 4274 23156 4284
rect 23548 4340 23604 4350
rect 23548 4246 23604 4284
rect 22652 4174 22654 4226
rect 22706 4174 22708 4226
rect 22652 4162 22708 4174
rect 22988 3668 23044 3678
rect 22988 3574 23044 3612
rect 24892 3668 24948 11004
rect 25004 9940 25060 9950
rect 25116 9940 25172 11116
rect 25004 9938 25172 9940
rect 25004 9886 25006 9938
rect 25058 9886 25172 9938
rect 25004 9884 25172 9886
rect 25564 9940 25620 12348
rect 25676 12178 25732 12190
rect 25676 12126 25678 12178
rect 25730 12126 25732 12178
rect 25676 11508 25732 12126
rect 25900 11620 25956 13470
rect 26012 13076 26068 14924
rect 26572 14420 26628 14430
rect 26684 14420 26740 19740
rect 26796 18452 26852 29036
rect 26908 28420 26964 35644
rect 27356 35588 27412 36428
rect 27244 35586 27412 35588
rect 27244 35534 27358 35586
rect 27410 35534 27412 35586
rect 27244 35532 27412 35534
rect 27132 35028 27188 35038
rect 27020 34914 27076 34926
rect 27020 34862 27022 34914
rect 27074 34862 27076 34914
rect 27020 34804 27076 34862
rect 27020 34738 27076 34748
rect 27020 34356 27076 34366
rect 27132 34356 27188 34972
rect 27020 34354 27188 34356
rect 27020 34302 27022 34354
rect 27074 34302 27188 34354
rect 27020 34300 27188 34302
rect 27020 31668 27076 34300
rect 27244 31892 27300 35532
rect 27356 35522 27412 35532
rect 27020 31602 27076 31612
rect 27132 31836 27300 31892
rect 27356 35364 27412 35374
rect 27020 30212 27076 30222
rect 27020 28754 27076 30156
rect 27020 28702 27022 28754
rect 27074 28702 27076 28754
rect 27020 28644 27076 28702
rect 27020 28578 27076 28588
rect 27020 28420 27076 28430
rect 26908 28364 27020 28420
rect 27020 28354 27076 28364
rect 27132 26964 27188 31836
rect 27244 31668 27300 31678
rect 27244 31218 27300 31612
rect 27244 31166 27246 31218
rect 27298 31166 27300 31218
rect 27244 31154 27300 31166
rect 27244 30212 27300 30222
rect 27244 30118 27300 30156
rect 27356 29988 27412 35308
rect 27468 33458 27524 33470
rect 27468 33406 27470 33458
rect 27522 33406 27524 33458
rect 27468 32340 27524 33406
rect 27468 32274 27524 32284
rect 27468 31668 27524 31678
rect 27468 31106 27524 31612
rect 27468 31054 27470 31106
rect 27522 31054 27524 31106
rect 27468 31042 27524 31054
rect 27580 30884 27636 43708
rect 27692 42756 27748 42766
rect 27692 42662 27748 42700
rect 27804 37604 27860 37614
rect 27692 37548 27804 37604
rect 27692 35028 27748 37548
rect 27804 37538 27860 37548
rect 27804 36594 27860 36606
rect 27804 36542 27806 36594
rect 27858 36542 27860 36594
rect 27804 36484 27860 36542
rect 27804 36418 27860 36428
rect 27804 35700 27860 35710
rect 27804 35606 27860 35644
rect 27916 35028 27972 50372
rect 28252 50260 28308 50270
rect 28028 49924 28084 49934
rect 28028 48804 28084 49868
rect 28028 48738 28084 48748
rect 28252 48242 28308 50204
rect 28364 49812 28420 50372
rect 28588 50372 28644 50382
rect 28588 50278 28644 50316
rect 28364 49746 28420 49756
rect 28588 49700 28644 49710
rect 28588 49606 28644 49644
rect 28252 48190 28254 48242
rect 28306 48190 28308 48242
rect 28252 48178 28308 48190
rect 28476 48466 28532 48478
rect 28476 48414 28478 48466
rect 28530 48414 28532 48466
rect 28252 47124 28308 47134
rect 28140 45332 28196 45342
rect 28028 42530 28084 42542
rect 28028 42478 28030 42530
rect 28082 42478 28084 42530
rect 28028 42420 28084 42478
rect 28028 42354 28084 42364
rect 28028 37268 28084 37278
rect 28028 37174 28084 37212
rect 28140 37266 28196 45276
rect 28252 37604 28308 47068
rect 28476 38668 28532 48414
rect 28588 48242 28644 48254
rect 28588 48190 28590 48242
rect 28642 48190 28644 48242
rect 28588 47124 28644 48190
rect 28588 47058 28644 47068
rect 28812 47012 28868 50876
rect 28924 50372 28980 51214
rect 29036 50484 29092 50522
rect 29036 50418 29092 50428
rect 28924 50306 28980 50316
rect 29148 49252 29204 53452
rect 29484 52836 29540 52846
rect 29260 52164 29316 52174
rect 29260 52070 29316 52108
rect 29372 51716 29428 51726
rect 29372 50594 29428 51660
rect 29372 50542 29374 50594
rect 29426 50542 29428 50594
rect 29372 50530 29428 50542
rect 29260 50482 29316 50494
rect 29260 50430 29262 50482
rect 29314 50430 29316 50482
rect 29260 50372 29316 50430
rect 29260 50306 29316 50316
rect 29148 49196 29316 49252
rect 29148 49028 29204 49038
rect 29148 48934 29204 48972
rect 28700 46956 28868 47012
rect 28700 45668 28756 46956
rect 29148 46788 29204 46798
rect 28252 37538 28308 37548
rect 28364 38612 28532 38668
rect 28588 45612 28756 45668
rect 28812 46732 29148 46788
rect 28364 37380 28420 38612
rect 28588 38276 28644 45612
rect 28700 45444 28756 45454
rect 28700 40628 28756 45388
rect 28700 40562 28756 40572
rect 28700 40404 28756 40414
rect 28700 40290 28756 40348
rect 28700 40238 28702 40290
rect 28754 40238 28756 40290
rect 28700 40226 28756 40238
rect 28700 40068 28756 40078
rect 28700 38500 28756 40012
rect 28700 38434 28756 38444
rect 28812 39058 28868 46732
rect 29148 46722 29204 46732
rect 29260 45668 29316 49196
rect 29260 45602 29316 45612
rect 29484 45444 29540 52780
rect 29596 46788 29652 57486
rect 29820 57484 29988 57540
rect 29708 56644 29764 56654
rect 29708 55748 29764 56588
rect 29708 55682 29764 55692
rect 29596 46722 29652 46732
rect 29708 52164 29764 52174
rect 29596 46564 29652 46574
rect 29596 46470 29652 46508
rect 29484 45378 29540 45388
rect 29596 45666 29652 45678
rect 29596 45614 29598 45666
rect 29650 45614 29652 45666
rect 29484 45108 29540 45118
rect 29260 45052 29484 45108
rect 29260 44994 29316 45052
rect 29484 45042 29540 45052
rect 29260 44942 29262 44994
rect 29314 44942 29316 44994
rect 29260 44930 29316 44942
rect 29596 44884 29652 45614
rect 29708 45556 29764 52108
rect 29820 51604 29876 57484
rect 30044 57428 30100 59052
rect 29932 57372 30100 57428
rect 30156 58434 30212 58446
rect 30156 58382 30158 58434
rect 30210 58382 30212 58434
rect 30156 57650 30212 58382
rect 30380 57764 30436 63756
rect 30492 63700 30548 63710
rect 30492 62356 30548 63644
rect 30604 62916 30660 65100
rect 31164 64482 31220 64494
rect 31164 64430 31166 64482
rect 31218 64430 31220 64482
rect 30940 63698 30996 63710
rect 30940 63646 30942 63698
rect 30994 63646 30996 63698
rect 30940 63364 30996 63646
rect 31164 63700 31220 64430
rect 31164 63634 31220 63644
rect 30940 63298 30996 63308
rect 31164 63026 31220 63038
rect 31164 62974 31166 63026
rect 31218 62974 31220 63026
rect 31052 62916 31108 62926
rect 30604 62914 31108 62916
rect 30604 62862 31054 62914
rect 31106 62862 31108 62914
rect 30604 62860 31108 62862
rect 31052 62850 31108 62860
rect 30492 62290 30548 62300
rect 31164 62244 31220 62974
rect 31164 62178 31220 62188
rect 31276 60788 31332 66220
rect 31836 65604 31892 66332
rect 32172 66388 32228 66398
rect 32172 66294 32228 66332
rect 32060 66276 32116 66286
rect 32060 66182 32116 66220
rect 32284 65828 32340 67172
rect 32508 67172 33236 67228
rect 32508 66386 32564 67172
rect 33180 67170 33236 67172
rect 33180 67118 33182 67170
rect 33234 67118 33236 67170
rect 33180 67106 33236 67118
rect 33404 67172 33684 67228
rect 34076 67732 34132 67742
rect 33404 67170 33460 67172
rect 33404 67118 33406 67170
rect 33458 67118 33460 67170
rect 33404 67106 33460 67118
rect 34076 67170 34132 67676
rect 34300 67228 34356 68684
rect 35644 68684 35812 68740
rect 36316 69300 36372 69310
rect 35196 68516 35252 68526
rect 35196 68422 35252 68460
rect 35084 68404 35140 68414
rect 34412 68402 35140 68404
rect 34412 68350 35086 68402
rect 35138 68350 35140 68402
rect 34412 68348 35140 68350
rect 34412 67842 34468 68348
rect 35084 68338 35140 68348
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 34412 67790 34414 67842
rect 34466 67790 34468 67842
rect 34412 67778 34468 67790
rect 35644 67508 35700 68684
rect 36316 68628 36372 69244
rect 36876 69300 36932 70140
rect 37660 70084 37716 70142
rect 37660 70018 37716 70028
rect 37772 70306 37828 70318
rect 37772 70254 37774 70306
rect 37826 70254 37828 70306
rect 37772 70196 37828 70254
rect 37100 69410 37156 69422
rect 37100 69358 37102 69410
rect 37154 69358 37156 69410
rect 37100 69300 37156 69358
rect 36876 69244 37156 69300
rect 37324 69410 37380 69422
rect 37324 69358 37326 69410
rect 37378 69358 37380 69410
rect 37324 69300 37380 69358
rect 36316 68572 36484 68628
rect 35756 68516 35812 68526
rect 35756 68422 35812 68460
rect 35756 67844 35812 67854
rect 35756 67842 36260 67844
rect 35756 67790 35758 67842
rect 35810 67790 36260 67842
rect 35756 67788 36260 67790
rect 35756 67778 35812 67788
rect 35644 67442 35700 67452
rect 34076 67118 34078 67170
rect 34130 67118 34132 67170
rect 34076 67106 34132 67118
rect 34188 67172 34356 67228
rect 36204 67282 36260 67788
rect 36204 67230 36206 67282
rect 36258 67230 36260 67282
rect 36204 67218 36260 67230
rect 33068 67060 33124 67070
rect 32508 66334 32510 66386
rect 32562 66334 32564 66386
rect 32508 66322 32564 66334
rect 32956 67058 33124 67060
rect 32956 67006 33070 67058
rect 33122 67006 33124 67058
rect 32956 67004 33124 67006
rect 32844 66276 32900 66286
rect 32844 66182 32900 66220
rect 31836 65538 31892 65548
rect 32172 65772 32340 65828
rect 31500 63810 31556 63822
rect 31500 63758 31502 63810
rect 31554 63758 31556 63810
rect 31500 63140 31556 63758
rect 31948 63812 32004 63822
rect 31948 63810 32116 63812
rect 31948 63758 31950 63810
rect 32002 63758 32116 63810
rect 31948 63756 32116 63758
rect 31948 63746 32004 63756
rect 31948 63364 32004 63374
rect 31948 63270 32004 63308
rect 31724 63140 31780 63150
rect 31500 63138 31780 63140
rect 31500 63086 31726 63138
rect 31778 63086 31780 63138
rect 31500 63084 31780 63086
rect 31388 62356 31444 62366
rect 31388 62262 31444 62300
rect 31724 62132 31780 63084
rect 31724 62066 31780 62076
rect 32060 62244 32116 63756
rect 32172 62468 32228 65772
rect 32396 65716 32452 65726
rect 32284 65602 32340 65614
rect 32284 65550 32286 65602
rect 32338 65550 32340 65602
rect 32284 65492 32340 65550
rect 32284 65426 32340 65436
rect 32396 65490 32452 65660
rect 32396 65438 32398 65490
rect 32450 65438 32452 65490
rect 32396 65426 32452 65438
rect 32508 65380 32564 65390
rect 32508 65266 32564 65324
rect 32508 65214 32510 65266
rect 32562 65214 32564 65266
rect 32284 63588 32340 63598
rect 32284 63362 32340 63532
rect 32284 63310 32286 63362
rect 32338 63310 32340 63362
rect 32284 63298 32340 63310
rect 32172 62412 32452 62468
rect 32172 62244 32228 62254
rect 32116 62242 32228 62244
rect 32116 62190 32174 62242
rect 32226 62190 32228 62242
rect 32116 62188 32228 62190
rect 31612 61684 31668 61694
rect 31500 61460 31556 61470
rect 31388 61012 31444 61022
rect 31388 60918 31444 60956
rect 31500 61010 31556 61404
rect 31612 61458 31668 61628
rect 31612 61406 31614 61458
rect 31666 61406 31668 61458
rect 31612 61394 31668 61406
rect 31948 61460 32004 61470
rect 32060 61460 32116 62188
rect 32172 62178 32228 62188
rect 31948 61458 32116 61460
rect 31948 61406 31950 61458
rect 32002 61406 32116 61458
rect 31948 61404 32116 61406
rect 31948 61394 32004 61404
rect 31500 60958 31502 61010
rect 31554 60958 31556 61010
rect 31500 60946 31556 60958
rect 31948 60900 32004 60910
rect 31164 60732 31332 60788
rect 31724 60844 31948 60900
rect 31052 59218 31108 59230
rect 31052 59166 31054 59218
rect 31106 59166 31108 59218
rect 30604 59108 30660 59118
rect 31052 59108 31108 59166
rect 30604 59106 31052 59108
rect 30604 59054 30606 59106
rect 30658 59054 31052 59106
rect 30604 59052 31052 59054
rect 30604 59042 30660 59052
rect 31052 59042 31108 59052
rect 30716 58436 30772 58446
rect 31164 58436 31220 60732
rect 31612 60564 31668 60574
rect 31612 60470 31668 60508
rect 31612 60228 31668 60238
rect 31724 60228 31780 60844
rect 31948 60806 32004 60844
rect 31836 60676 31892 60686
rect 31892 60620 32004 60676
rect 31836 60610 31892 60620
rect 31612 60226 31780 60228
rect 31612 60174 31614 60226
rect 31666 60174 31780 60226
rect 31612 60172 31780 60174
rect 31612 60162 31668 60172
rect 31724 59892 31780 59902
rect 31724 59798 31780 59836
rect 31276 59780 31332 59790
rect 31276 59686 31332 59724
rect 31612 59780 31668 59790
rect 31388 59668 31444 59678
rect 31276 59332 31332 59342
rect 31276 59238 31332 59276
rect 31388 58772 31444 59612
rect 31388 58716 31556 58772
rect 31388 58546 31444 58558
rect 31388 58494 31390 58546
rect 31442 58494 31444 58546
rect 30716 58434 31220 58436
rect 30716 58382 30718 58434
rect 30770 58382 31220 58434
rect 30716 58380 31220 58382
rect 31276 58434 31332 58446
rect 31276 58382 31278 58434
rect 31330 58382 31332 58434
rect 30716 58370 30772 58380
rect 31276 57764 31332 58382
rect 30380 57708 30884 57764
rect 30156 57598 30158 57650
rect 30210 57598 30212 57650
rect 30156 57428 30212 57598
rect 30156 57372 30324 57428
rect 29932 54740 29988 57372
rect 30268 57204 30324 57372
rect 30716 57426 30772 57438
rect 30716 57374 30718 57426
rect 30770 57374 30772 57426
rect 30492 57316 30548 57326
rect 30268 57138 30324 57148
rect 30380 57260 30492 57316
rect 30156 57092 30212 57102
rect 30044 56754 30100 56766
rect 30044 56702 30046 56754
rect 30098 56702 30100 56754
rect 30044 55972 30100 56702
rect 30156 56754 30212 57036
rect 30380 56866 30436 57260
rect 30492 57250 30548 57260
rect 30716 57204 30772 57374
rect 30716 57138 30772 57148
rect 30380 56814 30382 56866
rect 30434 56814 30436 56866
rect 30380 56802 30436 56814
rect 30156 56702 30158 56754
rect 30210 56702 30212 56754
rect 30156 56690 30212 56702
rect 30604 56754 30660 56766
rect 30604 56702 30606 56754
rect 30658 56702 30660 56754
rect 30156 55972 30212 55982
rect 30044 55970 30212 55972
rect 30044 55918 30158 55970
rect 30210 55918 30212 55970
rect 30044 55916 30212 55918
rect 29932 54684 30100 54740
rect 29932 53732 29988 53742
rect 29932 53638 29988 53676
rect 29820 50708 29876 51548
rect 29820 50614 29876 50652
rect 29932 48916 29988 48926
rect 29932 48822 29988 48860
rect 30044 48580 30100 54684
rect 30156 52836 30212 55916
rect 30604 55972 30660 56702
rect 30716 56642 30772 56654
rect 30716 56590 30718 56642
rect 30770 56590 30772 56642
rect 30716 56196 30772 56590
rect 30828 56308 30884 57708
rect 30940 57762 31332 57764
rect 30940 57710 31278 57762
rect 31330 57710 31332 57762
rect 30940 57708 31332 57710
rect 30940 56866 30996 57708
rect 31276 57698 31332 57708
rect 31052 57540 31108 57550
rect 31388 57540 31444 58494
rect 31052 57538 31444 57540
rect 31052 57486 31054 57538
rect 31106 57486 31444 57538
rect 31052 57484 31444 57486
rect 31052 57316 31108 57484
rect 31052 57250 31108 57260
rect 31276 57092 31332 57102
rect 31276 56978 31332 57036
rect 31276 56926 31278 56978
rect 31330 56926 31332 56978
rect 31276 56914 31332 56926
rect 30940 56814 30942 56866
rect 30994 56814 30996 56866
rect 30940 56802 30996 56814
rect 31500 56420 31556 58716
rect 31612 56644 31668 59724
rect 31612 56578 31668 56588
rect 31724 59108 31780 59118
rect 31724 56642 31780 59052
rect 31948 58658 32004 60620
rect 32060 59556 32116 61404
rect 32396 60788 32452 62412
rect 32508 61010 32564 65214
rect 32956 64148 33012 67004
rect 33068 66994 33124 67004
rect 34188 66386 34244 67172
rect 36316 67170 36372 67182
rect 36316 67118 36318 67170
rect 36370 67118 36372 67170
rect 35308 67060 35364 67070
rect 35308 66836 35364 67004
rect 35644 67060 35700 67070
rect 36092 67060 36148 67070
rect 35644 67058 36148 67060
rect 35644 67006 35646 67058
rect 35698 67006 36094 67058
rect 36146 67006 36148 67058
rect 35644 67004 36148 67006
rect 35308 66780 35588 66836
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 34188 66334 34190 66386
rect 34242 66334 34244 66386
rect 34188 66322 34244 66334
rect 34300 66388 34356 66398
rect 33404 66276 33460 66286
rect 33404 66182 33460 66220
rect 33740 66274 33796 66286
rect 33740 66222 33742 66274
rect 33794 66222 33796 66274
rect 33740 65716 33796 66222
rect 34300 66274 34356 66332
rect 34300 66222 34302 66274
rect 34354 66222 34356 66274
rect 34300 65940 34356 66222
rect 34412 66276 34468 66286
rect 34412 66162 34468 66220
rect 34412 66110 34414 66162
rect 34466 66110 34468 66162
rect 34412 66098 34468 66110
rect 33740 65650 33796 65660
rect 34076 65884 34356 65940
rect 34076 65602 34132 65884
rect 34076 65550 34078 65602
rect 34130 65550 34132 65602
rect 34076 65538 34132 65550
rect 34524 65604 34580 65614
rect 33628 65492 33684 65502
rect 33180 65380 33236 65390
rect 33180 65286 33236 65324
rect 33628 64708 33684 65436
rect 34412 64820 34468 64830
rect 33740 64708 33796 64718
rect 33628 64706 33796 64708
rect 33628 64654 33742 64706
rect 33794 64654 33796 64706
rect 33628 64652 33796 64654
rect 33740 64642 33796 64652
rect 32732 64092 33012 64148
rect 32732 61682 32788 64092
rect 34412 63362 34468 64764
rect 34412 63310 34414 63362
rect 34466 63310 34468 63362
rect 34412 63298 34468 63310
rect 34300 63250 34356 63262
rect 34300 63198 34302 63250
rect 34354 63198 34356 63250
rect 34188 63138 34244 63150
rect 34188 63086 34190 63138
rect 34242 63086 34244 63138
rect 34188 63028 34244 63086
rect 34188 62962 34244 62972
rect 34300 63140 34356 63198
rect 34524 63140 34580 65548
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35532 64932 35588 66780
rect 35644 66498 35700 67004
rect 36092 66994 36148 67004
rect 36316 67060 36372 67118
rect 36316 66994 36372 67004
rect 35644 66446 35646 66498
rect 35698 66446 35700 66498
rect 35644 66434 35700 66446
rect 36092 66386 36148 66398
rect 36092 66334 36094 66386
rect 36146 66334 36148 66386
rect 35868 66274 35924 66286
rect 35868 66222 35870 66274
rect 35922 66222 35924 66274
rect 35868 65602 35924 66222
rect 35868 65550 35870 65602
rect 35922 65550 35924 65602
rect 35756 64932 35812 64942
rect 35532 64930 35812 64932
rect 35532 64878 35758 64930
rect 35810 64878 35812 64930
rect 35532 64876 35812 64878
rect 35756 64866 35812 64876
rect 35420 64820 35476 64830
rect 35420 64726 35476 64764
rect 34636 64706 34692 64718
rect 34636 64654 34638 64706
rect 34690 64654 34692 64706
rect 34636 64596 34692 64654
rect 35196 64596 35252 64606
rect 34636 64594 35252 64596
rect 34636 64542 35198 64594
rect 35250 64542 35252 64594
rect 34636 64540 35252 64542
rect 33180 62356 33236 62366
rect 33180 62262 33236 62300
rect 32732 61630 32734 61682
rect 32786 61630 32788 61682
rect 32732 61618 32788 61630
rect 32844 61570 32900 61582
rect 32844 61518 32846 61570
rect 32898 61518 32900 61570
rect 32620 61460 32676 61470
rect 32620 61366 32676 61404
rect 32508 60958 32510 61010
rect 32562 60958 32564 61010
rect 32508 60946 32564 60958
rect 32620 60788 32676 60798
rect 32396 60732 32620 60788
rect 32172 60676 32228 60686
rect 32172 60582 32228 60620
rect 32508 60564 32564 60574
rect 32508 60114 32564 60508
rect 32508 60062 32510 60114
rect 32562 60062 32564 60114
rect 32508 60050 32564 60062
rect 32172 59892 32228 59902
rect 32172 59798 32228 59836
rect 32396 59780 32452 59790
rect 32396 59686 32452 59724
rect 32620 59778 32676 60732
rect 32844 60114 32900 61518
rect 33180 61460 33236 61470
rect 33740 61460 33796 61470
rect 33180 61458 33348 61460
rect 33180 61406 33182 61458
rect 33234 61406 33348 61458
rect 33180 61404 33348 61406
rect 33180 61394 33236 61404
rect 33180 61012 33236 61022
rect 33292 61012 33348 61404
rect 33740 61458 33908 61460
rect 33740 61406 33742 61458
rect 33794 61406 33908 61458
rect 33740 61404 33908 61406
rect 33740 61394 33796 61404
rect 33404 61348 33460 61358
rect 33404 61346 33572 61348
rect 33404 61294 33406 61346
rect 33458 61294 33572 61346
rect 33404 61292 33572 61294
rect 33404 61282 33460 61292
rect 33404 61012 33460 61022
rect 33292 61010 33460 61012
rect 33292 60958 33406 61010
rect 33458 60958 33460 61010
rect 33292 60956 33460 60958
rect 32956 60786 33012 60798
rect 32956 60734 32958 60786
rect 33010 60734 33012 60786
rect 32956 60564 33012 60734
rect 33180 60788 33236 60956
rect 33404 60946 33460 60956
rect 33292 60788 33348 60798
rect 33180 60786 33348 60788
rect 33180 60734 33294 60786
rect 33346 60734 33348 60786
rect 33180 60732 33348 60734
rect 33292 60722 33348 60732
rect 33516 60786 33572 61292
rect 33628 61346 33684 61358
rect 33628 61294 33630 61346
rect 33682 61294 33684 61346
rect 33628 60900 33684 61294
rect 33628 60834 33684 60844
rect 33516 60734 33518 60786
rect 33570 60734 33572 60786
rect 32956 60498 33012 60508
rect 33404 60564 33460 60574
rect 32844 60062 32846 60114
rect 32898 60062 32900 60114
rect 32844 60050 32900 60062
rect 33180 60340 33236 60350
rect 33180 60002 33236 60284
rect 33180 59950 33182 60002
rect 33234 59950 33236 60002
rect 33180 59938 33236 59950
rect 33404 60002 33460 60508
rect 33404 59950 33406 60002
rect 33458 59950 33460 60002
rect 32620 59726 32622 59778
rect 32674 59726 32676 59778
rect 32060 59500 32452 59556
rect 31948 58606 31950 58658
rect 32002 58606 32004 58658
rect 31948 58594 32004 58606
rect 32172 59108 32228 59118
rect 31724 56590 31726 56642
rect 31778 56590 31780 56642
rect 31276 56364 31556 56420
rect 30828 56252 31220 56308
rect 30716 56130 30772 56140
rect 30604 55878 30660 55916
rect 30604 55748 30660 55758
rect 30156 52770 30212 52780
rect 30268 52834 30324 52846
rect 30268 52782 30270 52834
rect 30322 52782 30324 52834
rect 30268 52388 30324 52782
rect 30268 52322 30324 52332
rect 30268 51268 30324 51278
rect 30268 51174 30324 51212
rect 30268 50596 30324 50606
rect 30268 50502 30324 50540
rect 30044 48514 30100 48524
rect 30380 50260 30436 50270
rect 30268 47348 30324 47358
rect 30268 45778 30324 47292
rect 30268 45726 30270 45778
rect 30322 45726 30324 45778
rect 30268 45714 30324 45726
rect 29708 45490 29764 45500
rect 29932 45666 29988 45678
rect 29932 45614 29934 45666
rect 29986 45614 29988 45666
rect 29932 45330 29988 45614
rect 29932 45278 29934 45330
rect 29986 45278 29988 45330
rect 29820 45106 29876 45118
rect 29820 45054 29822 45106
rect 29874 45054 29876 45106
rect 29708 44884 29764 44894
rect 29820 44884 29876 45054
rect 29932 45108 29988 45278
rect 30268 45444 30324 45454
rect 29932 45042 29988 45052
rect 30044 45220 30100 45230
rect 29596 44828 29708 44884
rect 29764 44828 29876 44884
rect 29708 44818 29764 44828
rect 29708 44548 29764 44558
rect 29708 44210 29764 44492
rect 30044 44322 30100 45164
rect 30156 45108 30212 45118
rect 30156 45014 30212 45052
rect 30268 44884 30324 45388
rect 30044 44270 30046 44322
rect 30098 44270 30100 44322
rect 30044 44258 30100 44270
rect 30156 44828 30324 44884
rect 29708 44158 29710 44210
rect 29762 44158 29764 44210
rect 29372 44100 29428 44110
rect 29708 44100 29764 44158
rect 29372 44098 29764 44100
rect 29372 44046 29374 44098
rect 29426 44046 29764 44098
rect 29372 44044 29764 44046
rect 29372 44034 29428 44044
rect 29708 43652 29764 44044
rect 29708 43586 29764 43596
rect 29820 44098 29876 44110
rect 29820 44046 29822 44098
rect 29874 44046 29876 44098
rect 29820 43988 29876 44046
rect 30156 43988 30212 44828
rect 29820 43932 30212 43988
rect 29372 43428 29428 43438
rect 29820 43428 29876 43932
rect 29372 43426 29876 43428
rect 29372 43374 29374 43426
rect 29426 43374 29876 43426
rect 29372 43372 29876 43374
rect 29372 43362 29428 43372
rect 29820 41972 29876 41982
rect 29596 41860 29652 41870
rect 29596 41766 29652 41804
rect 28812 39006 28814 39058
rect 28866 39006 28868 39058
rect 28588 38210 28644 38220
rect 28476 38164 28532 38174
rect 28476 38070 28532 38108
rect 28812 38052 28868 39006
rect 29596 38948 29652 38958
rect 29596 38854 29652 38892
rect 29820 38946 29876 41916
rect 30380 41186 30436 50204
rect 30604 48916 30660 55692
rect 31052 52946 31108 52958
rect 31052 52894 31054 52946
rect 31106 52894 31108 52946
rect 30716 52836 30772 52846
rect 31052 52836 31108 52894
rect 30772 52780 31108 52836
rect 30716 52742 30772 52780
rect 30716 51380 30772 51390
rect 30716 51378 31108 51380
rect 30716 51326 30718 51378
rect 30770 51326 31108 51378
rect 30716 51324 31108 51326
rect 30716 51314 30772 51324
rect 31052 50482 31108 51324
rect 31052 50430 31054 50482
rect 31106 50430 31108 50482
rect 31052 50372 31108 50430
rect 30604 48850 30660 48860
rect 30716 49698 30772 49710
rect 30716 49646 30718 49698
rect 30770 49646 30772 49698
rect 30716 48804 30772 49646
rect 30716 48738 30772 48748
rect 30716 47348 30772 47358
rect 30716 46786 30772 47292
rect 30716 46734 30718 46786
rect 30770 46734 30772 46786
rect 30716 46722 30772 46734
rect 30604 46450 30660 46462
rect 30604 46398 30606 46450
rect 30658 46398 30660 46450
rect 30604 46340 30660 46398
rect 30492 46284 30660 46340
rect 30492 45332 30548 46284
rect 31052 46116 31108 50316
rect 30492 45266 30548 45276
rect 30604 46060 31108 46116
rect 30380 41134 30382 41186
rect 30434 41134 30436 41186
rect 30380 41122 30436 41134
rect 30156 40962 30212 40974
rect 30156 40910 30158 40962
rect 30210 40910 30212 40962
rect 30156 40740 30212 40910
rect 30156 40674 30212 40684
rect 30492 40962 30548 40974
rect 30492 40910 30494 40962
rect 30546 40910 30548 40962
rect 30380 40402 30436 40414
rect 30380 40350 30382 40402
rect 30434 40350 30436 40402
rect 30380 40292 30436 40350
rect 30380 40068 30436 40236
rect 30380 40002 30436 40012
rect 30492 39844 30548 40910
rect 30604 40962 30660 46060
rect 30828 45780 30884 45790
rect 30828 45686 30884 45724
rect 31052 45778 31108 45790
rect 31052 45726 31054 45778
rect 31106 45726 31108 45778
rect 30940 45666 30996 45678
rect 30940 45614 30942 45666
rect 30994 45614 30996 45666
rect 30828 45220 30884 45230
rect 30716 45108 30772 45118
rect 30716 44994 30772 45052
rect 30828 45106 30884 45164
rect 30828 45054 30830 45106
rect 30882 45054 30884 45106
rect 30828 45042 30884 45054
rect 30716 44942 30718 44994
rect 30770 44942 30772 44994
rect 30716 44930 30772 44942
rect 30716 44324 30772 44334
rect 30716 44230 30772 44268
rect 30940 44322 30996 45614
rect 31052 44884 31108 45726
rect 31164 45556 31220 56252
rect 31276 48468 31332 56364
rect 31724 56308 31780 56590
rect 31500 56252 31780 56308
rect 31500 56196 31556 56252
rect 31388 54402 31444 54414
rect 31388 54350 31390 54402
rect 31442 54350 31444 54402
rect 31388 53284 31444 54350
rect 31388 53218 31444 53228
rect 31388 53058 31444 53070
rect 31388 53006 31390 53058
rect 31442 53006 31444 53058
rect 31388 52836 31444 53006
rect 31388 52770 31444 52780
rect 31500 51156 31556 56140
rect 31612 56084 31668 56094
rect 31612 53620 31668 56028
rect 32172 55412 32228 59052
rect 32172 55346 32228 55356
rect 32060 54404 32116 54414
rect 32060 53842 32116 54348
rect 32284 54402 32340 54414
rect 32284 54350 32286 54402
rect 32338 54350 32340 54402
rect 32284 54290 32340 54350
rect 32284 54238 32286 54290
rect 32338 54238 32340 54290
rect 32284 54226 32340 54238
rect 32060 53790 32062 53842
rect 32114 53790 32116 53842
rect 32060 53778 32116 53790
rect 31612 53554 31668 53564
rect 31836 53508 31892 53518
rect 31724 53452 31836 53508
rect 31724 52164 31780 53452
rect 31836 53442 31892 53452
rect 31724 52070 31780 52108
rect 31836 53116 32340 53172
rect 31500 51090 31556 51100
rect 31612 52052 31668 52062
rect 31388 50372 31444 50382
rect 31388 50370 31556 50372
rect 31388 50318 31390 50370
rect 31442 50318 31556 50370
rect 31388 50316 31556 50318
rect 31388 50306 31444 50316
rect 31388 49698 31444 49710
rect 31388 49646 31390 49698
rect 31442 49646 31444 49698
rect 31388 49140 31444 49646
rect 31500 49700 31556 50316
rect 31612 49810 31668 51996
rect 31836 51716 31892 53116
rect 32284 53058 32340 53116
rect 32284 53006 32286 53058
rect 32338 53006 32340 53058
rect 32284 52994 32340 53006
rect 32172 52946 32228 52958
rect 32172 52894 32174 52946
rect 32226 52894 32228 52946
rect 32172 52836 32228 52894
rect 32172 52770 32228 52780
rect 32284 52276 32340 52286
rect 32284 52182 32340 52220
rect 31724 51660 31892 51716
rect 32172 52164 32228 52174
rect 31724 50372 31780 51660
rect 32172 50428 32228 52108
rect 32396 51380 32452 59500
rect 32620 59332 32676 59726
rect 32620 59266 32676 59276
rect 32956 59890 33012 59902
rect 32956 59838 32958 59890
rect 33010 59838 33012 59890
rect 32956 59108 33012 59838
rect 32956 59042 33012 59052
rect 33180 59780 33236 59790
rect 33180 59218 33236 59724
rect 33180 59166 33182 59218
rect 33234 59166 33236 59218
rect 32844 56644 32900 56654
rect 33068 56644 33124 56654
rect 32844 56642 33124 56644
rect 32844 56590 32846 56642
rect 32898 56590 33070 56642
rect 33122 56590 33124 56642
rect 32844 56588 33124 56590
rect 32844 55972 32900 56588
rect 33068 56578 33124 56588
rect 33180 56308 33236 59166
rect 33404 58828 33460 59950
rect 33516 60004 33572 60734
rect 33740 60674 33796 60686
rect 33740 60622 33742 60674
rect 33794 60622 33796 60674
rect 33740 60340 33796 60622
rect 33740 60274 33796 60284
rect 33852 60676 33908 61404
rect 34188 61346 34244 61358
rect 34188 61294 34190 61346
rect 34242 61294 34244 61346
rect 33628 60004 33684 60014
rect 33516 60002 33684 60004
rect 33516 59950 33630 60002
rect 33682 59950 33684 60002
rect 33516 59948 33684 59950
rect 33628 59938 33684 59948
rect 33852 60002 33908 60620
rect 33852 59950 33854 60002
rect 33906 59950 33908 60002
rect 33852 59938 33908 59950
rect 33964 60788 34020 60798
rect 34188 60788 34244 61294
rect 33964 60786 34244 60788
rect 33964 60734 33966 60786
rect 34018 60734 34244 60786
rect 33964 60732 34244 60734
rect 33516 59108 33572 59118
rect 33516 59014 33572 59052
rect 33964 59108 34020 60732
rect 34188 60562 34244 60574
rect 34188 60510 34190 60562
rect 34242 60510 34244 60562
rect 34188 59890 34244 60510
rect 34188 59838 34190 59890
rect 34242 59838 34244 59890
rect 34076 59780 34132 59790
rect 34076 59686 34132 59724
rect 34076 59218 34132 59230
rect 34076 59166 34078 59218
rect 34130 59166 34132 59218
rect 34076 59108 34132 59166
rect 34020 59052 34132 59108
rect 34188 59108 34244 59838
rect 33964 59042 34020 59052
rect 34188 59042 34244 59052
rect 33404 58772 33796 58828
rect 33740 57874 33796 58772
rect 33740 57822 33742 57874
rect 33794 57822 33796 57874
rect 33740 57810 33796 57822
rect 33964 57762 34020 57774
rect 33964 57710 33966 57762
rect 34018 57710 34020 57762
rect 33516 57652 33572 57662
rect 33516 57540 33572 57596
rect 33404 57538 33572 57540
rect 33404 57486 33518 57538
rect 33570 57486 33572 57538
rect 33404 57484 33572 57486
rect 33404 56644 33460 57484
rect 33516 57474 33572 57484
rect 32508 55300 32564 55310
rect 32508 53170 32564 55244
rect 32508 53118 32510 53170
rect 32562 53118 32564 53170
rect 32508 53106 32564 53118
rect 32620 54292 32676 54302
rect 32844 54292 32900 55916
rect 32620 54290 32900 54292
rect 32620 54238 32622 54290
rect 32674 54238 32900 54290
rect 32620 54236 32900 54238
rect 33068 56252 33236 56308
rect 33292 56642 33460 56644
rect 33292 56590 33406 56642
rect 33458 56590 33460 56642
rect 33292 56588 33460 56590
rect 32620 53506 32676 54236
rect 33068 54180 33124 56252
rect 33292 56196 33348 56588
rect 33404 56578 33460 56588
rect 32620 53454 32622 53506
rect 32674 53454 32676 53506
rect 32620 52724 32676 53454
rect 32508 52668 32676 52724
rect 32732 54124 33124 54180
rect 33180 56140 33348 56196
rect 33516 56194 33572 56206
rect 33516 56142 33518 56194
rect 33570 56142 33572 56194
rect 32508 51716 32564 52668
rect 32732 52612 32788 54124
rect 32956 53844 33012 53854
rect 32956 53618 33012 53788
rect 32956 53566 32958 53618
rect 33010 53566 33012 53618
rect 32956 53554 33012 53566
rect 33180 53396 33236 56140
rect 33292 55970 33348 55982
rect 33292 55918 33294 55970
rect 33346 55918 33348 55970
rect 33292 55298 33348 55918
rect 33516 55468 33572 56142
rect 33516 55412 33796 55468
rect 33292 55246 33294 55298
rect 33346 55246 33348 55298
rect 33292 55188 33348 55246
rect 33516 55300 33572 55310
rect 33516 55206 33572 55244
rect 33292 53956 33348 55132
rect 33516 54964 33572 54974
rect 33516 54738 33572 54908
rect 33516 54686 33518 54738
rect 33570 54686 33572 54738
rect 33516 54674 33572 54686
rect 33740 54852 33796 55412
rect 33740 54738 33796 54796
rect 33740 54686 33742 54738
rect 33794 54686 33796 54738
rect 33740 54674 33796 54686
rect 33852 55074 33908 55086
rect 33852 55022 33854 55074
rect 33906 55022 33908 55074
rect 33852 54740 33908 55022
rect 33964 54964 34020 57710
rect 34076 57652 34132 57662
rect 34076 57558 34132 57596
rect 34188 55188 34244 55198
rect 34188 55094 34244 55132
rect 33964 54898 34020 54908
rect 34076 55076 34132 55086
rect 33964 54740 34020 54750
rect 33852 54738 34020 54740
rect 33852 54686 33966 54738
rect 34018 54686 34020 54738
rect 33852 54684 34020 54686
rect 33964 54674 34020 54684
rect 34076 54738 34132 55020
rect 34076 54686 34078 54738
rect 34130 54686 34132 54738
rect 34076 54674 34132 54686
rect 34188 54852 34244 54862
rect 34188 54738 34244 54796
rect 34188 54686 34190 54738
rect 34242 54686 34244 54738
rect 34188 54674 34244 54686
rect 33404 54514 33460 54526
rect 33404 54462 33406 54514
rect 33458 54462 33460 54514
rect 33404 54180 33460 54462
rect 33404 54124 33908 54180
rect 33404 53956 33460 53966
rect 33292 53954 33460 53956
rect 33292 53902 33406 53954
rect 33458 53902 33460 53954
rect 33292 53900 33460 53902
rect 33404 53890 33460 53900
rect 33516 53844 33572 53854
rect 33516 53730 33572 53788
rect 33516 53678 33518 53730
rect 33570 53678 33572 53730
rect 33516 53666 33572 53678
rect 33404 53508 33460 53518
rect 33404 53414 33460 53452
rect 33852 53396 33908 54124
rect 33964 53506 34020 53518
rect 33964 53454 33966 53506
rect 34018 53454 34020 53506
rect 33964 53396 34020 53454
rect 32620 52556 32788 52612
rect 32956 53340 33236 53396
rect 33516 53340 34020 53396
rect 32620 52052 32676 52556
rect 32844 52164 32900 52174
rect 32620 51958 32676 51996
rect 32732 52162 32900 52164
rect 32732 52110 32846 52162
rect 32898 52110 32900 52162
rect 32732 52108 32900 52110
rect 32732 51940 32788 52108
rect 32844 52098 32900 52108
rect 32508 51660 32676 51716
rect 32508 51380 32564 51390
rect 32396 51324 32508 51380
rect 32508 51314 32564 51324
rect 32508 50594 32564 50606
rect 32508 50542 32510 50594
rect 32562 50542 32564 50594
rect 32172 50372 32340 50428
rect 31724 50306 31780 50316
rect 31612 49758 31614 49810
rect 31666 49758 31668 49810
rect 31612 49746 31668 49758
rect 31500 49634 31556 49644
rect 31388 49074 31444 49084
rect 31948 49586 32004 49598
rect 31948 49534 31950 49586
rect 32002 49534 32004 49586
rect 31724 48916 31780 48926
rect 31276 48412 31668 48468
rect 31500 48242 31556 48254
rect 31500 48190 31502 48242
rect 31554 48190 31556 48242
rect 31276 46562 31332 46574
rect 31276 46510 31278 46562
rect 31330 46510 31332 46562
rect 31276 45892 31332 46510
rect 31500 46564 31556 48190
rect 31388 45892 31444 45902
rect 31276 45890 31444 45892
rect 31276 45838 31390 45890
rect 31442 45838 31444 45890
rect 31276 45836 31444 45838
rect 31164 45490 31220 45500
rect 31388 45332 31444 45836
rect 31500 45778 31556 46508
rect 31500 45726 31502 45778
rect 31554 45726 31556 45778
rect 31500 45714 31556 45726
rect 31388 45266 31444 45276
rect 31052 44882 31556 44884
rect 31052 44830 31054 44882
rect 31106 44830 31556 44882
rect 31052 44828 31556 44830
rect 31052 44818 31108 44828
rect 31500 44434 31556 44828
rect 31500 44382 31502 44434
rect 31554 44382 31556 44434
rect 31500 44370 31556 44382
rect 30940 44270 30942 44322
rect 30994 44270 30996 44322
rect 30940 44258 30996 44270
rect 31052 44212 31108 44222
rect 31612 44212 31668 48412
rect 31052 44210 31220 44212
rect 31052 44158 31054 44210
rect 31106 44158 31220 44210
rect 31052 44156 31220 44158
rect 31052 44146 31108 44156
rect 31052 41858 31108 41870
rect 31052 41806 31054 41858
rect 31106 41806 31108 41858
rect 30604 40910 30606 40962
rect 30658 40910 30660 40962
rect 30604 40068 30660 40910
rect 30940 41186 30996 41198
rect 30940 41134 30942 41186
rect 30994 41134 30996 41186
rect 30940 40740 30996 41134
rect 31052 41076 31108 41806
rect 31052 41010 31108 41020
rect 31164 40852 31220 44156
rect 30940 40674 30996 40684
rect 31052 40796 31220 40852
rect 31276 44156 31668 44212
rect 31724 47572 31780 48860
rect 31836 48692 31892 48702
rect 31836 48466 31892 48636
rect 31836 48414 31838 48466
rect 31890 48414 31892 48466
rect 31836 48402 31892 48414
rect 30828 40404 30884 40414
rect 30828 40310 30884 40348
rect 30604 40012 30884 40068
rect 29820 38894 29822 38946
rect 29874 38894 29876 38946
rect 29372 38834 29428 38846
rect 29372 38782 29374 38834
rect 29426 38782 29428 38834
rect 29036 38388 29092 38398
rect 28812 37986 28868 37996
rect 28924 38276 28980 38286
rect 28140 37214 28142 37266
rect 28194 37214 28196 37266
rect 28140 37044 28196 37214
rect 28028 36988 28196 37044
rect 28252 37324 28420 37380
rect 28028 36482 28084 36988
rect 28028 36430 28030 36482
rect 28082 36430 28084 36482
rect 28028 36418 28084 36430
rect 28252 35812 28308 37324
rect 28588 37268 28644 37278
rect 28364 37156 28420 37166
rect 28364 36706 28420 37100
rect 28588 37154 28644 37212
rect 28588 37102 28590 37154
rect 28642 37102 28644 37154
rect 28588 37090 28644 37102
rect 28364 36654 28366 36706
rect 28418 36654 28420 36706
rect 28364 36642 28420 36654
rect 28476 37042 28532 37054
rect 28476 36990 28478 37042
rect 28530 36990 28532 37042
rect 28140 35756 28308 35812
rect 28476 35812 28532 36990
rect 27748 34972 27860 35028
rect 27916 34972 28084 35028
rect 27692 34962 27748 34972
rect 27804 34804 27860 34972
rect 27916 34804 27972 34814
rect 27804 34802 27972 34804
rect 27804 34750 27918 34802
rect 27970 34750 27972 34802
rect 27804 34748 27972 34750
rect 27916 34738 27972 34748
rect 27916 34580 27972 34590
rect 27916 34130 27972 34524
rect 27916 34078 27918 34130
rect 27970 34078 27972 34130
rect 27916 34066 27972 34078
rect 26908 26908 27188 26964
rect 27244 29932 27412 29988
rect 27468 30828 27636 30884
rect 27244 26908 27300 29932
rect 27356 29540 27412 29550
rect 27356 29446 27412 29484
rect 27468 28980 27524 30828
rect 28028 30436 28084 34972
rect 27580 30380 28084 30436
rect 27580 30210 27636 30380
rect 28140 30324 28196 35756
rect 28476 35746 28532 35756
rect 28700 36372 28756 36382
rect 28252 35586 28308 35598
rect 28252 35534 28254 35586
rect 28306 35534 28308 35586
rect 28252 35364 28308 35534
rect 28252 35298 28308 35308
rect 28700 35586 28756 36316
rect 28700 35534 28702 35586
rect 28754 35534 28756 35586
rect 28476 35026 28532 35038
rect 28476 34974 28478 35026
rect 28530 34974 28532 35026
rect 28364 34804 28420 34814
rect 28252 34748 28364 34804
rect 28252 34018 28308 34748
rect 28364 34738 28420 34748
rect 28476 34580 28532 34974
rect 28476 34514 28532 34524
rect 28588 34020 28644 34030
rect 28252 33966 28254 34018
rect 28306 33966 28308 34018
rect 28252 33954 28308 33966
rect 28364 34018 28644 34020
rect 28364 33966 28590 34018
rect 28642 33966 28644 34018
rect 28364 33964 28644 33966
rect 28252 32788 28308 32798
rect 28252 32694 28308 32732
rect 27580 30158 27582 30210
rect 27634 30158 27636 30210
rect 27580 30146 27636 30158
rect 27804 30268 28196 30324
rect 27356 28924 27524 28980
rect 27356 27748 27412 28924
rect 27580 28868 27636 28906
rect 27580 28802 27636 28812
rect 27468 28754 27524 28766
rect 27468 28702 27470 28754
rect 27522 28702 27524 28754
rect 27468 27972 27524 28702
rect 27580 28644 27636 28654
rect 27580 28550 27636 28588
rect 27580 27972 27636 27982
rect 27468 27970 27636 27972
rect 27468 27918 27582 27970
rect 27634 27918 27636 27970
rect 27468 27916 27636 27918
rect 27580 27906 27636 27916
rect 27356 27692 27636 27748
rect 26908 22148 26964 26908
rect 27244 26852 27412 26908
rect 26908 22082 26964 22092
rect 27020 26740 27076 26750
rect 27020 21924 27076 26684
rect 27132 26178 27188 26190
rect 27132 26126 27134 26178
rect 27186 26126 27188 26178
rect 27132 25508 27188 26126
rect 27132 25442 27188 25452
rect 27132 24836 27188 24846
rect 27132 24742 27188 24780
rect 27356 23380 27412 26852
rect 27468 26068 27524 26078
rect 27468 25974 27524 26012
rect 27580 25844 27636 27692
rect 27692 26852 27748 26862
rect 27692 26758 27748 26796
rect 27468 25788 27636 25844
rect 27692 26290 27748 26302
rect 27692 26238 27694 26290
rect 27746 26238 27748 26290
rect 27468 25508 27524 25788
rect 27468 25442 27524 25452
rect 27580 25620 27636 25630
rect 27692 25620 27748 26238
rect 27580 25618 27748 25620
rect 27580 25566 27582 25618
rect 27634 25566 27748 25618
rect 27580 25564 27748 25566
rect 27580 24948 27636 25564
rect 26908 21868 27076 21924
rect 27132 23324 27412 23380
rect 27468 24892 27636 24948
rect 27692 24948 27748 24958
rect 26908 21140 26964 21868
rect 26908 21074 26964 21084
rect 27020 21474 27076 21486
rect 27020 21422 27022 21474
rect 27074 21422 27076 21474
rect 27020 21028 27076 21422
rect 27020 20934 27076 20972
rect 26796 18386 26852 18396
rect 26628 14364 26740 14420
rect 26908 14420 26964 14430
rect 26572 14326 26628 14364
rect 26908 14326 26964 14364
rect 27132 13972 27188 23324
rect 27244 23156 27300 23166
rect 27468 23156 27524 24892
rect 27580 24722 27636 24734
rect 27580 24670 27582 24722
rect 27634 24670 27636 24722
rect 27580 23380 27636 24670
rect 27580 23314 27636 23324
rect 27244 23154 27524 23156
rect 27244 23102 27246 23154
rect 27298 23102 27524 23154
rect 27244 23100 27524 23102
rect 27580 23156 27636 23166
rect 27244 23090 27300 23100
rect 27580 23062 27636 23100
rect 27244 22372 27300 22382
rect 27244 22278 27300 22316
rect 27244 22148 27300 22158
rect 27580 22148 27636 22158
rect 27244 21364 27300 22092
rect 27356 22146 27636 22148
rect 27356 22094 27582 22146
rect 27634 22094 27636 22146
rect 27356 22092 27636 22094
rect 27356 21586 27412 22092
rect 27580 22082 27636 22092
rect 27356 21534 27358 21586
rect 27410 21534 27412 21586
rect 27356 21522 27412 21534
rect 27244 21308 27524 21364
rect 27244 21140 27300 21150
rect 27244 20802 27300 21084
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 27244 20738 27300 20750
rect 27356 20914 27412 20926
rect 27356 20862 27358 20914
rect 27410 20862 27412 20914
rect 27356 20692 27412 20862
rect 27356 20626 27412 20636
rect 27244 20132 27300 20142
rect 27244 20038 27300 20076
rect 27468 18676 27524 21308
rect 27468 18340 27524 18620
rect 27468 18274 27524 18284
rect 27692 15148 27748 24892
rect 27804 24836 27860 30268
rect 28252 30212 28308 30222
rect 28252 30118 28308 30156
rect 28028 30100 28084 30110
rect 28084 30044 28196 30100
rect 28028 30034 28084 30044
rect 28028 29314 28084 29326
rect 28028 29262 28030 29314
rect 28082 29262 28084 29314
rect 28028 28420 28084 29262
rect 28028 27858 28084 28364
rect 28028 27806 28030 27858
rect 28082 27806 28084 27858
rect 28028 27794 28084 27806
rect 28140 26962 28196 30044
rect 28252 29538 28308 29550
rect 28252 29486 28254 29538
rect 28306 29486 28308 29538
rect 28252 28644 28308 29486
rect 28252 28578 28308 28588
rect 28252 27076 28308 27086
rect 28364 27076 28420 33964
rect 28588 33954 28644 33964
rect 28700 31892 28756 35534
rect 28476 31836 28756 31892
rect 28476 31444 28532 31836
rect 28588 31668 28644 31678
rect 28644 31612 28756 31668
rect 28588 31574 28644 31612
rect 28476 31388 28644 31444
rect 28476 30994 28532 31006
rect 28476 30942 28478 30994
rect 28530 30942 28532 30994
rect 28476 30884 28532 30942
rect 28476 30818 28532 30828
rect 28476 30210 28532 30222
rect 28476 30158 28478 30210
rect 28530 30158 28532 30210
rect 28476 30100 28532 30158
rect 28476 30034 28532 30044
rect 28476 27972 28532 27982
rect 28476 27858 28532 27916
rect 28476 27806 28478 27858
rect 28530 27806 28532 27858
rect 28476 27794 28532 27806
rect 28252 27074 28420 27076
rect 28252 27022 28254 27074
rect 28306 27022 28420 27074
rect 28252 27020 28420 27022
rect 28252 27010 28308 27020
rect 28140 26910 28142 26962
rect 28194 26910 28196 26962
rect 28140 26908 28196 26910
rect 27916 26850 27972 26862
rect 27916 26798 27918 26850
rect 27970 26798 27972 26850
rect 27916 26292 27972 26798
rect 28028 26852 28196 26908
rect 28588 26908 28644 31388
rect 28700 30436 28756 31612
rect 28812 31220 28868 31230
rect 28812 30994 28868 31164
rect 28812 30942 28814 30994
rect 28866 30942 28868 30994
rect 28812 30930 28868 30942
rect 28924 30996 28980 38220
rect 29036 35028 29092 38332
rect 29148 37940 29204 37950
rect 29372 37940 29428 38782
rect 29596 38052 29652 38090
rect 29596 37986 29652 37996
rect 29820 38050 29876 38894
rect 30268 39788 30548 39844
rect 30268 38668 30324 39788
rect 30716 39732 30772 39742
rect 30604 39676 30716 39732
rect 30492 38722 30548 38734
rect 30492 38670 30494 38722
rect 30546 38670 30548 38722
rect 30492 38668 30548 38670
rect 29820 37998 29822 38050
rect 29874 37998 29876 38050
rect 29820 37986 29876 37998
rect 29932 38612 30324 38668
rect 30380 38612 30548 38668
rect 29932 38050 29988 38612
rect 29932 37998 29934 38050
rect 29986 37998 29988 38050
rect 29484 37940 29540 37950
rect 29372 37938 29540 37940
rect 29372 37886 29486 37938
rect 29538 37886 29540 37938
rect 29372 37884 29540 37886
rect 29148 35812 29204 37884
rect 29260 37156 29316 37166
rect 29260 37062 29316 37100
rect 29484 37156 29540 37884
rect 29932 37940 29988 37998
rect 29932 37874 29988 37884
rect 30044 38052 30100 38062
rect 29596 37828 29652 37838
rect 29596 37268 29652 37772
rect 29596 37174 29652 37212
rect 30044 37156 30100 37996
rect 29484 37090 29540 37100
rect 29932 37100 30100 37156
rect 30156 37154 30212 37166
rect 30156 37102 30158 37154
rect 30210 37102 30212 37154
rect 29932 36594 29988 37100
rect 30156 37044 30212 37102
rect 30156 36978 30212 36988
rect 29932 36542 29934 36594
rect 29986 36542 29988 36594
rect 29932 36530 29988 36542
rect 30044 36932 30100 36942
rect 30044 36482 30100 36876
rect 30044 36430 30046 36482
rect 30098 36430 30100 36482
rect 29372 35812 29428 35822
rect 29148 35810 29428 35812
rect 29148 35758 29374 35810
rect 29426 35758 29428 35810
rect 29148 35756 29428 35758
rect 29372 35746 29428 35756
rect 29484 35810 29540 35822
rect 29484 35758 29486 35810
rect 29538 35758 29540 35810
rect 29484 35700 29540 35758
rect 29932 35812 29988 35822
rect 29932 35718 29988 35756
rect 29484 35634 29540 35644
rect 30044 35700 30100 36430
rect 30044 35634 30100 35644
rect 30156 36708 30212 36718
rect 29484 35476 29540 35486
rect 30044 35476 30100 35486
rect 29484 35474 29652 35476
rect 29484 35422 29486 35474
rect 29538 35422 29652 35474
rect 29484 35420 29652 35422
rect 29484 35410 29540 35420
rect 29036 34962 29092 34972
rect 29484 34804 29540 34814
rect 29260 34690 29316 34702
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29036 34580 29092 34590
rect 29036 34354 29092 34524
rect 29260 34580 29316 34638
rect 29260 34514 29316 34524
rect 29036 34302 29038 34354
rect 29090 34302 29092 34354
rect 29036 34290 29092 34302
rect 29484 34354 29540 34748
rect 29484 34302 29486 34354
rect 29538 34302 29540 34354
rect 29484 34290 29540 34302
rect 29260 32564 29316 32574
rect 29260 31890 29316 32508
rect 29260 31838 29262 31890
rect 29314 31838 29316 31890
rect 29260 31826 29316 31838
rect 29484 31668 29540 31678
rect 29484 31574 29540 31612
rect 29036 30996 29092 31006
rect 28924 30940 29036 30996
rect 29036 30902 29092 30940
rect 28700 30370 28756 30380
rect 29148 30770 29204 30782
rect 29148 30718 29150 30770
rect 29202 30718 29204 30770
rect 29148 30212 29204 30718
rect 29260 30212 29316 30222
rect 29148 30156 29260 30212
rect 29260 30098 29316 30156
rect 29260 30046 29262 30098
rect 29314 30046 29316 30098
rect 29260 30034 29316 30046
rect 29372 30100 29428 30110
rect 29372 30006 29428 30044
rect 29036 29988 29092 29998
rect 28700 29986 29092 29988
rect 28700 29934 29038 29986
rect 29090 29934 29092 29986
rect 28700 29932 29092 29934
rect 28700 28642 28756 29932
rect 29036 29922 29092 29932
rect 29596 29876 29652 35420
rect 29596 29810 29652 29820
rect 29708 35364 29764 35374
rect 29708 29652 29764 35308
rect 29932 35140 29988 35150
rect 29820 34804 29876 34814
rect 29820 34710 29876 34748
rect 29932 33346 29988 35084
rect 29932 33294 29934 33346
rect 29986 33294 29988 33346
rect 29932 33282 29988 33294
rect 30044 32676 30100 35420
rect 30156 34020 30212 36652
rect 30380 35140 30436 38612
rect 30492 37828 30548 37838
rect 30492 37734 30548 37772
rect 30492 36370 30548 36382
rect 30492 36318 30494 36370
rect 30546 36318 30548 36370
rect 30492 35474 30548 36318
rect 30492 35422 30494 35474
rect 30546 35422 30548 35474
rect 30492 35410 30548 35422
rect 30492 35140 30548 35150
rect 30380 35084 30492 35140
rect 30492 35074 30548 35084
rect 30156 33954 30212 33964
rect 30604 33572 30660 39676
rect 30716 39666 30772 39676
rect 30828 38668 30884 40012
rect 30940 38948 30996 38958
rect 30940 38854 30996 38892
rect 31052 38668 31108 40796
rect 30716 38612 30884 38668
rect 30940 38612 31108 38668
rect 31164 40404 31220 40414
rect 30716 37938 30772 38612
rect 30716 37886 30718 37938
rect 30770 37886 30772 37938
rect 30716 37874 30772 37886
rect 30828 37938 30884 37950
rect 30828 37886 30830 37938
rect 30882 37886 30884 37938
rect 30828 37268 30884 37886
rect 30828 37202 30884 37212
rect 30828 37042 30884 37054
rect 30828 36990 30830 37042
rect 30882 36990 30884 37042
rect 30716 35700 30772 35710
rect 30716 34804 30772 35644
rect 30828 35028 30884 36990
rect 30940 36594 30996 38612
rect 30940 36542 30942 36594
rect 30994 36542 30996 36594
rect 30940 35252 30996 36542
rect 31052 37156 31108 37166
rect 31052 36372 31108 37100
rect 31164 36596 31220 40348
rect 31276 38164 31332 44156
rect 31500 41972 31556 41982
rect 31500 41878 31556 41916
rect 31388 41076 31444 41086
rect 31388 40982 31444 41020
rect 31612 40964 31668 40974
rect 31500 40962 31668 40964
rect 31500 40910 31614 40962
rect 31666 40910 31668 40962
rect 31500 40908 31668 40910
rect 31388 40852 31444 40862
rect 31388 40402 31444 40796
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31388 40338 31444 40350
rect 31500 39732 31556 40908
rect 31612 40898 31668 40908
rect 31612 40740 31668 40750
rect 31612 40402 31668 40684
rect 31612 40350 31614 40402
rect 31666 40350 31668 40402
rect 31612 40338 31668 40350
rect 31500 39666 31556 39676
rect 31724 38948 31780 47516
rect 31948 46004 32004 49534
rect 32060 49140 32116 49150
rect 32060 49046 32116 49084
rect 32284 47348 32340 50372
rect 32508 49252 32564 50542
rect 32620 49812 32676 51660
rect 32732 50482 32788 51884
rect 32732 50430 32734 50482
rect 32786 50430 32788 50482
rect 32732 50418 32788 50430
rect 32844 51380 32900 51390
rect 32732 49812 32788 49822
rect 32620 49756 32732 49812
rect 32732 49746 32788 49756
rect 32508 49196 32788 49252
rect 32620 49028 32676 49038
rect 32396 48916 32452 48926
rect 32396 48822 32452 48860
rect 32284 47282 32340 47292
rect 31948 45948 32564 46004
rect 32060 45780 32116 45790
rect 32116 45724 32228 45780
rect 32060 45686 32116 45724
rect 32060 45220 32116 45230
rect 32060 45126 32116 45164
rect 31836 45108 31892 45118
rect 31836 45014 31892 45052
rect 31948 44994 32004 45006
rect 31948 44942 31950 44994
rect 32002 44942 32004 44994
rect 31836 44322 31892 44334
rect 31836 44270 31838 44322
rect 31890 44270 31892 44322
rect 31836 44100 31892 44270
rect 31948 44324 32004 44942
rect 31948 44258 32004 44268
rect 32172 44100 32228 45724
rect 31836 44044 32228 44100
rect 32284 45556 32340 45566
rect 31948 43540 32004 44044
rect 31948 43484 32116 43540
rect 31948 42084 32004 42094
rect 31948 41970 32004 42028
rect 31948 41918 31950 41970
rect 32002 41918 32004 41970
rect 31948 41860 32004 41918
rect 31948 41794 32004 41804
rect 31836 41186 31892 41198
rect 31836 41134 31838 41186
rect 31890 41134 31892 41186
rect 31836 40628 31892 41134
rect 31948 40628 32004 40638
rect 31836 40572 31948 40628
rect 31948 40534 32004 40572
rect 32060 39956 32116 43484
rect 32284 40404 32340 45500
rect 32396 44436 32452 44446
rect 32396 44342 32452 44380
rect 32396 41972 32452 41982
rect 32396 41858 32452 41916
rect 32396 41806 32398 41858
rect 32450 41806 32452 41858
rect 32396 41300 32452 41806
rect 32396 41234 32452 41244
rect 32396 40740 32452 40750
rect 32396 40626 32452 40684
rect 32396 40574 32398 40626
rect 32450 40574 32452 40626
rect 32396 40562 32452 40574
rect 32396 40404 32452 40414
rect 32284 40348 32396 40404
rect 32508 40404 32564 45948
rect 32620 40852 32676 48972
rect 32732 48804 32788 49196
rect 32732 45668 32788 48748
rect 32732 45602 32788 45612
rect 32732 42530 32788 42542
rect 32732 42478 32734 42530
rect 32786 42478 32788 42530
rect 32732 41412 32788 42478
rect 32844 41972 32900 51324
rect 32956 50428 33012 53340
rect 33404 53060 33460 53070
rect 33404 52276 33460 53004
rect 33292 52220 33404 52276
rect 33292 51044 33348 52220
rect 33404 52210 33460 52220
rect 33516 51268 33572 53340
rect 33964 53172 34020 53182
rect 34300 53172 34356 63084
rect 34412 63084 34580 63140
rect 34636 63812 34692 63822
rect 34412 56308 34468 63084
rect 34524 60674 34580 60686
rect 34524 60622 34526 60674
rect 34578 60622 34580 60674
rect 34524 60562 34580 60622
rect 34524 60510 34526 60562
rect 34578 60510 34580 60562
rect 34524 60498 34580 60510
rect 34636 56308 34692 63756
rect 34860 60900 34916 60910
rect 34860 60806 34916 60844
rect 34748 60788 34804 60798
rect 34748 60694 34804 60732
rect 34972 60788 35028 60798
rect 34860 60004 34916 60014
rect 34860 59910 34916 59948
rect 34972 59556 35028 60732
rect 34972 59490 35028 59500
rect 34972 56308 35028 56318
rect 34412 56252 34580 56308
rect 34636 56306 35028 56308
rect 34636 56254 34974 56306
rect 35026 56254 35028 56306
rect 34636 56252 35028 56254
rect 34412 55300 34468 55310
rect 34412 55206 34468 55244
rect 33964 53170 34356 53172
rect 33964 53118 33966 53170
rect 34018 53118 34356 53170
rect 33964 53116 34356 53118
rect 33964 53106 34020 53116
rect 33740 53060 33796 53070
rect 33740 52966 33796 53004
rect 33628 52946 33684 52958
rect 33628 52894 33630 52946
rect 33682 52894 33684 52946
rect 33628 52724 33684 52894
rect 34300 52834 34356 52846
rect 34300 52782 34302 52834
rect 34354 52782 34356 52834
rect 34300 52724 34356 52782
rect 33684 52668 33796 52724
rect 33628 52658 33684 52668
rect 33628 51268 33684 51278
rect 33516 51266 33684 51268
rect 33516 51214 33630 51266
rect 33682 51214 33684 51266
rect 33516 51212 33684 51214
rect 33180 50988 33348 51044
rect 33180 50484 33236 50988
rect 33292 50818 33348 50830
rect 33292 50766 33294 50818
rect 33346 50766 33348 50818
rect 33292 50708 33348 50766
rect 33292 50642 33348 50652
rect 33292 50484 33348 50494
rect 33180 50482 33348 50484
rect 33180 50430 33294 50482
rect 33346 50430 33348 50482
rect 33180 50428 33348 50430
rect 32956 50372 33124 50428
rect 33068 50148 33124 50372
rect 33180 50372 33236 50428
rect 33292 50418 33348 50428
rect 33404 50484 33460 50494
rect 33628 50484 33684 51212
rect 33404 50482 33684 50484
rect 33404 50430 33406 50482
rect 33458 50430 33684 50482
rect 33404 50428 33684 50430
rect 33740 50428 33796 52668
rect 34300 52658 34356 52668
rect 34412 51380 34468 51390
rect 33964 50708 34020 50718
rect 33964 50614 34020 50652
rect 34300 50594 34356 50606
rect 34300 50542 34302 50594
rect 34354 50542 34356 50594
rect 33180 50306 33236 50316
rect 33404 50372 33460 50428
rect 33740 50372 33908 50428
rect 33404 50306 33460 50316
rect 33068 50092 33348 50148
rect 33180 49978 33236 49990
rect 33180 49926 33182 49978
rect 33234 49926 33236 49978
rect 33068 49812 33124 49822
rect 32956 48916 33012 48926
rect 32956 48822 33012 48860
rect 33068 47796 33124 49756
rect 33068 47730 33124 47740
rect 33180 49700 33236 49926
rect 32956 47682 33012 47694
rect 32956 47630 32958 47682
rect 33010 47630 33012 47682
rect 32956 47572 33012 47630
rect 32956 47506 33012 47516
rect 32956 47348 33012 47358
rect 32956 47254 33012 47292
rect 33068 47346 33124 47358
rect 33068 47294 33070 47346
rect 33122 47294 33124 47346
rect 33068 45108 33124 47294
rect 33180 46788 33236 49644
rect 33292 49028 33348 50092
rect 33404 49924 33460 49934
rect 33404 49830 33460 49868
rect 33740 49812 33796 49822
rect 33740 49718 33796 49756
rect 33292 48972 33460 49028
rect 33292 48804 33348 48814
rect 33292 48710 33348 48748
rect 33180 46722 33236 46732
rect 33404 45892 33460 48972
rect 33628 48916 33684 48926
rect 33628 48822 33684 48860
rect 33852 48356 33908 50372
rect 33852 48290 33908 48300
rect 34188 50372 34244 50382
rect 33628 47572 33684 47582
rect 33628 47478 33684 47516
rect 33852 47460 33908 47470
rect 33908 47404 34020 47460
rect 33852 47366 33908 47404
rect 33852 47124 33908 47134
rect 33628 46788 33684 46798
rect 33740 46788 33796 46798
rect 33684 46786 33796 46788
rect 33684 46734 33742 46786
rect 33794 46734 33796 46786
rect 33684 46732 33796 46734
rect 33404 45836 33572 45892
rect 33068 42978 33124 45052
rect 33068 42926 33070 42978
rect 33122 42926 33124 42978
rect 33068 42914 33124 42926
rect 33404 45668 33460 45678
rect 33292 42756 33348 42766
rect 33180 42754 33348 42756
rect 33180 42702 33294 42754
rect 33346 42702 33348 42754
rect 33180 42700 33348 42702
rect 33180 42084 33236 42700
rect 33292 42690 33348 42700
rect 33404 42420 33460 45612
rect 33516 42644 33572 45836
rect 33628 45444 33684 46732
rect 33740 46722 33796 46732
rect 33852 46786 33908 47068
rect 33852 46734 33854 46786
rect 33906 46734 33908 46786
rect 33852 46722 33908 46734
rect 33740 46452 33796 46462
rect 33964 46452 34020 47404
rect 33740 46450 34020 46452
rect 33740 46398 33742 46450
rect 33794 46398 34020 46450
rect 33740 46396 34020 46398
rect 33740 46386 33796 46396
rect 34188 45668 34244 50316
rect 34300 49924 34356 50542
rect 34300 49830 34356 49868
rect 34300 48804 34356 48814
rect 34412 48804 34468 51324
rect 34524 50932 34580 56252
rect 34972 56242 35028 56252
rect 34636 56082 34692 56094
rect 34636 56030 34638 56082
rect 34690 56030 34692 56082
rect 34636 55300 34692 56030
rect 34636 55234 34692 55244
rect 34748 55076 34804 55086
rect 34636 55074 34804 55076
rect 34636 55022 34750 55074
rect 34802 55022 34804 55074
rect 34636 55020 34804 55022
rect 34636 54514 34692 55020
rect 34748 55010 34804 55020
rect 34636 54462 34638 54514
rect 34690 54462 34692 54514
rect 34636 54450 34692 54462
rect 34972 52388 35028 52398
rect 35084 52388 35140 64540
rect 35196 64530 35252 64540
rect 35756 64036 35812 64046
rect 35644 63980 35756 64036
rect 35644 63922 35700 63980
rect 35644 63870 35646 63922
rect 35698 63870 35700 63922
rect 35644 63858 35700 63870
rect 35196 63812 35252 63822
rect 35196 63718 35252 63756
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35756 63362 35812 63980
rect 35756 63310 35758 63362
rect 35810 63310 35812 63362
rect 35756 63298 35812 63310
rect 35420 63140 35476 63150
rect 35420 63046 35476 63084
rect 35196 63028 35252 63038
rect 35196 62934 35252 62972
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35756 60898 35812 60910
rect 35756 60846 35758 60898
rect 35810 60846 35812 60898
rect 35308 60788 35364 60798
rect 35644 60788 35700 60798
rect 35308 60786 35700 60788
rect 35308 60734 35310 60786
rect 35362 60734 35646 60786
rect 35698 60734 35700 60786
rect 35308 60732 35700 60734
rect 35308 60564 35364 60732
rect 35644 60722 35700 60732
rect 35756 60788 35812 60846
rect 35756 60722 35812 60732
rect 35308 60498 35364 60508
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 60228 35252 60238
rect 35196 59890 35252 60172
rect 35196 59838 35198 59890
rect 35250 59838 35252 59890
rect 35196 59826 35252 59838
rect 35868 59332 35924 65550
rect 36092 65490 36148 66334
rect 36092 65438 36094 65490
rect 36146 65438 36148 65490
rect 36092 63810 36148 65438
rect 36428 65378 36484 68572
rect 36876 65716 36932 69244
rect 37324 69234 37380 69244
rect 37772 69188 37828 70140
rect 39004 70306 39060 70318
rect 39004 70254 39006 70306
rect 39058 70254 39060 70306
rect 39004 70196 39060 70254
rect 39004 70130 39060 70140
rect 37996 69972 38052 69982
rect 37996 69522 38052 69916
rect 38780 69972 38836 69982
rect 38780 69878 38836 69916
rect 39116 69748 39172 70700
rect 40348 70756 40404 73948
rect 42028 72324 42084 76302
rect 45500 76354 45556 76366
rect 45500 76302 45502 76354
rect 45554 76302 45556 76354
rect 42028 72258 42084 72268
rect 44380 75012 44436 75022
rect 40348 70690 40404 70700
rect 41804 70308 41860 70318
rect 39564 70196 39620 70206
rect 39564 70102 39620 70140
rect 41692 70196 41748 70206
rect 39004 69692 39172 69748
rect 38444 69636 38500 69646
rect 38444 69542 38500 69580
rect 37996 69470 37998 69522
rect 38050 69470 38052 69522
rect 37996 69458 38052 69470
rect 39004 69524 39060 69692
rect 37772 69122 37828 69132
rect 38668 68628 38724 68638
rect 38668 68534 38724 68572
rect 37436 68516 37492 68526
rect 37436 67228 37492 68460
rect 38780 68404 38836 68414
rect 38780 68310 38836 68348
rect 39004 67228 39060 69468
rect 39116 69522 39172 69534
rect 39116 69470 39118 69522
rect 39170 69470 39172 69522
rect 39116 68514 39172 69470
rect 39228 69412 39284 69422
rect 39228 69410 39844 69412
rect 39228 69358 39230 69410
rect 39282 69358 39844 69410
rect 39228 69356 39844 69358
rect 39228 69346 39284 69356
rect 39116 68462 39118 68514
rect 39170 68462 39172 68514
rect 39116 67842 39172 68462
rect 39116 67790 39118 67842
rect 39170 67790 39172 67842
rect 39116 67778 39172 67790
rect 39228 68628 39284 68638
rect 36428 65326 36430 65378
rect 36482 65326 36484 65378
rect 36428 65314 36484 65326
rect 36540 65660 36932 65716
rect 37324 67172 37492 67228
rect 38892 67172 39060 67228
rect 39228 67282 39284 68572
rect 39564 68628 39620 68638
rect 39564 68534 39620 68572
rect 39788 67954 39844 69356
rect 40012 68516 40068 68526
rect 40012 68514 40516 68516
rect 40012 68462 40014 68514
rect 40066 68462 40516 68514
rect 40012 68460 40516 68462
rect 40012 68450 40068 68460
rect 39788 67902 39790 67954
rect 39842 67902 39844 67954
rect 39340 67844 39396 67854
rect 39676 67844 39732 67854
rect 39340 67842 39732 67844
rect 39340 67790 39342 67842
rect 39394 67790 39678 67842
rect 39730 67790 39732 67842
rect 39340 67788 39732 67790
rect 39340 67778 39396 67788
rect 39676 67778 39732 67788
rect 39228 67230 39230 67282
rect 39282 67230 39284 67282
rect 39228 67218 39284 67230
rect 39788 67228 39844 67902
rect 39340 67172 39844 67228
rect 40460 67954 40516 68460
rect 40460 67902 40462 67954
rect 40514 67902 40516 67954
rect 40460 67228 40516 67902
rect 40572 68404 40628 68414
rect 40572 67842 40628 68348
rect 40572 67790 40574 67842
rect 40626 67790 40628 67842
rect 40572 67778 40628 67790
rect 40908 67732 40964 67742
rect 40908 67638 40964 67676
rect 41692 67228 41748 70140
rect 41804 69522 41860 70252
rect 41804 69470 41806 69522
rect 41858 69470 41860 69522
rect 41804 69458 41860 69470
rect 42252 69410 42308 69422
rect 42252 69358 42254 69410
rect 42306 69358 42308 69410
rect 42252 67732 42308 69358
rect 42700 69412 42756 69422
rect 42700 69410 43204 69412
rect 42700 69358 42702 69410
rect 42754 69358 43204 69410
rect 42700 69356 43204 69358
rect 42700 69346 42756 69356
rect 42252 67666 42308 67676
rect 43148 67842 43204 69356
rect 43148 67790 43150 67842
rect 43202 67790 43204 67842
rect 43148 67228 43204 67790
rect 43596 67732 43652 67742
rect 43596 67638 43652 67676
rect 43820 67730 43876 67742
rect 43820 67678 43822 67730
rect 43874 67678 43876 67730
rect 40460 67172 41076 67228
rect 41692 67172 41860 67228
rect 37324 65716 37380 67172
rect 37548 66498 37604 66510
rect 37548 66446 37550 66498
rect 37602 66446 37604 66498
rect 37548 66388 37604 66446
rect 37548 66322 37604 66332
rect 38556 66386 38612 66398
rect 38556 66334 38558 66386
rect 38610 66334 38612 66386
rect 37436 66276 37492 66286
rect 37436 66164 37492 66220
rect 38332 66276 38388 66286
rect 37548 66164 37604 66174
rect 37436 66108 37548 66164
rect 37548 66070 37604 66108
rect 37660 66164 37716 66174
rect 37660 66162 37828 66164
rect 37660 66110 37662 66162
rect 37714 66110 37828 66162
rect 37660 66108 37828 66110
rect 37660 66098 37716 66108
rect 37324 65660 37604 65716
rect 36092 63758 36094 63810
rect 36146 63758 36148 63810
rect 36092 63746 36148 63758
rect 36428 63812 36484 63822
rect 36428 63718 36484 63756
rect 36316 60898 36372 60910
rect 36316 60846 36318 60898
rect 36370 60846 36372 60898
rect 35980 60788 36036 60798
rect 36204 60788 36260 60798
rect 35980 60786 36260 60788
rect 35980 60734 35982 60786
rect 36034 60734 36206 60786
rect 36258 60734 36260 60786
rect 35980 60732 36260 60734
rect 35980 60722 36036 60732
rect 36204 60722 36260 60732
rect 36316 60788 36372 60846
rect 36316 60722 36372 60732
rect 36316 60564 36372 60574
rect 36316 60470 36372 60508
rect 35980 59778 36036 59790
rect 35980 59726 35982 59778
rect 36034 59726 36036 59778
rect 35980 59556 36036 59726
rect 35980 59490 36036 59500
rect 36316 59778 36372 59790
rect 36316 59726 36318 59778
rect 36370 59726 36372 59778
rect 35868 59276 36148 59332
rect 35644 59220 35700 59230
rect 35644 59126 35700 59164
rect 35980 59108 36036 59118
rect 35980 59014 36036 59052
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35756 56868 35812 56878
rect 35644 56866 35812 56868
rect 35644 56814 35758 56866
rect 35810 56814 35812 56866
rect 35644 56812 35812 56814
rect 35644 56308 35700 56812
rect 35756 56802 35812 56812
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35532 55412 35588 55422
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35532 53396 35588 55356
rect 35644 54852 35700 56252
rect 35756 56644 35812 56654
rect 35756 55522 35812 56588
rect 35756 55470 35758 55522
rect 35810 55470 35812 55522
rect 35756 55458 35812 55470
rect 35868 55970 35924 55982
rect 35868 55918 35870 55970
rect 35922 55918 35924 55970
rect 35868 55188 35924 55918
rect 35868 55186 36036 55188
rect 35868 55134 35870 55186
rect 35922 55134 36036 55186
rect 35868 55132 36036 55134
rect 35868 55122 35924 55132
rect 35756 55076 35812 55086
rect 35756 54982 35812 55020
rect 35644 54796 35924 54852
rect 35532 53330 35588 53340
rect 35868 53058 35924 54796
rect 35868 53006 35870 53058
rect 35922 53006 35924 53058
rect 35868 52994 35924 53006
rect 35644 52948 35700 52958
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34972 52386 35140 52388
rect 34972 52334 34974 52386
rect 35026 52334 35140 52386
rect 34972 52332 35140 52334
rect 34972 52322 35028 52332
rect 35084 52164 35140 52174
rect 34524 50866 34580 50876
rect 34636 52162 35140 52164
rect 34636 52110 35086 52162
rect 35138 52110 35140 52162
rect 34636 52108 35140 52110
rect 34636 51938 34692 52108
rect 35084 52098 35140 52108
rect 35532 52162 35588 52174
rect 35532 52110 35534 52162
rect 35586 52110 35588 52162
rect 34636 51886 34638 51938
rect 34690 51886 34692 51938
rect 34524 50708 34580 50718
rect 34524 49810 34580 50652
rect 34524 49758 34526 49810
rect 34578 49758 34580 49810
rect 34524 49746 34580 49758
rect 34412 48748 34580 48804
rect 34300 48468 34356 48748
rect 34412 48468 34468 48478
rect 34300 48466 34468 48468
rect 34300 48414 34414 48466
rect 34466 48414 34468 48466
rect 34300 48412 34468 48414
rect 34412 48402 34468 48412
rect 34524 48242 34580 48748
rect 34524 48190 34526 48242
rect 34578 48190 34580 48242
rect 34412 48132 34468 48142
rect 34300 48020 34356 48030
rect 34300 47572 34356 47964
rect 34412 48018 34468 48076
rect 34412 47966 34414 48018
rect 34466 47966 34468 48018
rect 34412 47954 34468 47966
rect 34412 47572 34468 47582
rect 34300 47570 34468 47572
rect 34300 47518 34414 47570
rect 34466 47518 34468 47570
rect 34300 47516 34468 47518
rect 34412 46674 34468 47516
rect 34412 46622 34414 46674
rect 34466 46622 34468 46674
rect 34412 46610 34468 46622
rect 34524 46676 34580 48190
rect 34524 46610 34580 46620
rect 34636 46452 34692 51886
rect 34972 51940 35028 51950
rect 34972 51846 35028 51884
rect 35532 51940 35588 52110
rect 35532 51602 35588 51884
rect 35532 51550 35534 51602
rect 35586 51550 35588 51602
rect 35532 51538 35588 51550
rect 35420 51380 35476 51390
rect 35420 51286 35476 51324
rect 35532 51156 35588 51166
rect 35644 51156 35700 52892
rect 35756 52162 35812 52174
rect 35756 52110 35758 52162
rect 35810 52110 35812 52162
rect 35756 51268 35812 52110
rect 35756 51202 35812 51212
rect 35532 51154 35700 51156
rect 35532 51102 35534 51154
rect 35586 51102 35700 51154
rect 35532 51100 35700 51102
rect 35532 51090 35588 51100
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35980 50818 36036 55132
rect 36092 52386 36148 59276
rect 36316 58996 36372 59726
rect 36428 59220 36484 59230
rect 36428 59126 36484 59164
rect 36316 58930 36372 58940
rect 36428 56980 36484 56990
rect 36540 56980 36596 65660
rect 36764 65490 36820 65502
rect 36764 65438 36766 65490
rect 36818 65438 36820 65490
rect 36652 64036 36708 64046
rect 36652 63942 36708 63980
rect 36764 63810 36820 65438
rect 36764 63758 36766 63810
rect 36818 63758 36820 63810
rect 36764 63746 36820 63758
rect 36876 65492 36932 65502
rect 36876 63588 36932 65436
rect 36764 63532 36932 63588
rect 37436 65490 37492 65502
rect 37436 65438 37438 65490
rect 37490 65438 37492 65490
rect 36764 62578 36820 63532
rect 36764 62526 36766 62578
rect 36818 62526 36820 62578
rect 36764 62514 36820 62526
rect 37436 62580 37492 65438
rect 37548 65380 37604 65660
rect 37660 65492 37716 65502
rect 37660 65398 37716 65436
rect 37548 64818 37604 65324
rect 37548 64766 37550 64818
rect 37602 64766 37604 64818
rect 37548 64754 37604 64766
rect 37772 64820 37828 66108
rect 38332 65714 38388 66220
rect 38332 65662 38334 65714
rect 38386 65662 38388 65714
rect 38332 65650 38388 65662
rect 38444 66274 38500 66286
rect 38444 66222 38446 66274
rect 38498 66222 38500 66274
rect 38444 66164 38500 66222
rect 38444 65602 38500 66108
rect 38556 65828 38612 66334
rect 38556 65772 38724 65828
rect 38444 65550 38446 65602
rect 38498 65550 38500 65602
rect 38444 65538 38500 65550
rect 38668 65490 38724 65772
rect 38668 65438 38670 65490
rect 38722 65438 38724 65490
rect 37884 64820 37940 64830
rect 37772 64764 37884 64820
rect 37884 64726 37940 64764
rect 38220 64818 38276 64830
rect 38220 64766 38222 64818
rect 38274 64766 38276 64818
rect 38220 64148 38276 64766
rect 38668 64820 38724 65438
rect 38668 64754 38724 64764
rect 38556 64706 38612 64718
rect 38556 64654 38558 64706
rect 38610 64654 38612 64706
rect 38444 64148 38500 64158
rect 38220 64146 38500 64148
rect 38220 64094 38446 64146
rect 38498 64094 38500 64146
rect 38220 64092 38500 64094
rect 38444 64082 38500 64092
rect 37884 63922 37940 63934
rect 37884 63870 37886 63922
rect 37938 63870 37940 63922
rect 37884 63812 37940 63870
rect 37436 62524 37716 62580
rect 36988 62354 37044 62366
rect 36988 62302 36990 62354
rect 37042 62302 37044 62354
rect 36652 62132 36708 62142
rect 36652 62130 36820 62132
rect 36652 62078 36654 62130
rect 36706 62078 36820 62130
rect 36652 62076 36820 62078
rect 36652 62066 36708 62076
rect 36764 60900 36820 62076
rect 36988 61796 37044 62302
rect 37660 62188 37716 62524
rect 36876 61740 37044 61796
rect 37100 62132 37716 62188
rect 36876 61012 36932 61740
rect 37100 61684 37156 62132
rect 37884 61796 37940 63756
rect 38556 63924 38612 64654
rect 38780 63924 38836 63934
rect 38556 63868 38780 63924
rect 38108 63700 38164 63710
rect 38220 63700 38276 63710
rect 38108 63698 38220 63700
rect 38108 63646 38110 63698
rect 38162 63646 38220 63698
rect 38108 63644 38220 63646
rect 38108 63634 38164 63644
rect 36988 61628 37156 61684
rect 37660 61794 37940 61796
rect 37660 61742 37886 61794
rect 37938 61742 37940 61794
rect 37660 61740 37940 61742
rect 36988 61012 37044 61628
rect 37212 61572 37268 61582
rect 37548 61572 37604 61582
rect 37212 61570 37604 61572
rect 37212 61518 37214 61570
rect 37266 61518 37550 61570
rect 37602 61518 37604 61570
rect 37212 61516 37604 61518
rect 37212 61506 37268 61516
rect 37548 61506 37604 61516
rect 37100 61458 37156 61470
rect 37100 61406 37102 61458
rect 37154 61406 37156 61458
rect 37100 61236 37156 61406
rect 37660 61348 37716 61740
rect 37884 61730 37940 61740
rect 38108 61572 38164 61582
rect 37884 61570 38164 61572
rect 37884 61518 38110 61570
rect 38162 61518 38164 61570
rect 37884 61516 38164 61518
rect 37772 61460 37828 61470
rect 37772 61366 37828 61404
rect 37100 61170 37156 61180
rect 37212 61292 37716 61348
rect 37100 61012 37156 61022
rect 36988 61010 37156 61012
rect 36988 60958 37102 61010
rect 37154 60958 37156 61010
rect 36988 60956 37156 60958
rect 36876 60900 36932 60956
rect 37100 60946 37156 60956
rect 37212 61010 37268 61292
rect 37212 60958 37214 61010
rect 37266 60958 37268 61010
rect 37212 60946 37268 60958
rect 36876 60844 37044 60900
rect 36764 60806 36820 60844
rect 36988 60786 37044 60844
rect 36988 60734 36990 60786
rect 37042 60734 37044 60786
rect 36988 60722 37044 60734
rect 37212 60788 37268 60798
rect 37100 59892 37156 59902
rect 37100 59778 37156 59836
rect 37100 59726 37102 59778
rect 37154 59726 37156 59778
rect 37100 59668 37156 59726
rect 36428 56978 36596 56980
rect 36428 56926 36430 56978
rect 36482 56926 36596 56978
rect 36428 56924 36596 56926
rect 36764 59612 37156 59668
rect 36764 59108 36820 59612
rect 37100 59444 37156 59454
rect 37212 59444 37268 60732
rect 37324 60786 37380 60798
rect 37324 60734 37326 60786
rect 37378 60734 37380 60786
rect 37324 60564 37380 60734
rect 37324 60498 37380 60508
rect 37100 59442 37268 59444
rect 37100 59390 37102 59442
rect 37154 59390 37268 59442
rect 37100 59388 37268 59390
rect 37436 60002 37492 60014
rect 37436 59950 37438 60002
rect 37490 59950 37492 60002
rect 37100 59378 37156 59388
rect 36428 56914 36484 56924
rect 36316 56866 36372 56878
rect 36316 56814 36318 56866
rect 36370 56814 36372 56866
rect 36316 56196 36372 56814
rect 36652 56196 36708 56206
rect 36316 56140 36652 56196
rect 36652 56102 36708 56140
rect 36204 56082 36260 56094
rect 36204 56030 36206 56082
rect 36258 56030 36260 56082
rect 36204 55076 36260 56030
rect 36764 55972 36820 59052
rect 36876 59220 36932 59230
rect 36876 58772 36932 59164
rect 36988 59218 37044 59230
rect 36988 59166 36990 59218
rect 37042 59166 37044 59218
rect 36988 58996 37044 59166
rect 37212 59220 37268 59230
rect 37212 59126 37268 59164
rect 37324 59220 37380 59230
rect 37436 59220 37492 59950
rect 37884 60004 37940 61516
rect 38108 61506 38164 61516
rect 38220 60226 38276 63644
rect 38556 62188 38612 63868
rect 38780 63830 38836 63868
rect 38444 62132 38612 62188
rect 38892 62188 38948 67172
rect 39004 67060 39060 67070
rect 39004 66966 39060 67004
rect 39116 67058 39172 67070
rect 39116 67006 39118 67058
rect 39170 67006 39172 67058
rect 39116 66388 39172 67006
rect 39116 65716 39172 66332
rect 39340 66386 39396 67172
rect 41020 67170 41076 67172
rect 41020 67118 41022 67170
rect 41074 67118 41076 67170
rect 41020 67106 41076 67118
rect 39340 66334 39342 66386
rect 39394 66334 39396 66386
rect 39340 66322 39396 66334
rect 39452 67058 39508 67070
rect 39452 67006 39454 67058
rect 39506 67006 39508 67058
rect 39228 66276 39284 66286
rect 39228 66182 39284 66220
rect 39228 65716 39284 65726
rect 39452 65716 39508 67006
rect 39564 67060 39620 67070
rect 39620 67004 39732 67060
rect 39564 66994 39620 67004
rect 39116 65714 39284 65716
rect 39116 65662 39230 65714
rect 39282 65662 39284 65714
rect 39116 65660 39284 65662
rect 39228 65650 39284 65660
rect 39340 65714 39508 65716
rect 39340 65662 39454 65714
rect 39506 65662 39508 65714
rect 39340 65660 39508 65662
rect 39340 64146 39396 65660
rect 39452 65650 39508 65660
rect 39564 66162 39620 66174
rect 39564 66110 39566 66162
rect 39618 66110 39620 66162
rect 39564 65378 39620 66110
rect 39564 65326 39566 65378
rect 39618 65326 39620 65378
rect 39564 65314 39620 65326
rect 39676 65602 39732 67004
rect 41356 66946 41412 66958
rect 41356 66894 41358 66946
rect 41410 66894 41412 66946
rect 41356 66388 41412 66894
rect 41804 66388 41860 67172
rect 42924 67172 43204 67228
rect 43484 67618 43540 67630
rect 43484 67566 43486 67618
rect 43538 67566 43540 67618
rect 42924 67170 42980 67172
rect 42924 67118 42926 67170
rect 42978 67118 42980 67170
rect 42924 67106 42980 67118
rect 41916 67060 41972 67070
rect 42588 67060 42644 67070
rect 41916 67058 42420 67060
rect 41916 67006 41918 67058
rect 41970 67006 42420 67058
rect 41916 67004 42420 67006
rect 41916 66994 41972 67004
rect 41916 66388 41972 66398
rect 41804 66386 41972 66388
rect 41804 66334 41918 66386
rect 41970 66334 41972 66386
rect 41804 66332 41972 66334
rect 41356 66294 41412 66332
rect 40124 66052 40180 66062
rect 39676 65550 39678 65602
rect 39730 65550 39732 65602
rect 39676 64482 39732 65550
rect 40012 65996 40124 66052
rect 40012 65490 40068 65996
rect 40124 65986 40180 65996
rect 40572 66050 40628 66062
rect 40572 65998 40574 66050
rect 40626 65998 40628 66050
rect 40012 65438 40014 65490
rect 40066 65438 40068 65490
rect 40012 65426 40068 65438
rect 40236 65602 40292 65614
rect 40236 65550 40238 65602
rect 40290 65550 40292 65602
rect 39676 64430 39678 64482
rect 39730 64430 39732 64482
rect 39676 64418 39732 64430
rect 40012 65268 40068 65278
rect 40012 64706 40068 65212
rect 40012 64654 40014 64706
rect 40066 64654 40068 64706
rect 39340 64094 39342 64146
rect 39394 64094 39396 64146
rect 39340 64082 39396 64094
rect 39788 64148 39844 64158
rect 40012 64148 40068 64654
rect 40236 64708 40292 65550
rect 40348 65490 40404 65502
rect 40348 65438 40350 65490
rect 40402 65438 40404 65490
rect 40348 65268 40404 65438
rect 40572 65380 40628 65998
rect 41020 66052 41076 66062
rect 41244 66052 41300 66062
rect 41020 65958 41076 65996
rect 41132 66050 41300 66052
rect 41132 65998 41246 66050
rect 41298 65998 41300 66050
rect 41132 65996 41300 65998
rect 41132 65828 41188 65996
rect 41244 65986 41300 65996
rect 41468 66050 41524 66062
rect 41468 65998 41470 66050
rect 41522 65998 41524 66050
rect 41468 65828 41524 65998
rect 40572 65314 40628 65324
rect 41020 65772 41188 65828
rect 41244 65772 41524 65828
rect 41916 65828 41972 66332
rect 41020 65380 41076 65772
rect 41020 65314 41076 65324
rect 41132 65602 41188 65614
rect 41132 65550 41134 65602
rect 41186 65550 41188 65602
rect 40348 65202 40404 65212
rect 40908 65268 40964 65278
rect 40908 65174 40964 65212
rect 41132 64932 41188 65550
rect 41244 65378 41300 65772
rect 41916 65762 41972 65772
rect 41916 65604 41972 65614
rect 42028 65604 42084 67004
rect 42252 66388 42308 66398
rect 42252 66274 42308 66332
rect 42252 66222 42254 66274
rect 42306 66222 42308 66274
rect 42252 66210 42308 66222
rect 42364 66162 42420 67004
rect 42588 66274 42644 67004
rect 43372 67060 43428 67070
rect 43372 66966 43428 67004
rect 42588 66222 42590 66274
rect 42642 66222 42644 66274
rect 42588 66210 42644 66222
rect 43260 66946 43316 66958
rect 43260 66894 43262 66946
rect 43314 66894 43316 66946
rect 43260 66836 43316 66894
rect 42364 66110 42366 66162
rect 42418 66110 42420 66162
rect 42364 66098 42420 66110
rect 41916 65602 42084 65604
rect 41916 65550 41918 65602
rect 41970 65550 42084 65602
rect 41916 65548 42084 65550
rect 42364 65828 42420 65838
rect 41916 65538 41972 65548
rect 42364 65492 42420 65772
rect 42252 65490 42420 65492
rect 42252 65438 42366 65490
rect 42418 65438 42420 65490
rect 42252 65436 42420 65438
rect 41244 65326 41246 65378
rect 41298 65326 41300 65378
rect 41244 65314 41300 65326
rect 41356 65380 41412 65390
rect 40796 64876 41188 64932
rect 40684 64708 40740 64718
rect 40796 64708 40852 64876
rect 40236 64706 40852 64708
rect 40236 64654 40686 64706
rect 40738 64654 40852 64706
rect 40236 64652 40852 64654
rect 40684 64148 40740 64652
rect 40012 64092 40404 64148
rect 39788 64054 39844 64092
rect 39900 64034 39956 64046
rect 39900 63982 39902 64034
rect 39954 63982 39956 64034
rect 39900 63924 39956 63982
rect 39900 63858 39956 63868
rect 39004 63812 39060 63822
rect 39004 63718 39060 63756
rect 39676 63700 39732 63710
rect 39676 63606 39732 63644
rect 38892 62132 39396 62188
rect 38444 61010 38500 62132
rect 38444 60958 38446 61010
rect 38498 60958 38500 61010
rect 38444 60946 38500 60958
rect 38780 61570 38836 61582
rect 38780 61518 38782 61570
rect 38834 61518 38836 61570
rect 38668 60786 38724 60798
rect 38668 60734 38670 60786
rect 38722 60734 38724 60786
rect 38668 60340 38724 60734
rect 38668 60274 38724 60284
rect 38220 60174 38222 60226
rect 38274 60174 38276 60226
rect 38220 60162 38276 60174
rect 38780 60116 38836 61518
rect 37660 59892 37716 59902
rect 37660 59798 37716 59836
rect 37772 59444 37828 59454
rect 37884 59444 37940 59948
rect 38332 60060 38836 60116
rect 39116 60116 39172 60126
rect 38332 60002 38388 60060
rect 38332 59950 38334 60002
rect 38386 59950 38388 60002
rect 38332 59938 38388 59950
rect 37772 59442 37940 59444
rect 37772 59390 37774 59442
rect 37826 59390 37940 59442
rect 37772 59388 37940 59390
rect 37772 59378 37828 59388
rect 37324 59218 37492 59220
rect 37324 59166 37326 59218
rect 37378 59166 37492 59218
rect 37324 59164 37492 59166
rect 38108 59220 38164 59230
rect 38556 59220 38612 59230
rect 38164 59218 38612 59220
rect 38164 59166 38558 59218
rect 38610 59166 38612 59218
rect 38164 59164 38612 59166
rect 36988 58930 37044 58940
rect 36876 58716 37044 58772
rect 36988 58212 37044 58716
rect 36988 58146 37044 58156
rect 37324 57428 37380 59164
rect 38108 59126 38164 59164
rect 38556 59108 38612 59164
rect 37884 58322 37940 58334
rect 37884 58270 37886 58322
rect 37938 58270 37940 58322
rect 37884 58212 37940 58270
rect 37996 58212 38052 58222
rect 37884 58156 37996 58212
rect 37996 58146 38052 58156
rect 37324 57362 37380 57372
rect 38332 57762 38388 57774
rect 38332 57710 38334 57762
rect 38386 57710 38388 57762
rect 38332 57428 38388 57710
rect 38332 57362 38388 57372
rect 36204 55010 36260 55020
rect 36652 55916 36820 55972
rect 36988 56754 37044 56766
rect 36988 56702 36990 56754
rect 37042 56702 37044 56754
rect 36316 52948 36372 52958
rect 36316 52854 36372 52892
rect 36092 52334 36094 52386
rect 36146 52334 36148 52386
rect 36092 52322 36148 52334
rect 35980 50766 35982 50818
rect 36034 50766 36036 50818
rect 35980 50754 36036 50766
rect 36316 51268 36372 51278
rect 35308 50708 35364 50718
rect 35084 50706 35364 50708
rect 35084 50654 35310 50706
rect 35362 50654 35364 50706
rect 35084 50652 35364 50654
rect 34748 50484 34804 50494
rect 35084 50484 35140 50652
rect 35308 50642 35364 50652
rect 36316 50708 36372 51212
rect 36316 50642 36372 50652
rect 34748 50482 35140 50484
rect 34748 50430 34750 50482
rect 34802 50430 35140 50482
rect 34748 50428 35140 50430
rect 34748 50418 34804 50428
rect 34860 49588 34916 49598
rect 34860 49494 34916 49532
rect 35084 49026 35140 50428
rect 35756 50594 35812 50606
rect 35756 50542 35758 50594
rect 35810 50542 35812 50594
rect 35756 50034 35812 50542
rect 35756 49982 35758 50034
rect 35810 49982 35812 50034
rect 35756 49970 35812 49982
rect 35980 49924 36036 49934
rect 35868 49922 36036 49924
rect 35868 49870 35982 49922
rect 36034 49870 36036 49922
rect 35868 49868 36036 49870
rect 35868 49812 35924 49868
rect 35980 49858 36036 49868
rect 35532 49756 35924 49812
rect 36092 49812 36148 49822
rect 36092 49810 36260 49812
rect 36092 49758 36094 49810
rect 36146 49758 36260 49810
rect 36092 49756 36260 49758
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35084 48974 35086 49026
rect 35138 48974 35140 49026
rect 35084 48962 35140 48974
rect 34972 48916 35028 48926
rect 34860 48804 34916 48814
rect 34860 48710 34916 48748
rect 34972 48356 35028 48860
rect 35532 48916 35588 49756
rect 36092 49746 36148 49756
rect 36204 49700 36260 49756
rect 36540 49700 36596 49710
rect 36204 49698 36596 49700
rect 36204 49646 36542 49698
rect 36594 49646 36596 49698
rect 36204 49644 36596 49646
rect 35868 49588 35924 49598
rect 35868 49138 35924 49532
rect 35868 49086 35870 49138
rect 35922 49086 35924 49138
rect 35868 49074 35924 49086
rect 36092 49026 36148 49038
rect 36092 48974 36094 49026
rect 36146 48974 36148 49026
rect 35532 48822 35588 48860
rect 35644 48916 35700 48926
rect 36092 48916 36148 48974
rect 35644 48914 36148 48916
rect 35644 48862 35646 48914
rect 35698 48862 36148 48914
rect 35644 48860 36148 48862
rect 35644 48850 35700 48860
rect 35308 48804 35364 48814
rect 36204 48804 36260 49644
rect 36540 49634 36596 49644
rect 35308 48710 35364 48748
rect 36092 48748 36260 48804
rect 36428 48802 36484 48814
rect 36428 48750 36430 48802
rect 36482 48750 36484 48802
rect 35756 48692 35812 48702
rect 34972 48300 35140 48356
rect 34972 48132 35028 48142
rect 34972 48038 35028 48076
rect 34748 47572 34804 47582
rect 34748 47458 34804 47516
rect 34748 47406 34750 47458
rect 34802 47406 34804 47458
rect 34748 47394 34804 47406
rect 34972 47460 35028 47470
rect 34972 47366 35028 47404
rect 34860 47234 34916 47246
rect 35084 47236 35140 48300
rect 35196 48242 35252 48254
rect 35196 48190 35198 48242
rect 35250 48190 35252 48242
rect 35196 48020 35252 48190
rect 35196 47954 35252 47964
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34860 47182 34862 47234
rect 34914 47182 34916 47234
rect 34748 46676 34804 46686
rect 34748 46582 34804 46620
rect 34636 46386 34692 46396
rect 34860 46116 34916 47182
rect 34972 47180 35140 47236
rect 35196 47234 35252 47246
rect 35196 47182 35198 47234
rect 35250 47182 35252 47234
rect 34972 46898 35028 47180
rect 34972 46846 34974 46898
rect 35026 46846 35028 46898
rect 34972 46834 35028 46846
rect 35084 46900 35140 46910
rect 35196 46900 35252 47182
rect 35084 46898 35252 46900
rect 35084 46846 35086 46898
rect 35138 46846 35252 46898
rect 35084 46844 35252 46846
rect 35084 46834 35140 46844
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34748 46060 34916 46116
rect 34188 45612 34468 45668
rect 33628 45378 33684 45388
rect 34300 44996 34356 45006
rect 34076 44436 34132 44446
rect 34300 44436 34356 44940
rect 34076 44434 34244 44436
rect 34076 44382 34078 44434
rect 34130 44382 34244 44434
rect 34076 44380 34244 44382
rect 34076 44370 34132 44380
rect 34188 42868 34244 44380
rect 34300 44370 34356 44380
rect 34412 44324 34468 45612
rect 34748 45220 34804 46060
rect 35308 45332 35364 45342
rect 34748 45106 34804 45164
rect 35196 45276 35308 45332
rect 35196 45218 35252 45276
rect 35308 45266 35364 45276
rect 35196 45166 35198 45218
rect 35250 45166 35252 45218
rect 35196 45154 35252 45166
rect 35644 45220 35700 45230
rect 35644 45126 35700 45164
rect 34748 45054 34750 45106
rect 34802 45054 34804 45106
rect 34748 45042 34804 45054
rect 35532 45106 35588 45118
rect 35532 45054 35534 45106
rect 35586 45054 35588 45106
rect 35532 44996 35588 45054
rect 35532 44930 35588 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34412 44230 34468 44268
rect 34972 44324 35028 44334
rect 34972 44230 35028 44268
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34412 42868 34468 42878
rect 33516 42578 33572 42588
rect 33740 42866 34468 42868
rect 33740 42814 34414 42866
rect 34466 42814 34468 42866
rect 33740 42812 34468 42814
rect 33292 42364 33572 42420
rect 33292 42194 33348 42364
rect 33292 42142 33294 42194
rect 33346 42142 33348 42194
rect 33292 42130 33348 42142
rect 33404 42196 33460 42206
rect 33180 42018 33236 42028
rect 33404 42082 33460 42140
rect 33404 42030 33406 42082
rect 33458 42030 33460 42082
rect 33404 42018 33460 42030
rect 33068 41972 33124 41982
rect 32844 41906 32900 41916
rect 32956 41970 33124 41972
rect 32956 41918 33070 41970
rect 33122 41918 33124 41970
rect 32956 41916 33124 41918
rect 32732 41356 32900 41412
rect 32844 40964 32900 41356
rect 32956 41188 33012 41916
rect 33068 41906 33124 41916
rect 33292 41972 33348 41982
rect 33180 41860 33236 41870
rect 32956 41094 33012 41132
rect 33068 41298 33124 41310
rect 33068 41246 33070 41298
rect 33122 41246 33124 41298
rect 33068 40964 33124 41246
rect 32844 40908 33124 40964
rect 32620 40796 32900 40852
rect 32732 40404 32788 40414
rect 32508 40348 32676 40404
rect 32396 40338 32452 40348
rect 31724 38882 31780 38892
rect 31948 39900 32116 39956
rect 32284 40180 32340 40190
rect 32620 40180 32676 40348
rect 31276 38098 31332 38108
rect 31276 37266 31332 37278
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 36932 31332 37214
rect 31500 37266 31556 37278
rect 31500 37214 31502 37266
rect 31554 37214 31556 37266
rect 31500 37044 31556 37214
rect 31500 36978 31556 36988
rect 31836 37154 31892 37166
rect 31836 37102 31838 37154
rect 31890 37102 31892 37154
rect 31276 36866 31332 36876
rect 31836 36932 31892 37102
rect 31948 37156 32004 39900
rect 32060 39732 32116 39742
rect 32284 39732 32340 40124
rect 32508 40124 32676 40180
rect 32060 39730 32340 39732
rect 32060 39678 32062 39730
rect 32114 39678 32340 39730
rect 32060 39676 32340 39678
rect 32060 39666 32116 39676
rect 32284 39618 32340 39676
rect 32284 39566 32286 39618
rect 32338 39566 32340 39618
rect 32284 39554 32340 39566
rect 32396 40068 32452 40078
rect 32396 39394 32452 40012
rect 32396 39342 32398 39394
rect 32450 39342 32452 39394
rect 32396 39284 32452 39342
rect 32396 39218 32452 39228
rect 31948 37090 32004 37100
rect 32060 37044 32116 37054
rect 32396 37044 32452 37054
rect 32060 36950 32116 36988
rect 32284 37042 32452 37044
rect 32284 36990 32398 37042
rect 32450 36990 32452 37042
rect 32284 36988 32452 36990
rect 31836 36866 31892 36876
rect 31164 36540 31556 36596
rect 31164 36372 31220 36382
rect 31052 36370 31220 36372
rect 31052 36318 31166 36370
rect 31218 36318 31220 36370
rect 31052 36316 31220 36318
rect 30940 35186 30996 35196
rect 31052 35698 31108 35710
rect 31052 35646 31054 35698
rect 31106 35646 31108 35698
rect 31052 35028 31108 35646
rect 30828 34972 31108 35028
rect 31052 34916 31108 34972
rect 31052 34850 31108 34860
rect 31164 34914 31220 36316
rect 31388 35588 31444 35598
rect 31164 34862 31166 34914
rect 31218 34862 31220 34914
rect 31164 34850 31220 34862
rect 31276 35586 31444 35588
rect 31276 35534 31390 35586
rect 31442 35534 31444 35586
rect 31276 35532 31444 35534
rect 30828 34804 30884 34814
rect 30716 34802 30884 34804
rect 30716 34750 30830 34802
rect 30882 34750 30884 34802
rect 30716 34748 30884 34750
rect 30828 34738 30884 34748
rect 30268 33516 30660 33572
rect 30268 33124 30324 33516
rect 30380 33348 30436 33358
rect 30380 33346 30996 33348
rect 30380 33294 30382 33346
rect 30434 33294 30996 33346
rect 30380 33292 30996 33294
rect 30380 33282 30436 33292
rect 30268 33068 30436 33124
rect 30044 32620 30212 32676
rect 30044 32450 30100 32462
rect 30044 32398 30046 32450
rect 30098 32398 30100 32450
rect 29932 31780 29988 31790
rect 29932 31106 29988 31724
rect 29932 31054 29934 31106
rect 29986 31054 29988 31106
rect 29932 31042 29988 31054
rect 29820 30996 29876 31006
rect 29820 30324 29876 30940
rect 29932 30884 29988 30894
rect 30044 30884 30100 32398
rect 29988 30828 30100 30884
rect 29932 30818 29988 30828
rect 29932 30324 29988 30334
rect 29820 30322 29988 30324
rect 29820 30270 29934 30322
rect 29986 30270 29988 30322
rect 29820 30268 29988 30270
rect 29932 30258 29988 30268
rect 29708 29586 29764 29596
rect 30044 30100 30100 30110
rect 30044 29650 30100 30044
rect 30044 29598 30046 29650
rect 30098 29598 30100 29650
rect 30044 29586 30100 29598
rect 28700 28590 28702 28642
rect 28754 28590 28756 28642
rect 28700 28578 28756 28590
rect 29484 29428 29540 29438
rect 28588 26852 28868 26908
rect 28028 26786 28084 26796
rect 28700 26404 28756 26414
rect 27916 25394 27972 26236
rect 28140 26292 28196 26302
rect 28476 26292 28532 26302
rect 28140 26290 28532 26292
rect 28140 26238 28142 26290
rect 28194 26238 28478 26290
rect 28530 26238 28532 26290
rect 28140 26236 28532 26238
rect 28140 26226 28196 26236
rect 28476 26226 28532 26236
rect 28028 25508 28084 25518
rect 28028 25414 28084 25452
rect 28588 25508 28644 25518
rect 28700 25508 28756 26348
rect 28812 26180 28868 26852
rect 28924 26404 28980 26414
rect 28924 26310 28980 26348
rect 29036 26290 29092 26302
rect 29036 26238 29038 26290
rect 29090 26238 29092 26290
rect 28812 26124 28980 26180
rect 28588 25506 28756 25508
rect 28588 25454 28590 25506
rect 28642 25454 28756 25506
rect 28588 25452 28756 25454
rect 27916 25342 27918 25394
rect 27970 25342 27972 25394
rect 27916 25330 27972 25342
rect 28588 24948 28644 25452
rect 28700 24948 28756 24958
rect 28588 24946 28756 24948
rect 28588 24894 28702 24946
rect 28754 24894 28756 24946
rect 28588 24892 28756 24894
rect 28700 24882 28756 24892
rect 27804 24780 28308 24836
rect 28140 23492 28196 23502
rect 28140 23042 28196 23436
rect 28140 22990 28142 23042
rect 28194 22990 28196 23042
rect 28140 22978 28196 22990
rect 28028 21140 28084 21150
rect 28028 20690 28084 21084
rect 28028 20638 28030 20690
rect 28082 20638 28084 20690
rect 28028 20626 28084 20638
rect 28140 20692 28196 20702
rect 28140 20598 28196 20636
rect 27804 20580 27860 20590
rect 27804 20486 27860 20524
rect 27916 19908 27972 19918
rect 27916 19814 27972 19852
rect 28028 16212 28084 16222
rect 27468 15092 27748 15148
rect 27916 16210 28084 16212
rect 27916 16158 28030 16210
rect 28082 16158 28084 16210
rect 27916 16156 28084 16158
rect 27916 15540 27972 16156
rect 28028 16146 28084 16156
rect 27468 14644 27524 15092
rect 27468 14642 27636 14644
rect 27468 14590 27470 14642
rect 27522 14590 27636 14642
rect 27468 14588 27636 14590
rect 27468 14578 27524 14588
rect 27132 13916 27300 13972
rect 27132 13746 27188 13758
rect 27132 13694 27134 13746
rect 27186 13694 27188 13746
rect 27132 13636 27188 13694
rect 27132 13570 27188 13580
rect 26012 13074 26404 13076
rect 26012 13022 26014 13074
rect 26066 13022 26404 13074
rect 26012 13020 26404 13022
rect 26012 13010 26068 13020
rect 26348 12404 26404 13020
rect 26908 12404 26964 12414
rect 26404 12402 26964 12404
rect 26404 12350 26910 12402
rect 26962 12350 26964 12402
rect 26404 12348 26964 12350
rect 26348 12310 26404 12348
rect 26908 12338 26964 12348
rect 26236 12180 26292 12190
rect 26236 11844 26292 12124
rect 26572 12180 26628 12190
rect 26572 12178 26740 12180
rect 26572 12126 26574 12178
rect 26626 12126 26740 12178
rect 26572 12124 26740 12126
rect 26572 12114 26628 12124
rect 26236 11778 26292 11788
rect 25900 11564 26180 11620
rect 25676 11506 25844 11508
rect 25676 11454 25678 11506
rect 25730 11454 25844 11506
rect 25676 11452 25844 11454
rect 25676 11442 25732 11452
rect 25788 10612 25844 11452
rect 25900 11396 25956 11406
rect 25900 11394 26068 11396
rect 25900 11342 25902 11394
rect 25954 11342 26068 11394
rect 25900 11340 26068 11342
rect 25900 11330 25956 11340
rect 26012 10836 26068 11340
rect 25788 10610 25956 10612
rect 25788 10558 25790 10610
rect 25842 10558 25956 10610
rect 25788 10556 25956 10558
rect 25788 10546 25844 10556
rect 25004 9874 25060 9884
rect 25564 9874 25620 9884
rect 25900 9938 25956 10556
rect 26012 10500 26068 10780
rect 26124 10612 26180 11564
rect 26684 11396 26740 12124
rect 27132 11508 27188 11518
rect 27020 11506 27188 11508
rect 27020 11454 27134 11506
rect 27186 11454 27188 11506
rect 27020 11452 27188 11454
rect 26908 11396 26964 11406
rect 26684 11394 26964 11396
rect 26684 11342 26910 11394
rect 26962 11342 26964 11394
rect 26684 11340 26964 11342
rect 26908 11330 26964 11340
rect 26236 11172 26292 11182
rect 26236 11170 26852 11172
rect 26236 11118 26238 11170
rect 26290 11118 26852 11170
rect 26236 11116 26852 11118
rect 26236 11106 26292 11116
rect 26796 10834 26852 11116
rect 26796 10782 26798 10834
rect 26850 10782 26852 10834
rect 26796 10770 26852 10782
rect 26908 10836 26964 10846
rect 27020 10836 27076 11452
rect 27132 11442 27188 11452
rect 26908 10834 27076 10836
rect 26908 10782 26910 10834
rect 26962 10782 27076 10834
rect 26908 10780 27076 10782
rect 27244 10836 27300 13916
rect 27580 12516 27636 14588
rect 27916 14530 27972 15484
rect 28252 15148 28308 24780
rect 28812 24834 28868 24846
rect 28812 24782 28814 24834
rect 28866 24782 28868 24834
rect 28588 24612 28644 24622
rect 28476 23156 28532 23166
rect 28476 23062 28532 23100
rect 28364 21474 28420 21486
rect 28364 21422 28366 21474
rect 28418 21422 28420 21474
rect 28364 20692 28420 21422
rect 28588 21364 28644 24556
rect 28812 23380 28868 24782
rect 28812 22484 28868 23324
rect 28812 22418 28868 22428
rect 28588 21308 28756 21364
rect 28588 21140 28644 21150
rect 28588 20914 28644 21084
rect 28588 20862 28590 20914
rect 28642 20862 28644 20914
rect 28588 20850 28644 20862
rect 28588 20692 28644 20702
rect 28364 20636 28588 20692
rect 28588 20130 28644 20636
rect 28588 20078 28590 20130
rect 28642 20078 28644 20130
rect 28588 20066 28644 20078
rect 28700 19348 28756 21308
rect 28700 19282 28756 19292
rect 28812 18452 28868 18462
rect 28364 18396 28812 18452
rect 28364 17778 28420 18396
rect 28812 18358 28868 18396
rect 28364 17726 28366 17778
rect 28418 17726 28420 17778
rect 28364 17714 28420 17726
rect 28588 17108 28644 17118
rect 28588 17014 28644 17052
rect 28252 15092 28420 15148
rect 27916 14478 27918 14530
rect 27970 14478 27972 14530
rect 27916 14466 27972 14478
rect 27580 12460 28196 12516
rect 27580 12402 27636 12460
rect 27580 12350 27582 12402
rect 27634 12350 27636 12402
rect 27580 12338 27636 12350
rect 27804 12292 27860 12302
rect 27804 12198 27860 12236
rect 27468 12180 27524 12190
rect 27468 11060 27524 12124
rect 27580 11396 27636 11406
rect 27580 11394 27972 11396
rect 27580 11342 27582 11394
rect 27634 11342 27972 11394
rect 27580 11340 27972 11342
rect 27580 11330 27636 11340
rect 27804 11170 27860 11182
rect 27804 11118 27806 11170
rect 27858 11118 27860 11170
rect 27468 11004 27748 11060
rect 27244 10780 27636 10836
rect 26908 10770 26964 10780
rect 27020 10612 27076 10622
rect 26124 10556 26404 10612
rect 26012 10498 26180 10500
rect 26012 10446 26014 10498
rect 26066 10446 26180 10498
rect 26012 10444 26180 10446
rect 26012 10434 26068 10444
rect 26124 10050 26180 10444
rect 26124 9998 26126 10050
rect 26178 9998 26180 10050
rect 26124 9986 26180 9998
rect 25900 9886 25902 9938
rect 25954 9886 25956 9938
rect 25900 9874 25956 9886
rect 26236 7812 26292 7822
rect 25228 7474 25284 7486
rect 25228 7422 25230 7474
rect 25282 7422 25284 7474
rect 25228 6916 25284 7422
rect 25788 7476 25844 7486
rect 25788 7382 25844 7420
rect 25228 6850 25284 6860
rect 25676 7362 25732 7374
rect 25676 7310 25678 7362
rect 25730 7310 25732 7362
rect 25676 5908 25732 7310
rect 26236 6018 26292 7756
rect 26348 7588 26404 10556
rect 27020 10610 27188 10612
rect 27020 10558 27022 10610
rect 27074 10558 27188 10610
rect 27020 10556 27188 10558
rect 27020 10546 27076 10556
rect 26460 10500 26516 10510
rect 26460 10498 26852 10500
rect 26460 10446 26462 10498
rect 26514 10446 26852 10498
rect 26460 10444 26852 10446
rect 26460 10434 26516 10444
rect 26460 10164 26516 10174
rect 26460 10050 26516 10108
rect 26460 9998 26462 10050
rect 26514 9998 26516 10050
rect 26460 9986 26516 9998
rect 26796 8428 26852 10444
rect 27020 10388 27076 10398
rect 26908 10332 27020 10388
rect 26908 9826 26964 10332
rect 27020 10322 27076 10332
rect 26908 9774 26910 9826
rect 26962 9774 26964 9826
rect 26908 9762 26964 9774
rect 27020 9716 27076 9726
rect 27020 9622 27076 9660
rect 26796 8372 27076 8428
rect 26908 7924 26964 7934
rect 26348 7586 26628 7588
rect 26348 7534 26350 7586
rect 26402 7534 26628 7586
rect 26348 7532 26628 7534
rect 26348 7522 26404 7532
rect 26572 6802 26628 7532
rect 26908 7474 26964 7868
rect 26908 7422 26910 7474
rect 26962 7422 26964 7474
rect 26908 6916 26964 7422
rect 26908 6850 26964 6860
rect 26572 6750 26574 6802
rect 26626 6750 26628 6802
rect 26572 6132 26628 6750
rect 26572 6066 26628 6076
rect 26236 5966 26238 6018
rect 26290 5966 26292 6018
rect 26236 5954 26292 5966
rect 25676 5906 26180 5908
rect 25676 5854 25678 5906
rect 25730 5854 26180 5906
rect 25676 5852 26180 5854
rect 25676 5842 25732 5852
rect 25340 5794 25396 5806
rect 25340 5742 25342 5794
rect 25394 5742 25396 5794
rect 25004 5348 25060 5358
rect 25004 5254 25060 5292
rect 25340 5236 25396 5742
rect 25340 5012 25396 5180
rect 26012 5236 26068 5246
rect 26012 5142 26068 5180
rect 26124 5012 26180 5852
rect 25340 4226 25396 4956
rect 25900 5010 26180 5012
rect 25900 4958 26126 5010
rect 26178 4958 26180 5010
rect 25900 4956 26180 4958
rect 25900 4450 25956 4956
rect 26124 4946 26180 4956
rect 25900 4398 25902 4450
rect 25954 4398 25956 4450
rect 25900 4340 25956 4398
rect 25900 4274 25956 4284
rect 27020 4338 27076 8372
rect 27132 7812 27188 10556
rect 27356 10610 27412 10622
rect 27356 10558 27358 10610
rect 27410 10558 27412 10610
rect 27356 10164 27412 10558
rect 27356 10098 27412 10108
rect 27580 9716 27636 10780
rect 27692 10388 27748 11004
rect 27692 10322 27748 10332
rect 27580 9622 27636 9660
rect 27244 9602 27300 9614
rect 27244 9550 27246 9602
rect 27298 9550 27300 9602
rect 27244 8428 27300 9550
rect 27804 8428 27860 11118
rect 27916 10500 27972 11340
rect 28028 11284 28084 12460
rect 28140 12402 28196 12460
rect 28140 12350 28142 12402
rect 28194 12350 28196 12402
rect 28140 12338 28196 12350
rect 28252 12404 28308 12414
rect 28140 11396 28196 11406
rect 28252 11396 28308 12348
rect 28364 12180 28420 15092
rect 28924 14644 28980 26124
rect 29036 25508 29092 26238
rect 29148 26292 29204 26302
rect 29148 26198 29204 26236
rect 29036 25284 29092 25452
rect 29260 25284 29316 25294
rect 29036 25282 29316 25284
rect 29036 25230 29262 25282
rect 29314 25230 29316 25282
rect 29036 25228 29316 25230
rect 29260 25218 29316 25228
rect 29036 24892 29316 24948
rect 29036 21698 29092 24892
rect 29260 24836 29316 24892
rect 29484 24836 29540 29372
rect 29708 29426 29764 29438
rect 29708 29374 29710 29426
rect 29762 29374 29764 29426
rect 29260 24780 29540 24836
rect 29596 29316 29652 29326
rect 29148 24724 29204 24734
rect 29148 24050 29204 24668
rect 29484 24610 29540 24622
rect 29484 24558 29486 24610
rect 29538 24558 29540 24610
rect 29484 24500 29540 24558
rect 29148 23998 29150 24050
rect 29202 23998 29204 24050
rect 29148 23986 29204 23998
rect 29260 24444 29540 24500
rect 29148 23156 29204 23166
rect 29260 23156 29316 24444
rect 29596 24388 29652 29260
rect 29708 27972 29764 29374
rect 30156 29316 30212 32620
rect 30156 29250 30212 29260
rect 29708 27906 29764 27916
rect 30156 27858 30212 27870
rect 30156 27806 30158 27858
rect 30210 27806 30212 27858
rect 29204 23100 29316 23156
rect 29372 24332 29652 24388
rect 29708 27748 29764 27758
rect 29148 23062 29204 23100
rect 29372 22708 29428 24332
rect 29708 24276 29764 27692
rect 30156 27636 30212 27806
rect 30268 27636 30324 27646
rect 30156 27580 30268 27636
rect 30268 27570 30324 27580
rect 30268 26962 30324 26974
rect 30268 26910 30270 26962
rect 30322 26910 30324 26962
rect 30268 26908 30324 26910
rect 29708 24210 29764 24220
rect 29820 26852 30324 26908
rect 30380 26908 30436 33068
rect 30716 32674 30772 32686
rect 30716 32622 30718 32674
rect 30770 32622 30772 32674
rect 30716 31780 30772 32622
rect 30716 31686 30772 31724
rect 30828 30996 30884 31006
rect 30828 30902 30884 30940
rect 30828 28420 30884 28430
rect 30604 27748 30660 27758
rect 30604 27654 30660 27692
rect 30828 27074 30884 28364
rect 30828 27022 30830 27074
rect 30882 27022 30884 27074
rect 30828 27010 30884 27022
rect 30828 26908 30884 26918
rect 30380 26852 30772 26908
rect 29596 24052 29652 24062
rect 29596 24050 29764 24052
rect 29596 23998 29598 24050
rect 29650 23998 29764 24050
rect 29596 23996 29764 23998
rect 29596 23986 29652 23996
rect 29596 23716 29652 23726
rect 29596 23548 29652 23660
rect 29372 22642 29428 22652
rect 29484 23492 29652 23548
rect 29260 22484 29316 22494
rect 29260 22390 29316 22428
rect 29036 21646 29038 21698
rect 29090 21646 29092 21698
rect 29036 21634 29092 21646
rect 29036 19908 29092 19918
rect 29036 19814 29092 19852
rect 28924 14578 28980 14588
rect 29036 18562 29092 18574
rect 29036 18510 29038 18562
rect 29090 18510 29092 18562
rect 29036 14532 29092 18510
rect 29372 17780 29428 17790
rect 29372 16884 29428 17724
rect 29372 16210 29428 16828
rect 29372 16158 29374 16210
rect 29426 16158 29428 16210
rect 29372 16146 29428 16158
rect 29484 15148 29540 23492
rect 29708 23268 29764 23996
rect 29820 23938 29876 26852
rect 29820 23886 29822 23938
rect 29874 23886 29876 23938
rect 29820 23378 29876 23886
rect 29820 23326 29822 23378
rect 29874 23326 29876 23378
rect 29820 23314 29876 23326
rect 29932 24610 29988 24622
rect 29932 24558 29934 24610
rect 29986 24558 29988 24610
rect 29932 23380 29988 24558
rect 29932 23314 29988 23324
rect 29596 23266 29764 23268
rect 29596 23214 29710 23266
rect 29762 23214 29764 23266
rect 29596 23212 29764 23214
rect 29596 21026 29652 23212
rect 29708 23202 29764 23212
rect 30044 23156 30100 23166
rect 30044 23154 30660 23156
rect 30044 23102 30046 23154
rect 30098 23102 30660 23154
rect 30044 23100 30660 23102
rect 30044 23090 30100 23100
rect 30492 21700 30548 21710
rect 30380 21698 30548 21700
rect 30380 21646 30494 21698
rect 30546 21646 30548 21698
rect 30380 21644 30548 21646
rect 29708 21588 29764 21598
rect 29708 21494 29764 21532
rect 30268 21588 30324 21598
rect 30268 21494 30324 21532
rect 29932 21476 29988 21486
rect 29596 20974 29598 21026
rect 29650 20974 29652 21026
rect 29596 20962 29652 20974
rect 29820 21474 29988 21476
rect 29820 21422 29934 21474
rect 29986 21422 29988 21474
rect 29820 21420 29988 21422
rect 29820 16996 29876 21420
rect 29932 21410 29988 21420
rect 30380 21140 30436 21644
rect 30492 21634 30548 21644
rect 30604 21698 30660 23100
rect 30604 21646 30606 21698
rect 30658 21646 30660 21698
rect 30604 21634 30660 21646
rect 29932 21084 30436 21140
rect 29932 20130 29988 21084
rect 30716 21028 30772 26852
rect 30828 26516 30884 26852
rect 30940 26740 30996 33292
rect 31052 32564 31108 32574
rect 31052 32470 31108 32508
rect 30940 26674 30996 26684
rect 31052 27186 31108 27198
rect 31052 27134 31054 27186
rect 31106 27134 31108 27186
rect 30940 26516 30996 26526
rect 30828 26514 30996 26516
rect 30828 26462 30942 26514
rect 30994 26462 30996 26514
rect 30828 26460 30996 26462
rect 30940 26450 30996 26460
rect 31052 26514 31108 27134
rect 31052 26462 31054 26514
rect 31106 26462 31108 26514
rect 31052 26450 31108 26462
rect 31164 26628 31220 26638
rect 31164 26292 31220 26572
rect 31276 26404 31332 35532
rect 31388 35522 31444 35532
rect 31500 31332 31556 36540
rect 31836 35698 31892 35710
rect 31836 35646 31838 35698
rect 31890 35646 31892 35698
rect 31836 35140 31892 35646
rect 31836 35074 31892 35084
rect 32060 35252 32116 35262
rect 31836 34916 31892 34926
rect 31836 34822 31892 34860
rect 32060 34914 32116 35196
rect 32060 34862 32062 34914
rect 32114 34862 32116 34914
rect 32060 34850 32116 34862
rect 32172 35138 32228 35150
rect 32172 35086 32174 35138
rect 32226 35086 32228 35138
rect 32060 33124 32116 33134
rect 32060 32564 32116 33068
rect 32060 32470 32116 32508
rect 31948 32450 32004 32462
rect 31948 32398 31950 32450
rect 32002 32398 32004 32450
rect 31724 32340 31780 32350
rect 31612 32338 31780 32340
rect 31612 32286 31726 32338
rect 31778 32286 31780 32338
rect 31612 32284 31780 32286
rect 31612 31780 31668 32284
rect 31724 32274 31780 32284
rect 31724 31892 31780 31902
rect 31724 31798 31780 31836
rect 31612 31714 31668 31724
rect 31500 31266 31556 31276
rect 31948 31220 32004 32398
rect 31948 31154 32004 31164
rect 32060 31106 32116 31118
rect 32060 31054 32062 31106
rect 32114 31054 32116 31106
rect 31388 30996 31444 31006
rect 31444 30940 31668 30996
rect 31388 30930 31444 30940
rect 31612 29426 31668 30940
rect 31612 29374 31614 29426
rect 31666 29374 31668 29426
rect 31612 28532 31668 29374
rect 31836 30994 31892 31006
rect 31836 30942 31838 30994
rect 31890 30942 31892 30994
rect 31836 29428 31892 30942
rect 31948 30884 32004 30894
rect 31948 30210 32004 30828
rect 32060 30772 32116 31054
rect 32060 30706 32116 30716
rect 31948 30158 31950 30210
rect 32002 30158 32004 30210
rect 31948 30146 32004 30158
rect 32060 30098 32116 30110
rect 32060 30046 32062 30098
rect 32114 30046 32116 30098
rect 31948 29428 32004 29438
rect 31836 29372 31948 29428
rect 31948 29334 32004 29372
rect 31612 28466 31668 28476
rect 31948 28532 32004 28542
rect 31276 26338 31332 26348
rect 31388 27748 31444 27758
rect 31388 26404 31444 27692
rect 31612 27636 31668 27646
rect 31500 27580 31612 27636
rect 31500 26964 31556 27580
rect 31612 27570 31668 27580
rect 31948 27186 32004 28476
rect 32060 28420 32116 30046
rect 32060 28354 32116 28364
rect 31948 27134 31950 27186
rect 32002 27134 32004 27186
rect 31948 27122 32004 27134
rect 32060 28084 32116 28094
rect 31612 27076 31668 27086
rect 32060 27076 32116 28028
rect 31612 27074 31892 27076
rect 31612 27022 31614 27074
rect 31666 27022 31892 27074
rect 31612 27020 31892 27022
rect 31612 27010 31668 27020
rect 31500 26852 31668 26908
rect 31612 26514 31668 26852
rect 31612 26462 31614 26514
rect 31666 26462 31668 26514
rect 31612 26450 31668 26462
rect 31724 26852 31780 26862
rect 31500 26404 31556 26414
rect 31388 26402 31556 26404
rect 31388 26350 31502 26402
rect 31554 26350 31556 26402
rect 31388 26348 31556 26350
rect 31052 26236 31220 26292
rect 30940 23716 30996 23726
rect 31052 23716 31108 26236
rect 31388 26180 31444 26348
rect 31500 26338 31556 26348
rect 31164 26124 31444 26180
rect 31612 26292 31668 26302
rect 31164 26066 31220 26124
rect 31164 26014 31166 26066
rect 31218 26014 31220 26066
rect 31164 25956 31220 26014
rect 31164 25900 31332 25956
rect 31164 23938 31220 23950
rect 31164 23886 31166 23938
rect 31218 23886 31220 23938
rect 31164 23716 31220 23886
rect 30940 23714 31220 23716
rect 30940 23662 30942 23714
rect 30994 23662 31220 23714
rect 30940 23660 31220 23662
rect 30940 23650 30996 23660
rect 30716 20972 30884 21028
rect 30044 20914 30100 20926
rect 30044 20862 30046 20914
rect 30098 20862 30100 20914
rect 30044 20804 30100 20862
rect 30044 20738 30100 20748
rect 30156 20802 30212 20814
rect 30156 20750 30158 20802
rect 30210 20750 30212 20802
rect 29932 20078 29934 20130
rect 29986 20078 29988 20130
rect 29932 20066 29988 20078
rect 30156 20242 30212 20750
rect 30156 20190 30158 20242
rect 30210 20190 30212 20242
rect 30156 20020 30212 20190
rect 30716 20804 30772 20814
rect 30156 19954 30212 19964
rect 30268 20020 30324 20030
rect 30604 20020 30660 20030
rect 30268 20018 30660 20020
rect 30268 19966 30270 20018
rect 30322 19966 30606 20018
rect 30658 19966 30660 20018
rect 30268 19964 30660 19966
rect 30268 19954 30324 19964
rect 30604 19954 30660 19964
rect 30716 19908 30772 20748
rect 30828 20132 30884 20972
rect 30828 20066 30884 20076
rect 30940 19908 30996 19918
rect 30716 19906 30884 19908
rect 30716 19854 30718 19906
rect 30770 19854 30884 19906
rect 30716 19852 30884 19854
rect 30716 19842 30772 19852
rect 29932 18340 29988 18350
rect 29988 18284 30324 18340
rect 29932 18246 29988 18284
rect 30268 17666 30324 18284
rect 30268 17614 30270 17666
rect 30322 17614 30324 17666
rect 30268 17602 30324 17614
rect 29932 17444 29988 17454
rect 29932 17350 29988 17388
rect 30380 17442 30436 17454
rect 30380 17390 30382 17442
rect 30434 17390 30436 17442
rect 29596 16940 29876 16996
rect 29596 15876 29652 16940
rect 29932 16884 29988 16894
rect 30380 16884 30436 17390
rect 30492 17444 30548 17454
rect 30492 17350 30548 17388
rect 30716 17442 30772 17454
rect 30716 17390 30718 17442
rect 30770 17390 30772 17442
rect 30604 16884 30660 16894
rect 30380 16882 30660 16884
rect 30380 16830 30606 16882
rect 30658 16830 30660 16882
rect 30380 16828 30660 16830
rect 29820 16772 29876 16782
rect 29708 16770 29876 16772
rect 29708 16718 29822 16770
rect 29874 16718 29876 16770
rect 29708 16716 29876 16718
rect 29708 16212 29764 16716
rect 29820 16706 29876 16716
rect 29708 16098 29764 16156
rect 29708 16046 29710 16098
rect 29762 16046 29764 16098
rect 29708 16034 29764 16046
rect 29820 16100 29876 16110
rect 29820 16006 29876 16044
rect 29932 16098 29988 16828
rect 30604 16818 30660 16828
rect 29932 16046 29934 16098
rect 29986 16046 29988 16098
rect 29932 16034 29988 16046
rect 30268 16658 30324 16670
rect 30268 16606 30270 16658
rect 30322 16606 30324 16658
rect 29596 15820 30100 15876
rect 29820 15652 29876 15662
rect 29484 15092 29652 15148
rect 29260 14644 29316 14654
rect 29148 14532 29204 14542
rect 29036 14530 29204 14532
rect 29036 14478 29150 14530
rect 29202 14478 29204 14530
rect 29036 14476 29204 14478
rect 29148 14084 29204 14476
rect 29148 14018 29204 14028
rect 28476 12180 28532 12190
rect 28364 12124 28476 12180
rect 28476 12114 28532 12124
rect 28140 11394 28252 11396
rect 28140 11342 28142 11394
rect 28194 11342 28252 11394
rect 28140 11340 28252 11342
rect 28140 11330 28196 11340
rect 28252 11302 28308 11340
rect 29148 11508 29204 11518
rect 29148 11394 29204 11452
rect 29148 11342 29150 11394
rect 29202 11342 29204 11394
rect 29148 11330 29204 11342
rect 28028 11190 28084 11228
rect 28588 11284 28644 11294
rect 28588 11190 28644 11228
rect 29260 11284 29316 14588
rect 29596 13748 29652 15036
rect 29708 14644 29764 14654
rect 29708 14550 29764 14588
rect 29708 13748 29764 13758
rect 29596 13746 29764 13748
rect 29596 13694 29710 13746
rect 29762 13694 29764 13746
rect 29596 13692 29764 13694
rect 29708 13682 29764 13692
rect 29372 13522 29428 13534
rect 29372 13470 29374 13522
rect 29426 13470 29428 13522
rect 29372 13074 29428 13470
rect 29372 13022 29374 13074
rect 29426 13022 29428 13074
rect 29372 13010 29428 13022
rect 29708 12964 29764 12974
rect 29820 12964 29876 15596
rect 29708 12962 29876 12964
rect 29708 12910 29710 12962
rect 29762 12910 29876 12962
rect 29708 12908 29876 12910
rect 29932 15428 29988 15438
rect 29708 12898 29764 12908
rect 29820 11508 29876 11518
rect 29932 11508 29988 15372
rect 29876 11452 29988 11508
rect 29820 11414 29876 11452
rect 29260 11190 29316 11228
rect 29484 11170 29540 11182
rect 29484 11118 29486 11170
rect 29538 11118 29540 11170
rect 28476 10722 28532 10734
rect 28476 10670 28478 10722
rect 28530 10670 28532 10722
rect 28140 10500 28196 10510
rect 27916 10498 28196 10500
rect 27916 10446 28142 10498
rect 28194 10446 28196 10498
rect 27916 10444 28196 10446
rect 28140 10434 28196 10444
rect 28476 9044 28532 10670
rect 29484 10052 29540 11118
rect 30044 10834 30100 15820
rect 30156 15092 30212 15102
rect 30156 14642 30212 15036
rect 30156 14590 30158 14642
rect 30210 14590 30212 14642
rect 30156 14578 30212 14590
rect 30268 14084 30324 16606
rect 30716 16212 30772 17390
rect 30716 16146 30772 16156
rect 30380 16100 30436 16110
rect 30436 16044 30660 16100
rect 30380 16006 30436 16044
rect 30604 15538 30660 16044
rect 30604 15486 30606 15538
rect 30658 15486 30660 15538
rect 30604 15474 30660 15486
rect 30716 15986 30772 15998
rect 30716 15934 30718 15986
rect 30770 15934 30772 15986
rect 30492 15092 30548 15102
rect 30492 14756 30548 15036
rect 30492 14530 30548 14700
rect 30492 14478 30494 14530
rect 30546 14478 30548 14530
rect 30492 14466 30548 14478
rect 30604 14644 30660 14654
rect 30604 14418 30660 14588
rect 30604 14366 30606 14418
rect 30658 14366 30660 14418
rect 30604 14354 30660 14366
rect 30156 14028 30660 14084
rect 30156 13746 30212 14028
rect 30492 13860 30548 13870
rect 30492 13766 30548 13804
rect 30156 13694 30158 13746
rect 30210 13694 30212 13746
rect 30156 13682 30212 13694
rect 30604 13074 30660 14028
rect 30604 13022 30606 13074
rect 30658 13022 30660 13074
rect 30604 13010 30660 13022
rect 30044 10782 30046 10834
rect 30098 10782 30100 10834
rect 30044 10770 30100 10782
rect 30156 12850 30212 12862
rect 30156 12798 30158 12850
rect 30210 12798 30212 12850
rect 29484 9986 29540 9996
rect 29596 10610 29652 10622
rect 29596 10558 29598 10610
rect 29650 10558 29652 10610
rect 29484 9604 29540 9614
rect 29596 9604 29652 10558
rect 29484 9602 29652 9604
rect 29484 9550 29486 9602
rect 29538 9550 29652 9602
rect 29484 9548 29652 9550
rect 29820 9826 29876 9838
rect 29820 9774 29822 9826
rect 29874 9774 29876 9826
rect 29484 9538 29540 9548
rect 28476 8978 28532 8988
rect 27244 8372 27524 8428
rect 27804 8372 28196 8428
rect 27356 8260 27412 8270
rect 27132 7746 27188 7756
rect 27244 8258 27412 8260
rect 27244 8206 27358 8258
rect 27410 8206 27412 8258
rect 27244 8204 27412 8206
rect 27244 6914 27300 8204
rect 27356 8194 27412 8204
rect 27468 7924 27524 8372
rect 27468 7858 27524 7868
rect 27804 8034 27860 8046
rect 27804 7982 27806 8034
rect 27858 7982 27860 8034
rect 27804 7812 27860 7982
rect 27916 8036 27972 8046
rect 27916 7942 27972 7980
rect 28028 8034 28084 8046
rect 28028 7982 28030 8034
rect 28082 7982 28084 8034
rect 27804 7746 27860 7756
rect 28028 7700 28084 7982
rect 27356 7644 27636 7700
rect 27356 7474 27412 7644
rect 27580 7588 27636 7644
rect 28028 7634 28084 7644
rect 27580 7532 27972 7588
rect 27356 7422 27358 7474
rect 27410 7422 27412 7474
rect 27356 7410 27412 7422
rect 27916 7476 27972 7532
rect 28140 7476 28196 8372
rect 28252 7924 28308 7934
rect 28308 7868 28420 7924
rect 28252 7858 28308 7868
rect 27916 7474 28196 7476
rect 27916 7422 28142 7474
rect 28194 7422 28196 7474
rect 27916 7420 28196 7422
rect 27804 7364 27860 7374
rect 27692 7362 27860 7364
rect 27692 7310 27806 7362
rect 27858 7310 27860 7362
rect 27692 7308 27860 7310
rect 27244 6862 27246 6914
rect 27298 6862 27300 6914
rect 27244 6850 27300 6862
rect 27356 6916 27412 6926
rect 27580 6916 27636 6926
rect 27412 6914 27636 6916
rect 27412 6862 27582 6914
rect 27634 6862 27636 6914
rect 27412 6860 27636 6862
rect 27356 6850 27412 6860
rect 27580 6850 27636 6860
rect 27580 5124 27636 5134
rect 27692 5124 27748 7308
rect 27804 7298 27860 7308
rect 27804 6804 27860 6814
rect 27916 6804 27972 7420
rect 28140 7410 28196 7420
rect 28364 7474 28420 7868
rect 28700 7700 28756 7710
rect 28700 7606 28756 7644
rect 28364 7422 28366 7474
rect 28418 7422 28420 7474
rect 28364 7410 28420 7422
rect 29820 7140 29876 9774
rect 30156 8428 30212 12798
rect 30716 12180 30772 15934
rect 30828 15148 30884 19852
rect 30940 17892 30996 19852
rect 30940 17826 30996 17836
rect 30828 15092 30996 15148
rect 30828 14306 30884 14318
rect 30828 14254 30830 14306
rect 30882 14254 30884 14306
rect 30828 12964 30884 14254
rect 30828 12870 30884 12908
rect 30604 12124 30772 12180
rect 30268 11284 30324 11294
rect 30268 11190 30324 11228
rect 29820 7074 29876 7084
rect 29932 8372 30212 8428
rect 27804 6802 27972 6804
rect 27804 6750 27806 6802
rect 27858 6750 27972 6802
rect 27804 6748 27972 6750
rect 27804 6738 27860 6748
rect 29708 6692 29764 6702
rect 29260 6690 29764 6692
rect 29260 6638 29710 6690
rect 29762 6638 29764 6690
rect 29260 6636 29764 6638
rect 28700 6018 28756 6030
rect 28700 5966 28702 6018
rect 28754 5966 28756 6018
rect 28700 5348 28756 5966
rect 29260 5906 29316 6636
rect 29708 6626 29764 6636
rect 29260 5854 29262 5906
rect 29314 5854 29316 5906
rect 29260 5842 29316 5854
rect 29596 6466 29652 6478
rect 29596 6414 29598 6466
rect 29650 6414 29652 6466
rect 28700 5282 28756 5292
rect 29484 5236 29540 5246
rect 29596 5236 29652 6414
rect 29820 6466 29876 6478
rect 29820 6414 29822 6466
rect 29874 6414 29876 6466
rect 29820 6356 29876 6414
rect 29820 6290 29876 6300
rect 29932 5906 29988 8372
rect 30268 7140 30324 7150
rect 29932 5854 29934 5906
rect 29986 5854 29988 5906
rect 29932 5842 29988 5854
rect 30156 6690 30212 6702
rect 30156 6638 30158 6690
rect 30210 6638 30212 6690
rect 29484 5234 29652 5236
rect 29484 5182 29486 5234
rect 29538 5182 29652 5234
rect 29484 5180 29652 5182
rect 29484 5170 29540 5180
rect 27580 5122 27748 5124
rect 27580 5070 27582 5122
rect 27634 5070 27748 5122
rect 27580 5068 27748 5070
rect 29372 5124 29428 5134
rect 27580 5058 27636 5068
rect 28028 5010 28084 5022
rect 28028 4958 28030 5010
rect 28082 4958 28084 5010
rect 28028 4900 28084 4958
rect 29372 5010 29428 5068
rect 30044 5124 30100 5134
rect 29372 4958 29374 5010
rect 29426 4958 29428 5010
rect 29372 4946 29428 4958
rect 29596 5012 29652 5022
rect 29596 5010 29988 5012
rect 29596 4958 29598 5010
rect 29650 4958 29988 5010
rect 29596 4956 29988 4958
rect 29596 4946 29652 4956
rect 28028 4834 28084 4844
rect 29932 4452 29988 4956
rect 30044 4562 30100 5068
rect 30044 4510 30046 4562
rect 30098 4510 30100 4562
rect 30044 4498 30100 4510
rect 29932 4358 29988 4396
rect 27020 4286 27022 4338
rect 27074 4286 27076 4338
rect 27020 4274 27076 4286
rect 27468 4340 27524 4350
rect 27468 4246 27524 4284
rect 25340 4174 25342 4226
rect 25394 4174 25396 4226
rect 25340 4162 25396 4174
rect 30044 4116 30100 4126
rect 30156 4116 30212 6638
rect 30268 6130 30324 7084
rect 30268 6078 30270 6130
rect 30322 6078 30324 6130
rect 30268 6066 30324 6078
rect 30380 6356 30436 6366
rect 30380 5010 30436 6300
rect 30604 5124 30660 12124
rect 30716 10052 30772 10062
rect 30716 9714 30772 9996
rect 30716 9662 30718 9714
rect 30770 9662 30772 9714
rect 30716 9650 30772 9662
rect 30940 8428 30996 15092
rect 31052 14644 31108 23660
rect 31276 21026 31332 25900
rect 31500 24724 31556 24734
rect 31612 24724 31668 26236
rect 31500 24722 31668 24724
rect 31500 24670 31502 24722
rect 31554 24670 31668 24722
rect 31500 24668 31668 24670
rect 31500 24658 31556 24668
rect 31612 23940 31668 24668
rect 31612 23874 31668 23884
rect 31724 21924 31780 26796
rect 31836 26514 31892 27020
rect 32060 27010 32116 27020
rect 31836 26462 31838 26514
rect 31890 26462 31892 26514
rect 31836 26450 31892 26462
rect 32172 25844 32228 35086
rect 32284 35026 32340 36988
rect 32396 36978 32452 36988
rect 32508 35140 32564 40124
rect 32620 39620 32676 39630
rect 32620 39526 32676 39564
rect 32620 37044 32676 37054
rect 32620 36482 32676 36988
rect 32620 36430 32622 36482
rect 32674 36430 32676 36482
rect 32620 36418 32676 36430
rect 32732 35700 32788 40348
rect 32732 35634 32788 35644
rect 32284 34974 32286 35026
rect 32338 34974 32340 35026
rect 32284 34962 32340 34974
rect 32396 35084 32564 35140
rect 32396 26908 32452 35084
rect 32620 30212 32676 30222
rect 32508 30210 32676 30212
rect 32508 30158 32622 30210
rect 32674 30158 32676 30210
rect 32508 30156 32676 30158
rect 32508 29538 32564 30156
rect 32620 30146 32676 30156
rect 32508 29486 32510 29538
rect 32562 29486 32564 29538
rect 32508 29474 32564 29486
rect 32732 29428 32788 29438
rect 32620 28532 32676 28542
rect 32620 28438 32676 28476
rect 32732 28418 32788 29372
rect 32732 28366 32734 28418
rect 32786 28366 32788 28418
rect 32732 27300 32788 28366
rect 32844 27412 32900 40796
rect 33068 40514 33124 40908
rect 33068 40462 33070 40514
rect 33122 40462 33124 40514
rect 33068 40450 33124 40462
rect 33180 40628 33236 41804
rect 33180 40514 33236 40572
rect 33180 40462 33182 40514
rect 33234 40462 33236 40514
rect 33180 40404 33236 40462
rect 33180 40338 33236 40348
rect 33180 40178 33236 40190
rect 33180 40126 33182 40178
rect 33234 40126 33236 40178
rect 33180 39618 33236 40126
rect 33180 39566 33182 39618
rect 33234 39566 33236 39618
rect 33180 39554 33236 39566
rect 32956 36596 33012 36606
rect 32956 31892 33012 36540
rect 33068 36370 33124 36382
rect 33068 36318 33070 36370
rect 33122 36318 33124 36370
rect 33068 34916 33124 36318
rect 33292 35812 33348 41916
rect 33404 41074 33460 41086
rect 33404 41022 33406 41074
rect 33458 41022 33460 41074
rect 33404 39844 33460 41022
rect 33516 40852 33572 42364
rect 33740 42082 33796 42812
rect 34412 42802 34468 42812
rect 33964 42644 34020 42654
rect 34020 42588 34356 42644
rect 33964 42550 34020 42588
rect 33740 42030 33742 42082
rect 33794 42030 33796 42082
rect 33740 41412 33796 42030
rect 33852 42084 33908 42094
rect 33852 41990 33908 42028
rect 34300 42082 34356 42588
rect 34300 42030 34302 42082
rect 34354 42030 34356 42082
rect 34076 41972 34132 41982
rect 34076 41970 34244 41972
rect 34076 41918 34078 41970
rect 34130 41918 34244 41970
rect 34076 41916 34244 41918
rect 34076 41906 34132 41916
rect 34188 41412 34244 41916
rect 34300 41860 34356 42030
rect 34412 42084 34468 42094
rect 34412 41990 34468 42028
rect 35420 41972 35476 41982
rect 35420 41878 35476 41916
rect 35644 41860 35700 41870
rect 34300 41794 34356 41804
rect 35532 41858 35700 41860
rect 35532 41806 35646 41858
rect 35698 41806 35700 41858
rect 35532 41804 35700 41806
rect 34412 41748 34468 41758
rect 34412 41654 34468 41692
rect 35532 41748 35588 41804
rect 35644 41794 35700 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35084 41412 35140 41422
rect 33740 41356 34132 41412
rect 34188 41356 34468 41412
rect 33964 41188 34020 41198
rect 33964 41094 34020 41132
rect 33516 40786 33572 40796
rect 33740 41076 33796 41086
rect 33404 39788 33684 39844
rect 33628 39730 33684 39788
rect 33628 39678 33630 39730
rect 33682 39678 33684 39730
rect 33516 39620 33572 39630
rect 33516 38834 33572 39564
rect 33516 38782 33518 38834
rect 33570 38782 33572 38834
rect 33516 38770 33572 38782
rect 33628 38722 33684 39678
rect 33628 38670 33630 38722
rect 33682 38670 33684 38722
rect 33628 38658 33684 38670
rect 33292 35746 33348 35756
rect 33404 38610 33460 38622
rect 33404 38558 33406 38610
rect 33458 38558 33460 38610
rect 33404 35026 33460 38558
rect 33404 34974 33406 35026
rect 33458 34974 33460 35026
rect 33292 34916 33348 34926
rect 33068 34914 33348 34916
rect 33068 34862 33294 34914
rect 33346 34862 33348 34914
rect 33068 34860 33348 34862
rect 33292 34130 33348 34860
rect 33292 34078 33294 34130
rect 33346 34078 33348 34130
rect 33292 34066 33348 34078
rect 33404 34018 33460 34974
rect 33740 34244 33796 41020
rect 34076 40628 34132 41356
rect 34412 41186 34468 41356
rect 34972 41300 35028 41310
rect 34412 41134 34414 41186
rect 34466 41134 34468 41186
rect 34412 41122 34468 41134
rect 34524 41188 34580 41198
rect 34524 41074 34580 41132
rect 34524 41022 34526 41074
rect 34578 41022 34580 41074
rect 34524 41010 34580 41022
rect 34748 40964 34804 40974
rect 34748 40870 34804 40908
rect 34860 40628 34916 40638
rect 34972 40628 35028 41244
rect 34076 40626 34692 40628
rect 34076 40574 34078 40626
rect 34130 40574 34692 40626
rect 34076 40572 34692 40574
rect 34076 40562 34132 40572
rect 33964 39508 34020 39518
rect 33964 39506 34132 39508
rect 33964 39454 33966 39506
rect 34018 39454 34132 39506
rect 33964 39452 34132 39454
rect 33964 39442 34020 39452
rect 33404 33966 33406 34018
rect 33458 33966 33460 34018
rect 33404 33954 33460 33966
rect 33516 34188 33740 34244
rect 33516 32674 33572 34188
rect 33740 34178 33796 34188
rect 33852 37826 33908 37838
rect 33852 37774 33854 37826
rect 33906 37774 33908 37826
rect 33516 32622 33518 32674
rect 33570 32622 33572 32674
rect 33516 32610 33572 32622
rect 33852 33346 33908 37774
rect 34076 34020 34132 39452
rect 34188 38948 34244 38958
rect 34188 38274 34244 38892
rect 34188 38222 34190 38274
rect 34242 38222 34244 38274
rect 34188 38210 34244 38222
rect 34188 34916 34244 34926
rect 34188 34242 34244 34860
rect 34300 34356 34356 40572
rect 34636 40514 34692 40572
rect 34860 40626 35028 40628
rect 34860 40574 34862 40626
rect 34914 40574 35028 40626
rect 34860 40572 35028 40574
rect 35084 40628 35140 41356
rect 35420 41412 35476 41422
rect 35532 41412 35588 41692
rect 35756 41636 35812 48636
rect 35868 48132 35924 48142
rect 35868 48038 35924 48076
rect 35868 45220 35924 45230
rect 35868 45126 35924 45164
rect 36092 43988 36148 48748
rect 36428 48356 36484 48750
rect 36428 48290 36484 48300
rect 36204 45220 36260 45230
rect 36204 45126 36260 45164
rect 36316 45220 36372 45230
rect 36316 45218 36596 45220
rect 36316 45166 36318 45218
rect 36370 45166 36596 45218
rect 36316 45164 36596 45166
rect 36316 45154 36372 45164
rect 36540 45106 36596 45164
rect 36540 45054 36542 45106
rect 36594 45054 36596 45106
rect 36540 45042 36596 45054
rect 36092 43922 36148 43932
rect 36204 44882 36260 44894
rect 36204 44830 36206 44882
rect 36258 44830 36260 44882
rect 36092 41972 36148 41982
rect 36092 41878 36148 41916
rect 36204 41636 36260 44830
rect 36652 44548 36708 55916
rect 36988 55860 37044 56702
rect 37100 56644 37156 56654
rect 37100 56550 37156 56588
rect 37324 56644 37380 56654
rect 37324 56642 38052 56644
rect 37324 56590 37326 56642
rect 37378 56590 38052 56642
rect 37324 56588 38052 56590
rect 37324 56578 37380 56588
rect 37100 56308 37156 56318
rect 37100 56214 37156 56252
rect 37212 56196 37268 56206
rect 37212 56102 37268 56140
rect 37996 56084 38052 56588
rect 37996 56082 38164 56084
rect 37996 56030 37998 56082
rect 38050 56030 38164 56082
rect 37996 56028 38164 56030
rect 37996 56018 38052 56028
rect 37100 55860 37156 55870
rect 36988 55858 37156 55860
rect 36988 55806 37102 55858
rect 37154 55806 37156 55858
rect 36988 55804 37156 55806
rect 37100 55794 37156 55804
rect 37996 55298 38052 55310
rect 37996 55246 37998 55298
rect 38050 55246 38052 55298
rect 37436 55186 37492 55198
rect 37436 55134 37438 55186
rect 37490 55134 37492 55186
rect 37436 54068 37492 55134
rect 37996 54402 38052 55246
rect 37996 54350 37998 54402
rect 38050 54350 38052 54402
rect 37996 54292 38052 54350
rect 37436 54002 37492 54012
rect 37548 54236 38052 54292
rect 37436 53058 37492 53070
rect 37436 53006 37438 53058
rect 37490 53006 37492 53058
rect 37436 52948 37492 53006
rect 36764 52834 36820 52846
rect 36764 52782 36766 52834
rect 36818 52782 36820 52834
rect 36764 52724 36820 52782
rect 37212 52724 37268 52734
rect 36764 52722 37268 52724
rect 36764 52670 37214 52722
rect 37266 52670 37268 52722
rect 36764 52668 37268 52670
rect 37212 52276 37268 52668
rect 37212 52210 37268 52220
rect 37436 52164 37492 52892
rect 37548 52834 37604 54236
rect 37548 52782 37550 52834
rect 37602 52782 37604 52834
rect 37548 52770 37604 52782
rect 37884 54068 37940 54078
rect 37660 52164 37716 52174
rect 37436 52162 37716 52164
rect 37436 52110 37662 52162
rect 37714 52110 37716 52162
rect 37436 52108 37716 52110
rect 37660 52098 37716 52108
rect 37884 52162 37940 54012
rect 38108 53730 38164 56028
rect 38108 53678 38110 53730
rect 38162 53678 38164 53730
rect 38108 53666 38164 53678
rect 38220 55970 38276 55982
rect 38220 55918 38222 55970
rect 38274 55918 38276 55970
rect 38220 53844 38276 55918
rect 38332 54514 38388 54526
rect 38332 54462 38334 54514
rect 38386 54462 38388 54514
rect 38332 54068 38388 54462
rect 38332 54002 38388 54012
rect 38332 53844 38388 53854
rect 38220 53842 38388 53844
rect 38220 53790 38334 53842
rect 38386 53790 38388 53842
rect 38220 53788 38388 53790
rect 37884 52110 37886 52162
rect 37938 52110 37940 52162
rect 37884 52098 37940 52110
rect 37996 52276 38052 52286
rect 37660 51938 37716 51950
rect 37996 51940 38052 52220
rect 37660 51886 37662 51938
rect 37714 51886 37716 51938
rect 37660 50428 37716 51886
rect 37548 50372 37716 50428
rect 37772 51884 38052 51940
rect 36876 48804 36932 48814
rect 36876 45668 36932 48748
rect 37212 48356 37268 48366
rect 37212 48244 37268 48300
rect 37212 48242 37492 48244
rect 37212 48190 37214 48242
rect 37266 48190 37492 48242
rect 37212 48188 37492 48190
rect 37212 48178 37268 48188
rect 37100 48132 37156 48142
rect 37100 47460 37156 48076
rect 37212 47460 37268 47470
rect 37100 47458 37268 47460
rect 37100 47406 37214 47458
rect 37266 47406 37268 47458
rect 37100 47404 37268 47406
rect 37212 47394 37268 47404
rect 37436 47458 37492 48188
rect 37436 47406 37438 47458
rect 37490 47406 37492 47458
rect 37436 47394 37492 47406
rect 37324 47236 37380 47246
rect 37324 47234 37492 47236
rect 37324 47182 37326 47234
rect 37378 47182 37492 47234
rect 37324 47180 37492 47182
rect 37324 47170 37380 47180
rect 36876 45602 36932 45612
rect 36764 45444 36820 45454
rect 36764 45218 36820 45388
rect 37324 45332 37380 45342
rect 36764 45166 36766 45218
rect 36818 45166 36820 45218
rect 36764 45154 36820 45166
rect 36876 45164 37268 45220
rect 36876 45162 36932 45164
rect 36876 45110 36878 45162
rect 36930 45110 36932 45162
rect 36876 45098 36932 45110
rect 36540 44492 36708 44548
rect 36428 44324 36484 44334
rect 35420 41410 35588 41412
rect 35420 41358 35422 41410
rect 35474 41358 35588 41410
rect 35420 41356 35588 41358
rect 35644 41580 35812 41636
rect 36092 41580 36260 41636
rect 36316 42530 36372 42542
rect 36316 42478 36318 42530
rect 36370 42478 36372 42530
rect 36316 42308 36372 42478
rect 35420 41346 35476 41356
rect 34860 40562 34916 40572
rect 35084 40562 35140 40572
rect 35420 41076 35476 41086
rect 34636 40462 34638 40514
rect 34690 40462 34692 40514
rect 34636 40450 34692 40462
rect 34412 40402 34468 40414
rect 35420 40404 35476 41020
rect 34412 40350 34414 40402
rect 34466 40350 34468 40402
rect 34412 40292 34468 40350
rect 34972 40402 35476 40404
rect 34972 40350 35422 40402
rect 35474 40350 35476 40402
rect 34972 40348 35476 40350
rect 34412 40226 34468 40236
rect 34636 40292 34692 40302
rect 34636 39732 34692 40236
rect 34972 40290 35028 40348
rect 35420 40338 35476 40348
rect 35532 40962 35588 40974
rect 35532 40910 35534 40962
rect 35586 40910 35588 40962
rect 35532 40404 35588 40910
rect 35532 40338 35588 40348
rect 34972 40238 34974 40290
rect 35026 40238 35028 40290
rect 34972 40226 35028 40238
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39732 35140 39742
rect 34636 39676 34916 39732
rect 34412 39284 34468 39294
rect 34412 38162 34468 39228
rect 34636 39058 34692 39676
rect 34636 39006 34638 39058
rect 34690 39006 34692 39058
rect 34636 38994 34692 39006
rect 34748 39506 34804 39518
rect 34748 39454 34750 39506
rect 34802 39454 34804 39506
rect 34748 38836 34804 39454
rect 34860 39506 34916 39676
rect 35084 39618 35140 39676
rect 35084 39566 35086 39618
rect 35138 39566 35140 39618
rect 35084 39554 35140 39566
rect 34860 39454 34862 39506
rect 34914 39454 34916 39506
rect 34860 39442 34916 39454
rect 35084 39284 35140 39294
rect 34748 38770 34804 38780
rect 34972 38948 35028 38958
rect 34412 38110 34414 38162
rect 34466 38110 34468 38162
rect 34412 38098 34468 38110
rect 34972 38162 35028 38892
rect 34972 38110 34974 38162
rect 35026 38110 35028 38162
rect 34972 38098 35028 38110
rect 34972 37380 35028 37390
rect 34748 37268 34804 37278
rect 34748 37174 34804 37212
rect 34412 35812 34468 35822
rect 34412 35698 34468 35756
rect 34412 35646 34414 35698
rect 34466 35646 34468 35698
rect 34412 35634 34468 35646
rect 34860 35700 34916 35710
rect 34860 35586 34916 35644
rect 34860 35534 34862 35586
rect 34914 35534 34916 35586
rect 34860 35522 34916 35534
rect 34972 34914 35028 37324
rect 34972 34862 34974 34914
rect 35026 34862 35028 34914
rect 34972 34850 35028 34862
rect 34748 34692 34804 34702
rect 34748 34598 34804 34636
rect 34300 34300 34580 34356
rect 34188 34190 34190 34242
rect 34242 34190 34244 34242
rect 34188 34178 34244 34190
rect 34412 34020 34468 34030
rect 34076 33964 34356 34020
rect 33852 33294 33854 33346
rect 33906 33294 33908 33346
rect 33852 32562 33908 33294
rect 33852 32510 33854 32562
rect 33906 32510 33908 32562
rect 33852 32498 33908 32510
rect 34188 32788 34244 32798
rect 32956 31826 33012 31836
rect 33292 31666 33348 31678
rect 33292 31614 33294 31666
rect 33346 31614 33348 31666
rect 32956 31554 33012 31566
rect 32956 31502 32958 31554
rect 33010 31502 33012 31554
rect 32956 30212 33012 31502
rect 33292 30772 33348 31614
rect 33292 30706 33348 30716
rect 33068 30212 33124 30222
rect 32956 30210 33124 30212
rect 32956 30158 33070 30210
rect 33122 30158 33124 30210
rect 32956 30156 33124 30158
rect 33068 30146 33124 30156
rect 33852 29988 33908 29998
rect 33740 28868 33796 28878
rect 33180 28866 33796 28868
rect 33180 28814 33742 28866
rect 33794 28814 33796 28866
rect 33180 28812 33796 28814
rect 32956 28420 33012 28430
rect 32956 28418 33124 28420
rect 32956 28366 32958 28418
rect 33010 28366 33124 28418
rect 32956 28364 33124 28366
rect 32956 28354 33012 28364
rect 33068 27970 33124 28364
rect 33180 28082 33236 28812
rect 33740 28802 33796 28812
rect 33180 28030 33182 28082
rect 33234 28030 33236 28082
rect 33180 28018 33236 28030
rect 33628 28530 33684 28542
rect 33628 28478 33630 28530
rect 33682 28478 33684 28530
rect 33068 27918 33070 27970
rect 33122 27918 33124 27970
rect 33068 27906 33124 27918
rect 33180 27636 33236 27646
rect 33180 27542 33236 27580
rect 32844 27356 33572 27412
rect 32732 27234 32788 27244
rect 32620 27074 32676 27086
rect 32620 27022 32622 27074
rect 32674 27022 32676 27074
rect 32396 26852 32564 26908
rect 32172 25788 32452 25844
rect 32172 25506 32228 25788
rect 32172 25454 32174 25506
rect 32226 25454 32228 25506
rect 32172 25442 32228 25454
rect 32284 25618 32340 25630
rect 32284 25566 32286 25618
rect 32338 25566 32340 25618
rect 31836 24948 31892 24958
rect 31836 24722 31892 24892
rect 31948 24836 32004 24846
rect 32284 24836 32340 25566
rect 32396 24946 32452 25788
rect 32396 24894 32398 24946
rect 32450 24894 32452 24946
rect 32396 24882 32452 24894
rect 31948 24834 32340 24836
rect 31948 24782 31950 24834
rect 32002 24782 32286 24834
rect 32338 24782 32340 24834
rect 31948 24780 32340 24782
rect 31948 24770 32004 24780
rect 32284 24770 32340 24780
rect 31836 24670 31838 24722
rect 31890 24670 31892 24722
rect 31836 24050 31892 24670
rect 31836 23998 31838 24050
rect 31890 23998 31892 24050
rect 31836 23986 31892 23998
rect 31948 23940 32004 23950
rect 31948 23846 32004 23884
rect 31724 21868 31892 21924
rect 31724 21698 31780 21710
rect 31724 21646 31726 21698
rect 31778 21646 31780 21698
rect 31612 21364 31668 21374
rect 31276 20974 31278 21026
rect 31330 20974 31332 21026
rect 31276 20962 31332 20974
rect 31388 21362 31668 21364
rect 31388 21310 31614 21362
rect 31666 21310 31668 21362
rect 31388 21308 31668 21310
rect 31276 20244 31332 20254
rect 31388 20244 31444 21308
rect 31612 21298 31668 21308
rect 31724 20916 31780 21646
rect 31724 20850 31780 20860
rect 31276 20242 31444 20244
rect 31276 20190 31278 20242
rect 31330 20190 31444 20242
rect 31276 20188 31444 20190
rect 31612 20802 31668 20814
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 31612 20244 31668 20750
rect 31276 20178 31332 20188
rect 31612 20178 31668 20188
rect 31164 20132 31220 20142
rect 31164 18788 31220 20076
rect 31500 20132 31556 20142
rect 31500 20038 31556 20076
rect 31388 20020 31444 20030
rect 31388 19926 31444 19964
rect 31836 18788 31892 21868
rect 31948 21362 32004 21374
rect 31948 21310 31950 21362
rect 32002 21310 32004 21362
rect 31948 20244 32004 21310
rect 31948 20178 32004 20188
rect 32284 20916 32340 20926
rect 32284 20242 32340 20860
rect 32284 20190 32286 20242
rect 32338 20190 32340 20242
rect 32284 20178 32340 20190
rect 32396 20244 32452 20254
rect 32060 20130 32116 20142
rect 32060 20078 32062 20130
rect 32114 20078 32116 20130
rect 31948 20020 32004 20030
rect 32060 20020 32116 20078
rect 32396 20130 32452 20188
rect 32396 20078 32398 20130
rect 32450 20078 32452 20130
rect 32396 20066 32452 20078
rect 31948 20018 32116 20020
rect 31948 19966 31950 20018
rect 32002 19966 32116 20018
rect 31948 19964 32116 19966
rect 31948 19954 32004 19964
rect 32508 19348 32564 26852
rect 32620 26292 32676 27022
rect 32620 26226 32676 26236
rect 32844 27076 32900 27086
rect 32844 25508 32900 27020
rect 33068 27076 33124 27086
rect 33068 26402 33124 27020
rect 33068 26350 33070 26402
rect 33122 26350 33124 26402
rect 33068 26338 33124 26350
rect 33404 27074 33460 27086
rect 33404 27022 33406 27074
rect 33458 27022 33460 27074
rect 33404 26292 33460 27022
rect 33516 26516 33572 27356
rect 33628 27076 33684 28478
rect 33740 28532 33796 28542
rect 33852 28532 33908 29932
rect 33740 28530 33908 28532
rect 33740 28478 33742 28530
rect 33794 28478 33908 28530
rect 33740 28476 33908 28478
rect 33740 28466 33796 28476
rect 33628 27010 33684 27020
rect 33852 26962 33908 28476
rect 33964 29876 34020 29886
rect 33964 27970 34020 29820
rect 33964 27918 33966 27970
rect 34018 27918 34020 27970
rect 33964 27906 34020 27918
rect 33852 26910 33854 26962
rect 33906 26910 33908 26962
rect 33852 26898 33908 26910
rect 34188 26908 34244 32732
rect 33516 26450 33572 26460
rect 34076 26852 34244 26908
rect 33516 26292 33572 26302
rect 33404 26290 33572 26292
rect 33404 26238 33518 26290
rect 33570 26238 33572 26290
rect 33404 26236 33572 26238
rect 32844 25452 33236 25508
rect 32620 25396 32676 25406
rect 32620 25394 33124 25396
rect 32620 25342 32622 25394
rect 32674 25342 33124 25394
rect 32620 25340 33124 25342
rect 32620 25330 32676 25340
rect 32620 24724 32676 24734
rect 32956 24724 33012 24734
rect 32620 24722 33012 24724
rect 32620 24670 32622 24722
rect 32674 24670 32958 24722
rect 33010 24670 33012 24722
rect 32620 24668 33012 24670
rect 32620 24658 32676 24668
rect 32956 24658 33012 24668
rect 32956 23940 33012 23950
rect 33068 23940 33124 25340
rect 32956 23938 33124 23940
rect 32956 23886 32958 23938
rect 33010 23886 33124 23938
rect 32956 23884 33124 23886
rect 32956 23874 33012 23884
rect 32620 23828 32676 23838
rect 32620 23826 32788 23828
rect 32620 23774 32622 23826
rect 32674 23774 32788 23826
rect 32620 23772 32788 23774
rect 32620 23762 32676 23772
rect 32620 20916 32676 20926
rect 32620 20822 32676 20860
rect 32620 19348 32676 19358
rect 32284 19346 32676 19348
rect 32284 19294 32622 19346
rect 32674 19294 32676 19346
rect 32284 19292 32676 19294
rect 31164 18722 31220 18732
rect 31612 18732 31892 18788
rect 31948 18788 32004 18798
rect 31164 18338 31220 18350
rect 31164 18286 31166 18338
rect 31218 18286 31220 18338
rect 31164 17780 31220 18286
rect 31164 17714 31220 17724
rect 31276 17780 31332 17790
rect 31612 17780 31668 18732
rect 31948 18676 32004 18732
rect 31948 18674 32228 18676
rect 31948 18622 31950 18674
rect 32002 18622 32228 18674
rect 31948 18620 32228 18622
rect 31948 18610 32004 18620
rect 31724 18564 31780 18574
rect 31724 18470 31780 18508
rect 31836 18338 31892 18350
rect 31836 18286 31838 18338
rect 31890 18286 31892 18338
rect 31724 17780 31780 17790
rect 31276 17778 31724 17780
rect 31276 17726 31278 17778
rect 31330 17726 31724 17778
rect 31276 17724 31724 17726
rect 31276 17714 31332 17724
rect 31724 17686 31780 17724
rect 31164 17444 31220 17454
rect 31164 17350 31220 17388
rect 31164 16884 31220 16894
rect 31164 16098 31220 16828
rect 31836 16882 31892 18286
rect 32172 18004 32228 18620
rect 32284 18450 32340 19292
rect 32620 19282 32676 19292
rect 32284 18398 32286 18450
rect 32338 18398 32340 18450
rect 32284 18386 32340 18398
rect 32172 17948 32452 18004
rect 31836 16830 31838 16882
rect 31890 16830 31892 16882
rect 31276 16770 31332 16782
rect 31276 16718 31278 16770
rect 31330 16718 31332 16770
rect 31276 16212 31332 16718
rect 31276 16118 31332 16156
rect 31164 16046 31166 16098
rect 31218 16046 31220 16098
rect 31164 15314 31220 16046
rect 31164 15262 31166 15314
rect 31218 15262 31220 15314
rect 31164 15250 31220 15262
rect 31836 15314 31892 16830
rect 32060 16884 32116 16894
rect 32060 16790 32116 16828
rect 32060 16100 32116 16110
rect 32172 16100 32228 17948
rect 32284 17780 32340 17790
rect 32284 17108 32340 17724
rect 32396 17778 32452 17948
rect 32396 17726 32398 17778
rect 32450 17726 32452 17778
rect 32396 17714 32452 17726
rect 32284 17106 32564 17108
rect 32284 17054 32286 17106
rect 32338 17054 32564 17106
rect 32284 17052 32564 17054
rect 32284 17042 32340 17052
rect 32116 16044 32228 16100
rect 32396 16882 32452 16894
rect 32396 16830 32398 16882
rect 32450 16830 32452 16882
rect 32396 16322 32452 16830
rect 32396 16270 32398 16322
rect 32450 16270 32452 16322
rect 32060 16006 32116 16044
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31836 15250 31892 15262
rect 31948 15090 32004 15102
rect 31948 15038 31950 15090
rect 32002 15038 32004 15090
rect 31164 14644 31220 14654
rect 31612 14644 31668 14654
rect 31108 14642 31668 14644
rect 31108 14590 31166 14642
rect 31218 14590 31614 14642
rect 31666 14590 31668 14642
rect 31108 14588 31668 14590
rect 31052 13860 31108 14588
rect 31164 14578 31220 14588
rect 31612 14578 31668 14588
rect 31052 13794 31108 13804
rect 31836 13972 31892 13982
rect 31836 13746 31892 13916
rect 31836 13694 31838 13746
rect 31890 13694 31892 13746
rect 31836 13682 31892 13694
rect 31276 13524 31332 13534
rect 31612 13524 31668 13534
rect 31164 13522 31332 13524
rect 31164 13470 31278 13522
rect 31330 13470 31332 13522
rect 31164 13468 31332 13470
rect 31164 10276 31220 13468
rect 31276 13458 31332 13468
rect 31388 13522 31668 13524
rect 31388 13470 31614 13522
rect 31666 13470 31668 13522
rect 31388 13468 31668 13470
rect 31276 12404 31332 12414
rect 31388 12404 31444 13468
rect 31612 13458 31668 13468
rect 31948 13188 32004 15038
rect 32060 14756 32116 14766
rect 32060 14642 32116 14700
rect 32060 14590 32062 14642
rect 32114 14590 32116 14642
rect 32060 14578 32116 14590
rect 32396 14308 32452 16270
rect 32508 16210 32564 17052
rect 32508 16158 32510 16210
rect 32562 16158 32564 16210
rect 32508 16146 32564 16158
rect 32732 15148 32788 23772
rect 33068 23716 33124 23726
rect 33068 23622 33124 23660
rect 32956 20804 33012 20814
rect 33180 20804 33236 25452
rect 33516 24724 33572 26236
rect 33852 26292 33908 26302
rect 33852 26178 33908 26236
rect 33852 26126 33854 26178
rect 33906 26126 33908 26178
rect 33852 24836 33908 26126
rect 34076 25618 34132 26852
rect 34076 25566 34078 25618
rect 34130 25566 34132 25618
rect 34076 25554 34132 25566
rect 33964 25282 34020 25294
rect 33964 25230 33966 25282
rect 34018 25230 34020 25282
rect 33964 24948 34020 25230
rect 33964 24882 34020 24892
rect 33516 24658 33572 24668
rect 33628 24780 33908 24836
rect 33628 24610 33684 24780
rect 33628 24558 33630 24610
rect 33682 24558 33684 24610
rect 33292 20804 33348 20814
rect 32956 20802 33124 20804
rect 32956 20750 32958 20802
rect 33010 20750 33124 20802
rect 32956 20748 33124 20750
rect 33180 20748 33292 20804
rect 32956 20738 33012 20748
rect 33068 20132 33124 20748
rect 33292 20738 33348 20748
rect 33068 19348 33124 20076
rect 33068 19282 33124 19292
rect 33292 20244 33348 20254
rect 33292 18452 33348 20188
rect 33404 20244 33460 20254
rect 33628 20244 33684 24558
rect 33964 24724 34020 24734
rect 33740 24498 33796 24510
rect 33740 24446 33742 24498
rect 33794 24446 33796 24498
rect 33740 20916 33796 24446
rect 33852 23826 33908 23838
rect 33852 23774 33854 23826
rect 33906 23774 33908 23826
rect 33852 23268 33908 23774
rect 33964 23716 34020 24668
rect 34188 23938 34244 23950
rect 34188 23886 34190 23938
rect 34242 23886 34244 23938
rect 33964 23650 34020 23660
rect 34076 23828 34132 23838
rect 34188 23828 34244 23886
rect 34132 23772 34244 23828
rect 33852 23044 33908 23212
rect 33964 23154 34020 23166
rect 33964 23102 33966 23154
rect 34018 23102 34020 23154
rect 33964 23044 34020 23102
rect 33908 22988 34020 23044
rect 34076 23044 34132 23772
rect 33852 22978 33908 22988
rect 34076 22950 34132 22988
rect 33740 20850 33796 20860
rect 33852 21028 33908 21038
rect 33404 20242 33684 20244
rect 33404 20190 33406 20242
rect 33458 20190 33684 20242
rect 33404 20188 33684 20190
rect 33404 20178 33460 20188
rect 33740 19348 33796 19358
rect 33740 19254 33796 19292
rect 33404 19234 33460 19246
rect 33404 19182 33406 19234
rect 33458 19182 33460 19234
rect 33404 18674 33460 19182
rect 33628 19236 33684 19246
rect 33628 19142 33684 19180
rect 33852 19012 33908 20972
rect 34300 20356 34356 33964
rect 34412 33346 34468 33964
rect 34412 33294 34414 33346
rect 34466 33294 34468 33346
rect 34412 33282 34468 33294
rect 34524 32340 34580 34300
rect 34636 34244 34692 34254
rect 34636 34150 34692 34188
rect 34748 34018 34804 34030
rect 34748 33966 34750 34018
rect 34802 33966 34804 34018
rect 34748 33346 34804 33966
rect 34748 33294 34750 33346
rect 34802 33294 34804 33346
rect 34748 33282 34804 33294
rect 34860 33908 34916 33918
rect 34748 33122 34804 33134
rect 34748 33070 34750 33122
rect 34802 33070 34804 33122
rect 34748 32564 34804 33070
rect 34748 32498 34804 32508
rect 34860 32562 34916 33852
rect 34972 32788 35028 32798
rect 34972 32694 35028 32732
rect 34860 32510 34862 32562
rect 34914 32510 34916 32562
rect 34860 32498 34916 32510
rect 34524 32284 34916 32340
rect 34412 31892 34468 31902
rect 34412 31778 34468 31836
rect 34412 31726 34414 31778
rect 34466 31726 34468 31778
rect 34412 31714 34468 31726
rect 34524 31780 34580 31790
rect 34524 31666 34580 31724
rect 34524 31614 34526 31666
rect 34578 31614 34580 31666
rect 34524 31602 34580 31614
rect 34636 31668 34692 31678
rect 34412 31108 34468 31118
rect 34636 31108 34692 31612
rect 34412 31106 34692 31108
rect 34412 31054 34414 31106
rect 34466 31054 34692 31106
rect 34412 31052 34692 31054
rect 34748 31554 34804 31566
rect 34748 31502 34750 31554
rect 34802 31502 34804 31554
rect 34412 31042 34468 31052
rect 34524 30770 34580 30782
rect 34524 30718 34526 30770
rect 34578 30718 34580 30770
rect 34524 30100 34580 30718
rect 34748 30212 34804 31502
rect 34748 30146 34804 30156
rect 34524 30034 34580 30044
rect 34860 29988 34916 32284
rect 34748 29932 34916 29988
rect 34748 26908 34804 29932
rect 35084 29652 35140 39228
rect 35644 39172 35700 41580
rect 35756 41188 35812 41198
rect 35756 41094 35812 41132
rect 35980 40962 36036 40974
rect 35980 40910 35982 40962
rect 36034 40910 36036 40962
rect 35980 40516 36036 40910
rect 35868 40460 36036 40516
rect 35868 40402 35924 40460
rect 35868 40350 35870 40402
rect 35922 40350 35924 40402
rect 35868 39618 35924 40350
rect 35980 40290 36036 40302
rect 35980 40238 35982 40290
rect 36034 40238 36036 40290
rect 35980 39732 36036 40238
rect 35980 39638 36036 39676
rect 35868 39566 35870 39618
rect 35922 39566 35924 39618
rect 35868 39554 35924 39566
rect 35868 39172 35924 39182
rect 35644 39116 35868 39172
rect 35868 39106 35924 39116
rect 35196 38836 35252 38846
rect 35196 38742 35252 38780
rect 35868 38724 35924 38734
rect 35756 38668 35868 38724
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35532 35812 35588 35822
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 34916 35252 34926
rect 35532 34916 35588 35756
rect 35756 35308 35812 38668
rect 35868 38658 35924 38668
rect 36092 38724 36148 41580
rect 36204 41412 36260 41422
rect 36316 41412 36372 42252
rect 36260 41356 36372 41412
rect 36204 41346 36260 41356
rect 36316 41076 36372 41086
rect 36316 40982 36372 41020
rect 36204 40964 36260 40974
rect 36204 40870 36260 40908
rect 36092 38658 36148 38668
rect 36204 40178 36260 40190
rect 36204 40126 36206 40178
rect 36258 40126 36260 40178
rect 36204 38668 36260 40126
rect 36316 39732 36372 39742
rect 36428 39732 36484 44268
rect 36316 39730 36484 39732
rect 36316 39678 36318 39730
rect 36370 39678 36484 39730
rect 36316 39676 36484 39678
rect 36316 39666 36372 39676
rect 36428 39172 36484 39182
rect 36204 38612 36372 38668
rect 36092 38500 36148 38510
rect 35756 35252 35924 35308
rect 35196 34242 35252 34860
rect 35420 34860 35588 34916
rect 35868 34916 35924 35252
rect 35868 34860 36036 34916
rect 35308 34690 35364 34702
rect 35308 34638 35310 34690
rect 35362 34638 35364 34690
rect 35308 34356 35364 34638
rect 35308 34290 35364 34300
rect 35196 34190 35198 34242
rect 35250 34190 35252 34242
rect 35196 34178 35252 34190
rect 35420 34244 35476 34860
rect 35644 34804 35700 34814
rect 35644 34802 35812 34804
rect 35644 34750 35646 34802
rect 35698 34750 35812 34802
rect 35644 34748 35812 34750
rect 35644 34738 35700 34748
rect 35532 34690 35588 34702
rect 35532 34638 35534 34690
rect 35586 34638 35588 34690
rect 35532 34468 35588 34638
rect 35532 34402 35588 34412
rect 35756 34692 35812 34748
rect 35868 34692 35924 34702
rect 35756 34690 35924 34692
rect 35756 34638 35870 34690
rect 35922 34638 35924 34690
rect 35756 34636 35924 34638
rect 35532 34244 35588 34254
rect 35420 34188 35532 34244
rect 35532 34178 35588 34188
rect 35308 33908 35364 33918
rect 35756 33908 35812 34636
rect 35868 34626 35924 34636
rect 35868 34244 35924 34254
rect 35868 34150 35924 34188
rect 35308 33906 35700 33908
rect 35308 33854 35310 33906
rect 35362 33854 35700 33906
rect 35308 33852 35700 33854
rect 35308 33842 35364 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35644 31892 35700 33852
rect 35756 33842 35812 33852
rect 35980 31892 36036 34860
rect 36092 34802 36148 38444
rect 36092 34750 36094 34802
rect 36146 34750 36148 34802
rect 36092 34738 36148 34750
rect 36204 34802 36260 34814
rect 36204 34750 36206 34802
rect 36258 34750 36260 34802
rect 36204 34692 36260 34750
rect 36204 34626 36260 34636
rect 35644 31798 35700 31836
rect 35756 31836 36036 31892
rect 35532 31780 35588 31790
rect 35532 31668 35588 31724
rect 35756 31668 35812 31836
rect 35532 31612 35812 31668
rect 35980 31668 36036 31678
rect 35980 31574 36036 31612
rect 36204 30994 36260 31006
rect 36204 30942 36206 30994
rect 36258 30942 36260 30994
rect 35308 30772 35364 30810
rect 35308 30706 35364 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35420 30212 35476 30222
rect 35420 30118 35476 30156
rect 36204 30212 36260 30942
rect 36204 30146 36260 30156
rect 35084 28868 35140 29596
rect 35868 30100 35924 30110
rect 35868 29314 35924 30044
rect 36092 30098 36148 30110
rect 36092 30046 36094 30098
rect 36146 30046 36148 30098
rect 35980 29988 36036 29998
rect 36092 29988 36148 30046
rect 36204 29988 36260 29998
rect 36092 29932 36204 29988
rect 35980 29894 36036 29932
rect 36204 29922 36260 29932
rect 36316 29764 36372 38612
rect 36428 36932 36484 39116
rect 36540 38668 36596 44492
rect 37100 44324 37156 44334
rect 37212 44324 37268 45164
rect 37156 44268 37268 44324
rect 37324 44322 37380 45276
rect 37436 44996 37492 47180
rect 37548 46228 37604 50372
rect 37660 48802 37716 48814
rect 37660 48750 37662 48802
rect 37714 48750 37716 48802
rect 37660 47346 37716 48750
rect 37660 47294 37662 47346
rect 37714 47294 37716 47346
rect 37660 47282 37716 47294
rect 37548 46162 37604 46172
rect 37772 45892 37828 51884
rect 37884 50594 37940 50606
rect 37884 50542 37886 50594
rect 37938 50542 37940 50594
rect 37884 50428 37940 50542
rect 38108 50484 38164 50494
rect 37884 50372 38164 50428
rect 37996 48914 38052 48926
rect 37996 48862 37998 48914
rect 38050 48862 38052 48914
rect 37884 48802 37940 48814
rect 37884 48750 37886 48802
rect 37938 48750 37940 48802
rect 37884 48356 37940 48750
rect 37884 48262 37940 48300
rect 37996 48132 38052 48862
rect 37996 48066 38052 48076
rect 38108 48020 38164 50372
rect 38220 48354 38276 53788
rect 38332 53778 38388 53788
rect 38332 50596 38388 50606
rect 38556 50596 38612 59052
rect 38668 58996 38724 60060
rect 38892 60002 38948 60014
rect 38892 59950 38894 60002
rect 38946 59950 38948 60002
rect 38892 59108 38948 59950
rect 39004 59108 39060 59118
rect 38892 59052 39004 59108
rect 39004 59014 39060 59052
rect 38724 58940 38948 58996
rect 38668 58930 38724 58940
rect 38892 58322 38948 58940
rect 39116 58884 39172 60060
rect 38892 58270 38894 58322
rect 38946 58270 38948 58322
rect 38892 58258 38948 58270
rect 39004 58828 39172 58884
rect 38892 57876 38948 57886
rect 39004 57876 39060 58828
rect 39228 58212 39284 58222
rect 39228 58118 39284 58156
rect 38892 57874 39060 57876
rect 38892 57822 38894 57874
rect 38946 57822 39060 57874
rect 38892 57820 39060 57822
rect 38892 57810 38948 57820
rect 39116 57762 39172 57774
rect 39116 57710 39118 57762
rect 39170 57710 39172 57762
rect 38668 57652 38724 57662
rect 39116 57652 39172 57710
rect 38668 57650 39172 57652
rect 38668 57598 38670 57650
rect 38722 57598 39172 57650
rect 38668 57596 39172 57598
rect 38668 57586 38724 57596
rect 38892 56644 38948 56654
rect 39116 56644 39172 57596
rect 39228 57652 39284 57662
rect 39228 57558 39284 57596
rect 38892 56642 39172 56644
rect 38892 56590 38894 56642
rect 38946 56590 39172 56642
rect 38892 56588 39172 56590
rect 38892 56196 38948 56588
rect 38892 56130 38948 56140
rect 38668 55970 38724 55982
rect 38668 55918 38670 55970
rect 38722 55918 38724 55970
rect 38668 55300 38724 55918
rect 39340 55410 39396 62132
rect 40348 61794 40404 64092
rect 40684 64082 40740 64092
rect 41020 64596 41076 64606
rect 41020 63700 41076 64540
rect 41244 64596 41300 64606
rect 41356 64596 41412 65324
rect 41244 64594 41412 64596
rect 41244 64542 41246 64594
rect 41298 64542 41412 64594
rect 41244 64540 41412 64542
rect 41244 64530 41300 64540
rect 41020 63634 41076 63644
rect 42252 63252 42308 65436
rect 42364 65426 42420 65436
rect 42812 65380 42868 65390
rect 42812 65378 43092 65380
rect 42812 65326 42814 65378
rect 42866 65326 43092 65378
rect 42812 65324 43092 65326
rect 42812 65314 42868 65324
rect 43036 64148 43092 65324
rect 42924 64146 43092 64148
rect 42924 64094 43038 64146
rect 43090 64094 43092 64146
rect 42924 64092 43092 64094
rect 42924 63362 42980 64092
rect 43036 64082 43092 64092
rect 43148 63812 43204 63822
rect 42924 63310 42926 63362
rect 42978 63310 42980 63362
rect 42924 63298 42980 63310
rect 43036 63810 43204 63812
rect 43036 63758 43150 63810
rect 43202 63758 43204 63810
rect 43036 63756 43204 63758
rect 42252 63250 42420 63252
rect 42252 63198 42254 63250
rect 42306 63198 42420 63250
rect 42252 63196 42420 63198
rect 42252 63186 42308 63196
rect 42364 63028 42420 63196
rect 42364 62972 42756 63028
rect 42700 62914 42756 62972
rect 42700 62862 42702 62914
rect 42754 62862 42756 62914
rect 42700 62850 42756 62862
rect 42812 62916 42868 62926
rect 42812 62822 42868 62860
rect 43036 62692 43092 63756
rect 43148 63746 43204 63756
rect 43260 63250 43316 66780
rect 43484 63812 43540 67566
rect 43820 67228 43876 67678
rect 44380 67228 44436 74956
rect 45500 74004 45556 76302
rect 45500 73938 45556 73948
rect 43820 67172 44324 67228
rect 44380 67172 44548 67228
rect 44268 67060 44324 67172
rect 44380 67060 44436 67070
rect 44268 67058 44436 67060
rect 44268 67006 44382 67058
rect 44434 67006 44436 67058
rect 44268 67004 44436 67006
rect 44380 66994 44436 67004
rect 44268 66836 44324 66846
rect 44268 66742 44324 66780
rect 43484 63746 43540 63756
rect 44268 63700 44324 63710
rect 44268 63606 44324 63644
rect 43260 63198 43262 63250
rect 43314 63198 43316 63250
rect 43260 63186 43316 63198
rect 44044 63250 44100 63262
rect 44044 63198 44046 63250
rect 44098 63198 44100 63250
rect 42476 62636 43092 62692
rect 43932 63138 43988 63150
rect 43932 63086 43934 63138
rect 43986 63086 43988 63138
rect 42476 62466 42532 62636
rect 42476 62414 42478 62466
rect 42530 62414 42532 62466
rect 42476 62402 42532 62414
rect 43260 62468 43316 62478
rect 40348 61742 40350 61794
rect 40402 61742 40404 61794
rect 40348 61730 40404 61742
rect 41580 62354 41636 62366
rect 41580 62302 41582 62354
rect 41634 62302 41636 62354
rect 41020 61572 41076 61582
rect 41020 61478 41076 61516
rect 39452 61460 39508 61470
rect 39452 60788 39508 61404
rect 41020 61012 41076 61022
rect 41020 60918 41076 60956
rect 40012 60898 40068 60910
rect 41356 60900 41412 60910
rect 40012 60846 40014 60898
rect 40066 60846 40068 60898
rect 40012 60788 40068 60846
rect 41244 60898 41412 60900
rect 41244 60846 41358 60898
rect 41410 60846 41412 60898
rect 41244 60844 41412 60846
rect 40908 60788 40964 60798
rect 39452 60786 39620 60788
rect 39452 60734 39454 60786
rect 39506 60734 39620 60786
rect 39452 60732 39620 60734
rect 39452 60722 39508 60732
rect 39564 60116 39620 60732
rect 40012 60722 40068 60732
rect 40236 60786 40964 60788
rect 40236 60734 40910 60786
rect 40962 60734 40964 60786
rect 40236 60732 40964 60734
rect 39564 60022 39620 60060
rect 39788 60340 39844 60350
rect 39788 60226 39844 60284
rect 39788 60174 39790 60226
rect 39842 60174 39844 60226
rect 39564 59106 39620 59118
rect 39564 59054 39566 59106
rect 39618 59054 39620 59106
rect 39564 58212 39620 59054
rect 39788 58434 39844 60174
rect 40124 60228 40180 60238
rect 40236 60228 40292 60732
rect 40908 60722 40964 60732
rect 41132 60788 41188 60798
rect 41132 60694 41188 60732
rect 40124 60226 40292 60228
rect 40124 60174 40126 60226
rect 40178 60174 40292 60226
rect 40124 60172 40292 60174
rect 40348 60564 40404 60574
rect 40124 60162 40180 60172
rect 39900 59108 39956 59118
rect 39900 59014 39956 59052
rect 39788 58382 39790 58434
rect 39842 58382 39844 58434
rect 39788 58370 39844 58382
rect 40124 58324 40180 58334
rect 40124 58230 40180 58268
rect 40012 58212 40068 58222
rect 39564 58146 39620 58156
rect 39900 58156 40012 58212
rect 39676 57652 39732 57662
rect 39676 57558 39732 57596
rect 39340 55358 39342 55410
rect 39394 55358 39396 55410
rect 39340 55346 39396 55358
rect 39788 56196 39844 56206
rect 38668 55244 39172 55300
rect 39116 55188 39172 55244
rect 39116 55186 39396 55188
rect 39116 55134 39118 55186
rect 39170 55134 39396 55186
rect 39116 55132 39396 55134
rect 39116 55122 39172 55132
rect 38780 54684 39284 54740
rect 38780 54626 38836 54684
rect 38780 54574 38782 54626
rect 38834 54574 38836 54626
rect 38780 54562 38836 54574
rect 39228 54626 39284 54684
rect 39228 54574 39230 54626
rect 39282 54574 39284 54626
rect 39228 54562 39284 54574
rect 39340 54516 39396 55132
rect 39452 54516 39508 54526
rect 39340 54514 39508 54516
rect 39340 54462 39454 54514
rect 39506 54462 39508 54514
rect 39340 54460 39508 54462
rect 39452 54450 39508 54460
rect 39228 54402 39284 54414
rect 39228 54350 39230 54402
rect 39282 54350 39284 54402
rect 39228 54292 39284 54350
rect 39228 54226 39284 54236
rect 38780 54180 38836 54190
rect 38668 54124 38780 54180
rect 38668 53954 38724 54124
rect 38780 54114 38836 54124
rect 38668 53902 38670 53954
rect 38722 53902 38724 53954
rect 38668 53890 38724 53902
rect 39116 52836 39172 52846
rect 39116 52162 39172 52780
rect 39564 52724 39620 52734
rect 39564 52274 39620 52668
rect 39564 52222 39566 52274
rect 39618 52222 39620 52274
rect 39564 52210 39620 52222
rect 39116 52110 39118 52162
rect 39170 52110 39172 52162
rect 38892 51604 38948 51614
rect 38668 51156 38724 51166
rect 38724 51100 38836 51156
rect 38668 51090 38724 51100
rect 38388 50540 38612 50596
rect 38332 50502 38388 50540
rect 38780 49140 38836 51100
rect 38892 50484 38948 51548
rect 39116 51378 39172 52110
rect 39116 51326 39118 51378
rect 39170 51326 39172 51378
rect 39116 51314 39172 51326
rect 38892 50418 38948 50428
rect 39452 50708 39508 50718
rect 38892 49140 38948 49150
rect 38780 49138 39172 49140
rect 38780 49086 38894 49138
rect 38946 49086 39172 49138
rect 38780 49084 39172 49086
rect 38892 49074 38948 49084
rect 38668 49028 38724 49038
rect 39116 49028 39172 49084
rect 39228 49028 39284 49038
rect 38724 48972 38836 49028
rect 39116 49026 39284 49028
rect 39116 48974 39230 49026
rect 39282 48974 39284 49026
rect 39116 48972 39284 48974
rect 38668 48962 38724 48972
rect 38220 48302 38222 48354
rect 38274 48302 38276 48354
rect 38220 48290 38276 48302
rect 38668 48356 38724 48366
rect 38668 48242 38724 48300
rect 38668 48190 38670 48242
rect 38722 48190 38724 48242
rect 38668 48178 38724 48190
rect 38556 48132 38612 48142
rect 38108 47964 38276 48020
rect 37436 44930 37492 44940
rect 37548 45836 37828 45892
rect 38108 47236 38164 47246
rect 38108 46562 38164 47180
rect 38108 46510 38110 46562
rect 38162 46510 38164 46562
rect 37324 44270 37326 44322
rect 37378 44270 37380 44322
rect 37100 44230 37156 44268
rect 37324 44258 37380 44270
rect 37548 42866 37604 45836
rect 37772 45556 37828 45566
rect 37772 44884 37828 45500
rect 37772 44818 37828 44828
rect 37884 44996 37940 45006
rect 37772 44660 37828 44670
rect 37772 43764 37828 44604
rect 37772 43698 37828 43708
rect 37884 44324 37940 44940
rect 37996 44994 38052 45006
rect 37996 44942 37998 44994
rect 38050 44942 38052 44994
rect 37996 44884 38052 44942
rect 37996 44548 38052 44828
rect 38108 44660 38164 46510
rect 38220 44660 38276 47964
rect 38444 47236 38500 47246
rect 38444 47142 38500 47180
rect 38332 45218 38388 45230
rect 38332 45166 38334 45218
rect 38386 45166 38388 45218
rect 38332 45108 38388 45166
rect 38332 45042 38388 45052
rect 38444 44660 38500 44670
rect 38220 44604 38444 44660
rect 38108 44594 38164 44604
rect 38444 44594 38500 44604
rect 37996 44482 38052 44492
rect 37884 43538 37940 44268
rect 37996 44324 38052 44334
rect 38444 44324 38500 44334
rect 37996 44322 38500 44324
rect 37996 44270 37998 44322
rect 38050 44270 38446 44322
rect 38498 44270 38500 44322
rect 37996 44268 38500 44270
rect 37996 44258 38052 44268
rect 37884 43486 37886 43538
rect 37938 43486 37940 43538
rect 37884 43474 37940 43486
rect 37996 43764 38052 43774
rect 37548 42814 37550 42866
rect 37602 42814 37604 42866
rect 37548 42802 37604 42814
rect 37436 42754 37492 42766
rect 37436 42702 37438 42754
rect 37490 42702 37492 42754
rect 37212 42644 37268 42654
rect 37212 42642 37380 42644
rect 37212 42590 37214 42642
rect 37266 42590 37380 42642
rect 37212 42588 37380 42590
rect 37212 42578 37268 42588
rect 36652 42308 36708 42318
rect 36652 42194 36708 42252
rect 36652 42142 36654 42194
rect 36706 42142 36708 42194
rect 36652 42130 36708 42142
rect 36764 42084 36820 42094
rect 36764 41990 36820 42028
rect 37212 41858 37268 41870
rect 37212 41806 37214 41858
rect 37266 41806 37268 41858
rect 36652 41748 36708 41758
rect 37212 41748 37268 41806
rect 36652 41746 37268 41748
rect 36652 41694 36654 41746
rect 36706 41694 37268 41746
rect 36652 41692 37268 41694
rect 36652 41682 36708 41692
rect 37212 41410 37268 41692
rect 37212 41358 37214 41410
rect 37266 41358 37268 41410
rect 37212 41346 37268 41358
rect 37324 41300 37380 42588
rect 37436 42532 37492 42702
rect 37436 42466 37492 42476
rect 37324 41234 37380 41244
rect 37436 41972 37492 41982
rect 37436 41074 37492 41916
rect 37436 41022 37438 41074
rect 37490 41022 37492 41074
rect 37436 41010 37492 41022
rect 37324 40962 37380 40974
rect 37324 40910 37326 40962
rect 37378 40910 37380 40962
rect 37324 40290 37380 40910
rect 37436 40404 37492 40414
rect 37436 40310 37492 40348
rect 37324 40238 37326 40290
rect 37378 40238 37380 40290
rect 37324 40226 37380 40238
rect 37548 40292 37604 40302
rect 37324 38836 37380 38846
rect 37324 38668 37380 38780
rect 37548 38668 37604 40236
rect 37884 40180 37940 40190
rect 36540 38612 36820 38668
rect 37324 38612 37604 38668
rect 36428 35698 36484 36876
rect 36428 35646 36430 35698
rect 36482 35646 36484 35698
rect 36428 35634 36484 35646
rect 36540 32676 36596 32686
rect 35868 29262 35870 29314
rect 35922 29262 35924 29314
rect 35868 29250 35924 29262
rect 35980 29708 36372 29764
rect 36428 32564 36484 32574
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28802 35140 28812
rect 35308 28868 35364 28878
rect 34972 28532 35028 28542
rect 34972 27858 35028 28476
rect 35196 28532 35252 28542
rect 35196 28438 35252 28476
rect 35308 27972 35364 28812
rect 35532 28866 35588 28878
rect 35532 28814 35534 28866
rect 35586 28814 35588 28866
rect 35420 28644 35476 28654
rect 35420 28530 35476 28588
rect 35420 28478 35422 28530
rect 35474 28478 35476 28530
rect 35420 28466 35476 28478
rect 35308 27906 35364 27916
rect 34972 27806 34974 27858
rect 35026 27806 35028 27858
rect 34972 27794 35028 27806
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35308 27300 35364 27310
rect 35308 27206 35364 27244
rect 35532 27186 35588 28814
rect 35980 28756 36036 29708
rect 36428 29538 36484 32508
rect 36540 30994 36596 32620
rect 36540 30942 36542 30994
rect 36594 30942 36596 30994
rect 36540 30930 36596 30942
rect 36428 29486 36430 29538
rect 36482 29486 36484 29538
rect 36428 29474 36484 29486
rect 35756 28700 36036 28756
rect 35756 27858 35812 28700
rect 35980 28644 36036 28700
rect 35868 28532 35924 28542
rect 35868 28196 35924 28476
rect 35980 28530 36036 28588
rect 35980 28478 35982 28530
rect 36034 28478 36036 28530
rect 35980 28466 36036 28478
rect 36204 28418 36260 28430
rect 36204 28366 36206 28418
rect 36258 28366 36260 28418
rect 35868 28140 36036 28196
rect 35756 27806 35758 27858
rect 35810 27806 35812 27858
rect 35756 27794 35812 27806
rect 35868 27972 35924 27982
rect 35532 27134 35534 27186
rect 35586 27134 35588 27186
rect 35532 27122 35588 27134
rect 35644 27636 35700 27646
rect 35420 27074 35476 27086
rect 35420 27022 35422 27074
rect 35474 27022 35476 27074
rect 35420 26964 35476 27022
rect 35644 26964 35700 27580
rect 35420 26908 35700 26964
rect 35868 26908 35924 27916
rect 34300 20290 34356 20300
rect 34636 26852 34804 26908
rect 35756 26852 35924 26908
rect 35980 26908 36036 28140
rect 36092 27970 36148 27982
rect 36092 27918 36094 27970
rect 36146 27918 36148 27970
rect 36092 27636 36148 27918
rect 36092 27570 36148 27580
rect 36204 27074 36260 28366
rect 36204 27022 36206 27074
rect 36258 27022 36260 27074
rect 36204 27010 36260 27022
rect 35980 26852 36148 26908
rect 34300 20018 34356 20030
rect 34300 19966 34302 20018
rect 34354 19966 34356 20018
rect 34188 19348 34244 19358
rect 33964 19346 34244 19348
rect 33964 19294 34190 19346
rect 34242 19294 34244 19346
rect 33964 19292 34244 19294
rect 33964 19234 34020 19292
rect 34188 19282 34244 19292
rect 33964 19182 33966 19234
rect 34018 19182 34020 19234
rect 33964 19170 34020 19182
rect 33404 18622 33406 18674
rect 33458 18622 33460 18674
rect 33404 18610 33460 18622
rect 33628 18956 33908 19012
rect 33292 18396 33460 18452
rect 33292 16994 33348 17006
rect 33292 16942 33294 16994
rect 33346 16942 33348 16994
rect 32956 16324 33012 16334
rect 33292 16324 33348 16942
rect 32956 16322 33348 16324
rect 32956 16270 32958 16322
rect 33010 16270 33348 16322
rect 32956 16268 33348 16270
rect 32956 16258 33012 16268
rect 32844 16100 32900 16110
rect 32844 16006 32900 16044
rect 32396 14242 32452 14252
rect 32620 15092 32788 15148
rect 32284 13972 32340 13982
rect 32284 13878 32340 13916
rect 31948 13132 32452 13188
rect 31948 13076 32004 13132
rect 31612 13020 32004 13076
rect 32396 13074 32452 13132
rect 32396 13022 32398 13074
rect 32450 13022 32452 13074
rect 31276 12402 31444 12404
rect 31276 12350 31278 12402
rect 31330 12350 31444 12402
rect 31276 12348 31444 12350
rect 31500 12850 31556 12862
rect 31500 12798 31502 12850
rect 31554 12798 31556 12850
rect 31276 12338 31332 12348
rect 31500 11284 31556 12798
rect 31612 12178 31668 13020
rect 32396 13010 32452 13022
rect 32060 12964 32116 12974
rect 32172 12964 32228 12974
rect 31948 12908 32060 12964
rect 32116 12962 32228 12964
rect 32116 12910 32174 12962
rect 32226 12910 32228 12962
rect 32116 12908 32228 12910
rect 31948 12852 32004 12908
rect 32060 12870 32116 12908
rect 32172 12898 32228 12908
rect 31836 12796 32004 12852
rect 31836 12290 31892 12796
rect 31836 12238 31838 12290
rect 31890 12238 31892 12290
rect 31836 12226 31892 12238
rect 31612 12126 31614 12178
rect 31666 12126 31668 12178
rect 31612 12114 31668 12126
rect 32620 11508 32676 15092
rect 33292 14644 33348 14654
rect 33292 14530 33348 14588
rect 33292 14478 33294 14530
rect 33346 14478 33348 14530
rect 33292 14466 33348 14478
rect 32732 14420 32788 14430
rect 32732 14326 32788 14364
rect 32284 11452 32676 11508
rect 32844 12850 32900 12862
rect 32844 12798 32846 12850
rect 32898 12798 32900 12850
rect 32284 11396 32340 11452
rect 32844 11396 32900 12798
rect 33180 12292 33236 12302
rect 33068 12290 33236 12292
rect 33068 12238 33182 12290
rect 33234 12238 33236 12290
rect 33068 12236 33236 12238
rect 32172 11394 32340 11396
rect 32172 11342 32286 11394
rect 32338 11342 32340 11394
rect 32172 11340 32340 11342
rect 31500 11228 31892 11284
rect 31164 10220 31444 10276
rect 31276 9938 31332 9950
rect 31276 9886 31278 9938
rect 31330 9886 31332 9938
rect 31276 9266 31332 9886
rect 31276 9214 31278 9266
rect 31330 9214 31332 9266
rect 31276 9202 31332 9214
rect 31388 9266 31444 10220
rect 31836 9938 31892 11228
rect 32172 10500 32228 11340
rect 32284 11330 32340 11340
rect 32396 11394 32900 11396
rect 32396 11342 32846 11394
rect 32898 11342 32900 11394
rect 32396 11340 32900 11342
rect 32396 11172 32452 11340
rect 32844 11330 32900 11340
rect 32956 11396 33012 11406
rect 33068 11396 33124 12236
rect 33180 12226 33236 12236
rect 33292 12178 33348 12190
rect 33292 12126 33294 12178
rect 33346 12126 33348 12178
rect 33012 11340 33124 11396
rect 33180 11954 33236 11966
rect 33180 11902 33182 11954
rect 33234 11902 33236 11954
rect 32956 11302 33012 11340
rect 32284 11116 32452 11172
rect 32284 10722 32340 11116
rect 33180 11060 33236 11902
rect 33292 11508 33348 12126
rect 33292 11442 33348 11452
rect 33292 11284 33348 11294
rect 33404 11284 33460 18396
rect 33628 17332 33684 18956
rect 34300 18564 34356 19966
rect 34524 19234 34580 19246
rect 34524 19182 34526 19234
rect 34578 19182 34580 19234
rect 34524 18564 34580 19182
rect 34636 18788 34692 26852
rect 34748 26628 34804 26638
rect 34748 23548 34804 26572
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35420 24724 35476 24734
rect 35420 24722 35588 24724
rect 35420 24670 35422 24722
rect 35474 24670 35588 24722
rect 35420 24668 35588 24670
rect 35420 24658 35476 24668
rect 34972 24610 35028 24622
rect 34972 24558 34974 24610
rect 35026 24558 35028 24610
rect 34748 23492 34916 23548
rect 34748 22930 34804 22942
rect 34748 22878 34750 22930
rect 34802 22878 34804 22930
rect 34748 20244 34804 22878
rect 34860 21028 34916 23492
rect 34972 23044 35028 24558
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 23938 35252 23950
rect 35196 23886 35198 23938
rect 35250 23886 35252 23938
rect 35196 23268 35252 23886
rect 35532 23268 35588 24668
rect 35196 23212 35476 23268
rect 34972 22978 35028 22988
rect 35308 23044 35364 23054
rect 35308 22950 35364 22988
rect 35420 22932 35476 23212
rect 35532 23174 35588 23212
rect 35420 22876 35588 22932
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34860 20972 35028 21028
rect 34748 20178 34804 20188
rect 34860 20356 34916 20366
rect 34748 19348 34804 19358
rect 34860 19348 34916 20300
rect 34748 19346 34916 19348
rect 34748 19294 34750 19346
rect 34802 19294 34916 19346
rect 34748 19292 34916 19294
rect 34748 19282 34804 19292
rect 34636 18732 34804 18788
rect 33852 18508 34580 18564
rect 33516 17276 33684 17332
rect 33740 18228 33796 18238
rect 33852 18228 33908 18508
rect 33964 18340 34020 18350
rect 34412 18340 34468 18350
rect 34748 18340 34804 18732
rect 33964 18338 34468 18340
rect 33964 18286 33966 18338
rect 34018 18286 34414 18338
rect 34466 18286 34468 18338
rect 33964 18284 34468 18286
rect 33964 18274 34020 18284
rect 33740 18226 33908 18228
rect 33740 18174 33742 18226
rect 33794 18174 33908 18226
rect 33740 18172 33908 18174
rect 34412 18226 34468 18284
rect 34412 18174 34414 18226
rect 34466 18174 34468 18226
rect 33516 16884 33572 17276
rect 33628 17108 33684 17118
rect 33628 17014 33684 17052
rect 33516 16828 33684 16884
rect 33292 11282 33460 11284
rect 33292 11230 33294 11282
rect 33346 11230 33460 11282
rect 33292 11228 33460 11230
rect 33292 11218 33348 11228
rect 33180 11004 33348 11060
rect 32284 10670 32286 10722
rect 32338 10670 32340 10722
rect 32284 10658 32340 10670
rect 32396 10722 32452 10734
rect 32396 10670 32398 10722
rect 32450 10670 32452 10722
rect 32396 10500 32452 10670
rect 32620 10724 32676 10734
rect 33180 10724 33236 10734
rect 32620 10722 33236 10724
rect 32620 10670 32622 10722
rect 32674 10670 33182 10722
rect 33234 10670 33236 10722
rect 32620 10668 33236 10670
rect 32620 10658 32676 10668
rect 33180 10658 33236 10668
rect 33292 10722 33348 11004
rect 33292 10670 33294 10722
rect 33346 10670 33348 10722
rect 33292 10658 33348 10670
rect 32172 10444 32452 10500
rect 31836 9886 31838 9938
rect 31890 9886 31892 9938
rect 31836 9874 31892 9886
rect 33180 10386 33236 10398
rect 33180 10334 33182 10386
rect 33234 10334 33236 10386
rect 31388 9214 31390 9266
rect 31442 9214 31444 9266
rect 31164 9156 31220 9166
rect 31164 9062 31220 9100
rect 31388 8428 31444 9214
rect 31724 9602 31780 9614
rect 31724 9550 31726 9602
rect 31778 9550 31780 9602
rect 31724 9156 31780 9550
rect 30940 8372 31332 8428
rect 31388 8372 31556 8428
rect 31276 7700 31332 8372
rect 31500 8258 31556 8372
rect 31724 8370 31780 9100
rect 31724 8318 31726 8370
rect 31778 8318 31780 8370
rect 31724 8306 31780 8318
rect 31836 9042 31892 9054
rect 31836 8990 31838 9042
rect 31890 8990 31892 9042
rect 31500 8206 31502 8258
rect 31554 8206 31556 8258
rect 31500 8194 31556 8206
rect 31276 7644 31780 7700
rect 31612 7476 31668 7486
rect 31276 6692 31332 6702
rect 31276 6598 31332 6636
rect 31612 6690 31668 7420
rect 31612 6638 31614 6690
rect 31666 6638 31668 6690
rect 31612 6626 31668 6638
rect 31724 6692 31780 7644
rect 31836 7698 31892 8990
rect 31836 7646 31838 7698
rect 31890 7646 31892 7698
rect 31836 7634 31892 7646
rect 32172 8146 32228 8158
rect 32172 8094 32174 8146
rect 32226 8094 32228 8146
rect 32060 7588 32116 7598
rect 31948 7586 32116 7588
rect 31948 7534 32062 7586
rect 32114 7534 32116 7586
rect 31948 7532 32116 7534
rect 31836 6692 31892 6702
rect 31724 6690 31892 6692
rect 31724 6638 31838 6690
rect 31890 6638 31892 6690
rect 31724 6636 31892 6638
rect 31836 6626 31892 6636
rect 31388 6580 31444 6590
rect 31388 6486 31444 6524
rect 31948 5906 32004 7532
rect 32060 7522 32116 7532
rect 31948 5854 31950 5906
rect 32002 5854 32004 5906
rect 30604 5030 30660 5068
rect 31500 5122 31556 5134
rect 31500 5070 31502 5122
rect 31554 5070 31556 5122
rect 30380 4958 30382 5010
rect 30434 4958 30436 5010
rect 30380 4946 30436 4958
rect 30492 4452 30548 4462
rect 30492 4358 30548 4396
rect 30604 4340 30660 4350
rect 30604 4246 30660 4284
rect 31500 4340 31556 5070
rect 31948 4898 32004 5854
rect 32172 7474 32228 8094
rect 32172 7422 32174 7474
rect 32226 7422 32228 7474
rect 32172 5794 32228 7422
rect 32956 7476 33012 7486
rect 32956 7382 33012 7420
rect 32396 6692 32452 6702
rect 32396 6020 32452 6636
rect 33180 6580 33236 10334
rect 33628 9940 33684 16828
rect 33740 14308 33796 18172
rect 34412 18162 34468 18174
rect 34524 18284 34804 18340
rect 34524 17778 34580 18284
rect 34524 17726 34526 17778
rect 34578 17726 34580 17778
rect 34188 17108 34244 17118
rect 34188 17014 34244 17052
rect 34524 16996 34580 17726
rect 34748 17668 34804 18284
rect 34860 18674 34916 19292
rect 34860 18622 34862 18674
rect 34914 18622 34916 18674
rect 34860 18226 34916 18622
rect 34860 18174 34862 18226
rect 34914 18174 34916 18226
rect 34860 18162 34916 18174
rect 34860 17668 34916 17678
rect 34748 17666 34916 17668
rect 34748 17614 34862 17666
rect 34914 17614 34916 17666
rect 34748 17612 34916 17614
rect 34860 17602 34916 17612
rect 34524 16930 34580 16940
rect 34972 14644 35028 20972
rect 35196 20356 35252 20366
rect 35084 20130 35140 20142
rect 35084 20078 35086 20130
rect 35138 20078 35140 20130
rect 35084 19908 35140 20078
rect 35196 20018 35252 20300
rect 35196 19966 35198 20018
rect 35250 19966 35252 20018
rect 35196 19954 35252 19966
rect 35084 19236 35140 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19460 35588 22876
rect 35308 19404 35588 19460
rect 35308 19346 35364 19404
rect 35756 19348 35812 26852
rect 35868 24612 35924 24622
rect 35868 24518 35924 24556
rect 36092 24050 36148 26852
rect 36092 23998 36094 24050
rect 36146 23998 36148 24050
rect 36092 23986 36148 23998
rect 36092 20578 36148 20590
rect 36092 20526 36094 20578
rect 36146 20526 36148 20578
rect 36092 20356 36148 20526
rect 36092 20290 36148 20300
rect 36428 20244 36484 20254
rect 36428 20130 36484 20188
rect 36428 20078 36430 20130
rect 36482 20078 36484 20130
rect 36428 20066 36484 20078
rect 36204 20020 36260 20030
rect 35308 19294 35310 19346
rect 35362 19294 35364 19346
rect 35308 19282 35364 19294
rect 35420 19292 35812 19348
rect 36092 20018 36260 20020
rect 36092 19966 36206 20018
rect 36258 19966 36260 20018
rect 36092 19964 36260 19966
rect 35084 19170 35140 19180
rect 35420 18228 35476 19292
rect 35980 19236 36036 19246
rect 35532 19180 35980 19236
rect 35532 18450 35588 19180
rect 35980 19142 36036 19180
rect 36092 18674 36148 19964
rect 36204 19954 36260 19964
rect 36316 19908 36372 19918
rect 36316 19814 36372 19852
rect 36652 19908 36708 19918
rect 36092 18622 36094 18674
rect 36146 18622 36148 18674
rect 36092 18610 36148 18622
rect 36204 19348 36260 19358
rect 35532 18398 35534 18450
rect 35586 18398 35588 18450
rect 35532 18386 35588 18398
rect 35756 18452 35812 18462
rect 36204 18452 36260 19292
rect 36316 19236 36372 19246
rect 36316 18674 36372 19180
rect 36316 18622 36318 18674
rect 36370 18622 36372 18674
rect 36316 18610 36372 18622
rect 35756 18450 36260 18452
rect 35756 18398 35758 18450
rect 35810 18398 36260 18450
rect 35756 18396 36260 18398
rect 36540 18562 36596 18574
rect 36540 18510 36542 18562
rect 36594 18510 36596 18562
rect 36540 18452 36596 18510
rect 36652 18564 36708 19852
rect 36652 18470 36708 18508
rect 35756 18386 35812 18396
rect 35420 18172 35588 18228
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17780 35476 17790
rect 35532 17780 35588 18172
rect 36092 17890 36148 18396
rect 36540 18386 36596 18396
rect 36092 17838 36094 17890
rect 36146 17838 36148 17890
rect 36092 17826 36148 17838
rect 35420 17778 35700 17780
rect 35420 17726 35422 17778
rect 35474 17726 35700 17778
rect 35420 17724 35700 17726
rect 35420 17714 35476 17724
rect 35644 16772 35700 17724
rect 36204 17556 36260 17566
rect 36092 17444 36148 17454
rect 35980 17442 36148 17444
rect 35980 17390 36094 17442
rect 36146 17390 36148 17442
rect 35980 17388 36148 17390
rect 35980 16996 36036 17388
rect 36092 17378 36148 17388
rect 36204 17108 36260 17500
rect 36540 17108 36596 17118
rect 36204 17106 36596 17108
rect 36204 17054 36542 17106
rect 36594 17054 36596 17106
rect 36204 17052 36596 17054
rect 36540 17042 36596 17052
rect 35980 16930 36036 16940
rect 35644 16716 36260 16772
rect 35980 16548 36036 16558
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 15428 35364 15438
rect 35756 15428 35812 15438
rect 35308 15426 35812 15428
rect 35308 15374 35310 15426
rect 35362 15374 35758 15426
rect 35810 15374 35812 15426
rect 35308 15372 35812 15374
rect 35308 15148 35364 15372
rect 35756 15362 35812 15372
rect 35980 15426 36036 16492
rect 36204 16212 36260 16716
rect 36764 16212 36820 38612
rect 37212 35474 37268 35486
rect 37212 35422 37214 35474
rect 37266 35422 37268 35474
rect 37100 34692 37156 34702
rect 37100 34598 37156 34636
rect 36876 34130 36932 34142
rect 36876 34078 36878 34130
rect 36930 34078 36932 34130
rect 36876 33572 36932 34078
rect 36876 33516 37156 33572
rect 37100 33460 37156 33516
rect 37100 33366 37156 33404
rect 37212 33124 37268 35422
rect 37436 35476 37492 35486
rect 37436 33346 37492 35420
rect 37548 34020 37604 38612
rect 37772 40178 37940 40180
rect 37772 40126 37886 40178
rect 37938 40126 37940 40178
rect 37772 40124 37940 40126
rect 37772 35588 37828 40124
rect 37884 40114 37940 40124
rect 37996 39956 38052 43708
rect 38108 43538 38164 44268
rect 38444 44258 38500 44268
rect 38556 44100 38612 48076
rect 38780 47460 38836 48972
rect 39116 48804 39172 48814
rect 38668 47404 38836 47460
rect 39004 47572 39060 47582
rect 38668 45444 38724 47404
rect 38892 47348 38948 47358
rect 38780 47234 38836 47246
rect 38780 47182 38782 47234
rect 38834 47182 38836 47234
rect 38780 47124 38836 47182
rect 38780 47058 38836 47068
rect 38668 45378 38724 45388
rect 38668 45106 38724 45118
rect 38668 45054 38670 45106
rect 38722 45054 38724 45106
rect 38668 44996 38724 45054
rect 38668 44930 38724 44940
rect 38668 44660 38724 44670
rect 38724 44604 38836 44660
rect 38668 44594 38724 44604
rect 38668 44324 38724 44334
rect 38668 44230 38724 44268
rect 38108 43486 38110 43538
rect 38162 43486 38164 43538
rect 38108 43474 38164 43486
rect 38220 44044 38612 44100
rect 38108 42866 38164 42878
rect 38108 42814 38110 42866
rect 38162 42814 38164 42866
rect 38108 42532 38164 42814
rect 38108 42466 38164 42476
rect 38108 42084 38164 42094
rect 38220 42084 38276 44044
rect 38780 43540 38836 44604
rect 38556 43484 38836 43540
rect 38444 43316 38500 43326
rect 38108 42082 38276 42084
rect 38108 42030 38110 42082
rect 38162 42030 38276 42082
rect 38108 42028 38276 42030
rect 38332 43314 38500 43316
rect 38332 43262 38446 43314
rect 38498 43262 38500 43314
rect 38332 43260 38500 43262
rect 38108 42018 38164 42028
rect 38220 41298 38276 41310
rect 38220 41246 38222 41298
rect 38274 41246 38276 41298
rect 38220 40292 38276 41246
rect 38220 40226 38276 40236
rect 37884 39900 38052 39956
rect 37884 36708 37940 39900
rect 37996 39394 38052 39406
rect 37996 39342 37998 39394
rect 38050 39342 38052 39394
rect 37996 38836 38052 39342
rect 37996 38770 38052 38780
rect 38332 38668 38388 43260
rect 38444 43250 38500 43260
rect 38444 42756 38500 42766
rect 38556 42756 38612 43484
rect 38444 42754 38612 42756
rect 38444 42702 38446 42754
rect 38498 42702 38612 42754
rect 38444 42700 38612 42702
rect 38668 43316 38724 43326
rect 38444 42084 38500 42700
rect 38444 42018 38500 42028
rect 38556 41860 38612 41870
rect 38556 41186 38612 41804
rect 38556 41134 38558 41186
rect 38610 41134 38612 41186
rect 38556 40964 38612 41134
rect 38556 40898 38612 40908
rect 38668 40626 38724 43260
rect 38892 41188 38948 47292
rect 39004 43428 39060 47516
rect 39004 43362 39060 43372
rect 39004 42532 39060 42542
rect 39004 42438 39060 42476
rect 39116 41188 39172 48748
rect 39228 46004 39284 48972
rect 39340 48468 39396 48478
rect 39340 47348 39396 48412
rect 39340 47282 39396 47292
rect 39228 45938 39284 45948
rect 39340 45220 39396 45230
rect 39452 45220 39508 50652
rect 39564 49924 39620 49934
rect 39620 49868 39732 49924
rect 39564 49830 39620 49868
rect 39676 49140 39732 49868
rect 39676 49074 39732 49084
rect 39564 49028 39620 49038
rect 39564 48914 39620 48972
rect 39564 48862 39566 48914
rect 39618 48862 39620 48914
rect 39564 48850 39620 48862
rect 39564 48356 39620 48366
rect 39564 48242 39620 48300
rect 39564 48190 39566 48242
rect 39618 48190 39620 48242
rect 39564 47124 39620 48190
rect 39788 47460 39844 56140
rect 39900 50034 39956 58156
rect 40012 58118 40068 58156
rect 40124 57538 40180 57550
rect 40124 57486 40126 57538
rect 40178 57486 40180 57538
rect 40124 56196 40180 57486
rect 40124 56130 40180 56140
rect 40012 54514 40068 54526
rect 40012 54462 40014 54514
rect 40066 54462 40068 54514
rect 40012 54180 40068 54462
rect 40012 54114 40068 54124
rect 40348 53172 40404 60508
rect 40684 60340 40740 60350
rect 41244 60340 41300 60844
rect 41356 60834 41412 60844
rect 41468 60788 41524 60798
rect 41468 60564 41524 60732
rect 41580 60676 41636 62302
rect 41692 62356 41748 62366
rect 41692 62262 41748 62300
rect 41804 62354 41860 62366
rect 41804 62302 41806 62354
rect 41858 62302 41860 62354
rect 41804 62188 41860 62302
rect 42252 62354 42308 62366
rect 42252 62302 42254 62354
rect 42306 62302 42308 62354
rect 42252 62188 42308 62302
rect 42924 62356 42980 62366
rect 42924 62262 42980 62300
rect 41804 62132 42084 62188
rect 42252 62132 42868 62188
rect 41916 61684 41972 61694
rect 41916 61012 41972 61628
rect 41916 60918 41972 60956
rect 42028 61570 42084 62132
rect 42476 61684 42532 61694
rect 42476 61590 42532 61628
rect 42028 61518 42030 61570
rect 42082 61518 42084 61570
rect 41804 60676 41860 60686
rect 41580 60674 41860 60676
rect 41580 60622 41806 60674
rect 41858 60622 41860 60674
rect 41580 60620 41860 60622
rect 41804 60610 41860 60620
rect 42028 60564 42084 61518
rect 41468 60508 41748 60564
rect 40684 60226 40740 60284
rect 40684 60174 40686 60226
rect 40738 60174 40740 60226
rect 40684 60162 40740 60174
rect 41020 60284 41300 60340
rect 41020 60226 41076 60284
rect 41020 60174 41022 60226
rect 41074 60174 41076 60226
rect 41020 60162 41076 60174
rect 40460 60116 40516 60126
rect 40460 60022 40516 60060
rect 41132 58324 41188 58334
rect 40572 58212 40628 58222
rect 40572 58118 40628 58156
rect 41132 58210 41188 58268
rect 41132 58158 41134 58210
rect 41186 58158 41188 58210
rect 40460 56868 40516 56878
rect 40796 56868 40852 56878
rect 40460 56866 40740 56868
rect 40460 56814 40462 56866
rect 40514 56814 40740 56866
rect 40460 56812 40740 56814
rect 40460 56802 40516 56812
rect 40684 55300 40740 56812
rect 40796 56774 40852 56812
rect 41132 56420 41188 58158
rect 41468 56868 41524 56878
rect 40908 56364 41188 56420
rect 41244 56866 41524 56868
rect 41244 56814 41470 56866
rect 41522 56814 41524 56866
rect 41244 56812 41524 56814
rect 40908 56082 40964 56364
rect 41244 56306 41300 56812
rect 41468 56802 41524 56812
rect 41244 56254 41246 56306
rect 41298 56254 41300 56306
rect 41244 56242 41300 56254
rect 41020 56196 41076 56206
rect 41020 56102 41076 56140
rect 40908 56030 40910 56082
rect 40962 56030 40964 56082
rect 40908 55972 40964 56030
rect 40908 55906 40964 55916
rect 41580 55972 41636 55982
rect 41580 55878 41636 55916
rect 40796 55300 40852 55310
rect 40684 55298 40852 55300
rect 40684 55246 40798 55298
rect 40850 55246 40852 55298
rect 40684 55244 40852 55246
rect 40572 55074 40628 55086
rect 40572 55022 40574 55074
rect 40626 55022 40628 55074
rect 40460 53172 40516 53182
rect 40348 53170 40516 53172
rect 40348 53118 40462 53170
rect 40514 53118 40516 53170
rect 40348 53116 40516 53118
rect 40460 53106 40516 53116
rect 40236 53060 40292 53070
rect 40236 52966 40292 53004
rect 40124 52948 40180 52958
rect 40012 52946 40180 52948
rect 40012 52894 40126 52946
rect 40178 52894 40180 52946
rect 40012 52892 40180 52894
rect 40012 51604 40068 52892
rect 40124 52882 40180 52892
rect 40012 51538 40068 51548
rect 40348 52274 40404 52286
rect 40348 52222 40350 52274
rect 40402 52222 40404 52274
rect 40348 50820 40404 52222
rect 40348 50754 40404 50764
rect 39900 49982 39902 50034
rect 39954 49982 39956 50034
rect 39900 47572 39956 49982
rect 40124 49812 40180 49822
rect 40012 49810 40180 49812
rect 40012 49758 40126 49810
rect 40178 49758 40180 49810
rect 40012 49756 40180 49758
rect 40012 49028 40068 49756
rect 40124 49746 40180 49756
rect 40460 49140 40516 49150
rect 40572 49140 40628 55022
rect 40684 55076 40740 55086
rect 40684 54982 40740 55020
rect 40796 54738 40852 55244
rect 41020 55076 41076 55086
rect 40796 54686 40798 54738
rect 40850 54686 40852 54738
rect 40796 54674 40852 54686
rect 40908 55074 41076 55076
rect 40908 55022 41022 55074
rect 41074 55022 41076 55074
rect 40908 55020 41076 55022
rect 40796 54404 40852 54414
rect 40684 53844 40740 53854
rect 40684 53750 40740 53788
rect 40796 52388 40852 54348
rect 40908 52948 40964 55020
rect 41020 55010 41076 55020
rect 41692 54740 41748 60508
rect 42028 60498 42084 60508
rect 42140 61572 42196 61582
rect 42140 60562 42196 61516
rect 42812 61570 42868 62132
rect 42812 61518 42814 61570
rect 42866 61518 42868 61570
rect 42812 61506 42868 61518
rect 43036 61684 43092 61694
rect 43036 61458 43092 61628
rect 43148 61572 43204 61582
rect 43148 61478 43204 61516
rect 43036 61406 43038 61458
rect 43090 61406 43092 61458
rect 43036 61394 43092 61406
rect 42140 60510 42142 60562
rect 42194 60510 42196 60562
rect 41916 59444 41972 59454
rect 41916 57092 41972 59388
rect 41916 57026 41972 57036
rect 42140 57090 42196 60510
rect 43260 59332 43316 62412
rect 43708 62354 43764 62366
rect 43708 62302 43710 62354
rect 43762 62302 43764 62354
rect 43372 62244 43428 62254
rect 43708 62244 43764 62302
rect 43372 62242 43764 62244
rect 43372 62190 43374 62242
rect 43426 62190 43764 62242
rect 43372 62188 43764 62190
rect 43372 62178 43428 62188
rect 43260 59266 43316 59276
rect 43596 58546 43652 62188
rect 43932 61460 43988 63086
rect 44044 62580 44100 63198
rect 44044 62514 44100 62524
rect 44268 62916 44324 62926
rect 44044 62356 44100 62366
rect 44044 62262 44100 62300
rect 44268 62354 44324 62860
rect 44268 62302 44270 62354
rect 44322 62302 44324 62354
rect 44268 62290 44324 62302
rect 43932 61394 43988 61404
rect 44492 58828 44548 67172
rect 44604 67060 44660 67098
rect 44604 66994 44660 67004
rect 44940 63922 44996 63934
rect 44940 63870 44942 63922
rect 44994 63870 44996 63922
rect 44940 63140 44996 63870
rect 45948 63922 46004 63934
rect 45948 63870 45950 63922
rect 46002 63870 46004 63922
rect 45836 63812 45892 63822
rect 45836 63718 45892 63756
rect 45948 63364 46004 63870
rect 45500 63308 46004 63364
rect 44940 63074 44996 63084
rect 45388 63140 45444 63150
rect 45500 63140 45556 63308
rect 45948 63252 46004 63308
rect 45948 63186 46004 63196
rect 46060 63812 46116 63822
rect 45388 63138 45556 63140
rect 45388 63086 45390 63138
rect 45442 63086 45556 63138
rect 45388 63084 45556 63086
rect 45612 63140 45668 63150
rect 44604 62580 44660 62590
rect 45276 62580 45332 62590
rect 45388 62580 45444 63084
rect 45612 63046 45668 63084
rect 45948 62916 46004 62926
rect 44660 62524 44996 62580
rect 44604 62514 44660 62524
rect 44940 62354 44996 62524
rect 45276 62578 45444 62580
rect 45276 62526 45278 62578
rect 45330 62526 45444 62578
rect 45276 62524 45444 62526
rect 45724 62914 46004 62916
rect 45724 62862 45950 62914
rect 46002 62862 46004 62914
rect 45724 62860 46004 62862
rect 45724 62578 45780 62860
rect 45948 62850 46004 62860
rect 45724 62526 45726 62578
rect 45778 62526 45780 62578
rect 45276 62514 45332 62524
rect 45724 62514 45780 62526
rect 45948 62580 46004 62590
rect 46060 62580 46116 63756
rect 46844 63252 46900 63262
rect 46844 63158 46900 63196
rect 46620 63140 46676 63150
rect 45948 62578 46116 62580
rect 45948 62526 45950 62578
rect 46002 62526 46116 62578
rect 45948 62524 46116 62526
rect 46284 62914 46340 62926
rect 46284 62862 46286 62914
rect 46338 62862 46340 62914
rect 45948 62514 46004 62524
rect 44940 62302 44942 62354
rect 44994 62302 44996 62354
rect 44940 62290 44996 62302
rect 46284 62354 46340 62862
rect 46284 62302 46286 62354
rect 46338 62302 46340 62354
rect 46284 62290 46340 62302
rect 44716 62242 44772 62254
rect 44716 62190 44718 62242
rect 44770 62190 44772 62242
rect 44716 61796 44772 62190
rect 45836 62242 45892 62254
rect 45836 62190 45838 62242
rect 45890 62190 45892 62242
rect 45836 62188 45892 62190
rect 46620 62188 46676 63084
rect 45836 62132 46340 62188
rect 46620 62132 46788 62188
rect 44828 61796 44884 61806
rect 44716 61794 44884 61796
rect 44716 61742 44830 61794
rect 44882 61742 44884 61794
rect 44716 61740 44884 61742
rect 44828 61730 44884 61740
rect 44940 61460 44996 61470
rect 44492 58772 44660 58828
rect 43596 58494 43598 58546
rect 43650 58494 43652 58546
rect 43596 58482 43652 58494
rect 43148 58434 43204 58446
rect 43148 58382 43150 58434
rect 43202 58382 43204 58434
rect 42140 57038 42142 57090
rect 42194 57038 42196 57090
rect 42140 57026 42196 57038
rect 42924 57650 42980 57662
rect 42924 57598 42926 57650
rect 42978 57598 42980 57650
rect 42924 56532 42980 57598
rect 43036 57538 43092 57550
rect 43036 57486 43038 57538
rect 43090 57486 43092 57538
rect 43036 56756 43092 57486
rect 43148 56868 43204 58382
rect 43484 58434 43540 58446
rect 43484 58382 43486 58434
rect 43538 58382 43540 58434
rect 43372 58212 43428 58222
rect 43204 56812 43316 56868
rect 43148 56802 43204 56812
rect 43036 56662 43092 56700
rect 43148 56642 43204 56654
rect 43148 56590 43150 56642
rect 43202 56590 43204 56642
rect 43148 56532 43204 56590
rect 42924 56476 43204 56532
rect 42028 56196 42084 56206
rect 42028 56102 42084 56140
rect 41692 54674 41748 54684
rect 42140 55524 42196 55534
rect 41020 54626 41076 54638
rect 41020 54574 41022 54626
rect 41074 54574 41076 54626
rect 41020 54404 41076 54574
rect 42028 54628 42084 54638
rect 41020 54338 41076 54348
rect 41132 54514 41188 54526
rect 41132 54462 41134 54514
rect 41186 54462 41188 54514
rect 41132 53954 41188 54462
rect 41692 54404 41748 54414
rect 41132 53902 41134 53954
rect 41186 53902 41188 53954
rect 41132 53890 41188 53902
rect 41244 54180 41300 54190
rect 41244 53844 41300 54124
rect 41244 53788 41412 53844
rect 41356 53730 41412 53788
rect 41356 53678 41358 53730
rect 41410 53678 41412 53730
rect 41356 53666 41412 53678
rect 41692 53730 41748 54348
rect 42028 53956 42084 54572
rect 42140 54180 42196 55468
rect 43148 55076 43204 56476
rect 43148 55010 43204 55020
rect 43036 54628 43092 54638
rect 42812 54572 43036 54628
rect 42812 54516 42868 54572
rect 43036 54562 43092 54572
rect 43260 54626 43316 56812
rect 43372 56866 43428 58156
rect 43372 56814 43374 56866
rect 43426 56814 43428 56866
rect 43372 56802 43428 56814
rect 43484 57762 43540 58382
rect 43484 57710 43486 57762
rect 43538 57710 43540 57762
rect 43484 56868 43540 57710
rect 43932 58322 43988 58334
rect 43932 58270 43934 58322
rect 43986 58270 43988 58322
rect 43596 56868 43652 56878
rect 43484 56866 43652 56868
rect 43484 56814 43598 56866
rect 43650 56814 43652 56866
rect 43484 56812 43652 56814
rect 43596 56802 43652 56812
rect 43708 56868 43764 56878
rect 43708 56754 43764 56812
rect 43932 56866 43988 58270
rect 44044 58212 44100 58222
rect 44044 58118 44100 58156
rect 44268 58212 44324 58222
rect 44268 58210 44548 58212
rect 44268 58158 44270 58210
rect 44322 58158 44548 58210
rect 44268 58156 44548 58158
rect 44268 58146 44324 58156
rect 44492 57876 44548 58156
rect 44492 57650 44548 57820
rect 44492 57598 44494 57650
rect 44546 57598 44548 57650
rect 44492 57586 44548 57598
rect 44604 57652 44660 58772
rect 44828 58548 44884 58558
rect 44940 58548 44996 61404
rect 45836 59332 45892 59342
rect 45836 59238 45892 59276
rect 46284 59220 46340 62132
rect 46284 59218 46564 59220
rect 46284 59166 46286 59218
rect 46338 59166 46564 59218
rect 46284 59164 46564 59166
rect 46284 59154 46340 59164
rect 46172 59106 46228 59118
rect 46172 59054 46174 59106
rect 46226 59054 46228 59106
rect 44828 58546 44996 58548
rect 44828 58494 44830 58546
rect 44882 58494 44996 58546
rect 44828 58492 44996 58494
rect 45164 58546 45220 58558
rect 45164 58494 45166 58546
rect 45218 58494 45220 58546
rect 44828 58482 44884 58492
rect 45164 57764 45220 58494
rect 44604 57586 44660 57596
rect 44828 57762 45220 57764
rect 44828 57710 45166 57762
rect 45218 57710 45220 57762
rect 44828 57708 45220 57710
rect 44268 57540 44324 57550
rect 43932 56814 43934 56866
rect 43986 56814 43988 56866
rect 43932 56802 43988 56814
rect 44156 57484 44268 57540
rect 43708 56702 43710 56754
rect 43762 56702 43764 56754
rect 43708 56690 43764 56702
rect 43596 56644 43652 56654
rect 43260 54574 43262 54626
rect 43314 54574 43316 54626
rect 43260 54562 43316 54574
rect 43484 55188 43540 55198
rect 42140 54114 42196 54124
rect 42252 54514 42868 54516
rect 42252 54462 42814 54514
rect 42866 54462 42868 54514
rect 42252 54460 42868 54462
rect 42028 53900 42196 53956
rect 41916 53844 41972 53854
rect 41916 53732 41972 53788
rect 41692 53678 41694 53730
rect 41746 53678 41748 53730
rect 41692 53666 41748 53678
rect 41804 53730 41972 53732
rect 41804 53678 41918 53730
rect 41970 53678 41972 53730
rect 41804 53676 41972 53678
rect 41132 53620 41188 53630
rect 41132 53506 41188 53564
rect 41132 53454 41134 53506
rect 41186 53454 41188 53506
rect 41468 53620 41524 53630
rect 41468 53562 41524 53564
rect 41468 53510 41470 53562
rect 41522 53510 41524 53562
rect 41468 53498 41524 53510
rect 41132 53396 41188 53454
rect 40908 52882 40964 52892
rect 41020 53284 41076 53294
rect 41020 52946 41076 53228
rect 41020 52894 41022 52946
rect 41074 52894 41076 52946
rect 41020 52882 41076 52894
rect 41132 52388 41188 53340
rect 40796 52332 40964 52388
rect 40908 51602 40964 52332
rect 41132 52322 41188 52332
rect 41244 53060 41300 53070
rect 41020 52276 41076 52286
rect 41020 52162 41076 52220
rect 41244 52276 41300 53004
rect 41804 53058 41860 53676
rect 41916 53666 41972 53676
rect 42140 53620 42196 53900
rect 42252 53730 42308 54460
rect 42812 54450 42868 54460
rect 43148 54514 43204 54526
rect 43148 54462 43150 54514
rect 43202 54462 43204 54514
rect 43148 54404 43204 54462
rect 43148 54338 43204 54348
rect 42924 54068 42980 54078
rect 42252 53678 42254 53730
rect 42306 53678 42308 53730
rect 42252 53666 42308 53678
rect 42700 53730 42756 53742
rect 42700 53678 42702 53730
rect 42754 53678 42756 53730
rect 42140 53554 42196 53564
rect 42028 53506 42084 53518
rect 42028 53454 42030 53506
rect 42082 53454 42084 53506
rect 41916 53396 41972 53406
rect 41916 53170 41972 53340
rect 42028 53284 42084 53454
rect 42364 53396 42420 53406
rect 42084 53228 42308 53284
rect 42028 53218 42084 53228
rect 41916 53118 41918 53170
rect 41970 53118 41972 53170
rect 41916 53106 41972 53118
rect 41804 53006 41806 53058
rect 41858 53006 41860 53058
rect 41804 52994 41860 53006
rect 42140 52948 42196 52958
rect 42028 52946 42196 52948
rect 42028 52894 42142 52946
rect 42194 52894 42196 52946
rect 42028 52892 42196 52894
rect 41804 52724 41860 52734
rect 41692 52388 41748 52398
rect 41692 52294 41748 52332
rect 41244 52210 41300 52220
rect 41020 52110 41022 52162
rect 41074 52110 41076 52162
rect 41020 52098 41076 52110
rect 41804 52164 41860 52668
rect 41804 52050 41860 52108
rect 41804 51998 41806 52050
rect 41858 51998 41860 52050
rect 41804 51986 41860 51998
rect 41916 52276 41972 52286
rect 40908 51550 40910 51602
rect 40962 51550 40964 51602
rect 40908 51380 40964 51550
rect 40460 49138 40628 49140
rect 40460 49086 40462 49138
rect 40514 49086 40628 49138
rect 40460 49084 40628 49086
rect 40684 51324 40964 51380
rect 41020 51940 41076 51950
rect 40460 49074 40516 49084
rect 40012 48962 40068 48972
rect 40124 48916 40180 48926
rect 40180 48860 40292 48916
rect 40124 48822 40180 48860
rect 39900 47506 39956 47516
rect 40012 48804 40068 48814
rect 39788 47394 39844 47404
rect 39900 47346 39956 47358
rect 39900 47294 39902 47346
rect 39954 47294 39956 47346
rect 39676 47236 39732 47246
rect 39900 47236 39956 47294
rect 40012 47346 40068 48748
rect 40124 48132 40180 48142
rect 40124 48038 40180 48076
rect 40236 47908 40292 48860
rect 40012 47294 40014 47346
rect 40066 47294 40068 47346
rect 40012 47282 40068 47294
rect 40124 47852 40292 47908
rect 40348 48802 40404 48814
rect 40348 48750 40350 48802
rect 40402 48750 40404 48802
rect 39732 47180 39956 47236
rect 39676 47142 39732 47180
rect 39564 47058 39620 47068
rect 40124 46788 40180 47852
rect 40236 47684 40292 47694
rect 40236 47458 40292 47628
rect 40348 47572 40404 48750
rect 40460 48802 40516 48814
rect 40460 48750 40462 48802
rect 40514 48750 40516 48802
rect 40460 48356 40516 48750
rect 40684 48804 40740 51324
rect 40908 51156 40964 51166
rect 40796 51100 40908 51156
rect 40796 49138 40852 51100
rect 40908 51090 40964 51100
rect 41020 50428 41076 51884
rect 41692 51938 41748 51950
rect 41692 51886 41694 51938
rect 41746 51886 41748 51938
rect 41132 51716 41188 51726
rect 41132 51268 41188 51660
rect 41244 51492 41300 51502
rect 41692 51492 41748 51886
rect 41244 51490 41748 51492
rect 41244 51438 41246 51490
rect 41298 51438 41748 51490
rect 41244 51436 41748 51438
rect 41244 51426 41300 51436
rect 41132 51212 41300 51268
rect 40908 50372 41076 50428
rect 40908 50036 40964 50372
rect 40908 49922 40964 49980
rect 40908 49870 40910 49922
rect 40962 49870 40964 49922
rect 40908 49858 40964 49870
rect 41020 49924 41076 49934
rect 41020 49830 41076 49868
rect 41020 49588 41076 49598
rect 41020 49494 41076 49532
rect 40796 49086 40798 49138
rect 40850 49086 40852 49138
rect 40796 49074 40852 49086
rect 41132 49028 41188 49038
rect 40908 48916 40964 48926
rect 40684 48738 40740 48748
rect 40796 48914 40964 48916
rect 40796 48862 40910 48914
rect 40962 48862 40964 48914
rect 40796 48860 40964 48862
rect 40460 48290 40516 48300
rect 40796 47572 40852 48860
rect 40908 48850 40964 48860
rect 41132 48802 41188 48972
rect 41132 48750 41134 48802
rect 41186 48750 41188 48802
rect 41020 48468 41076 48478
rect 41132 48468 41188 48750
rect 41020 48466 41188 48468
rect 41020 48414 41022 48466
rect 41074 48414 41188 48466
rect 41020 48412 41188 48414
rect 41244 48466 41300 51212
rect 41244 48414 41246 48466
rect 41298 48414 41300 48466
rect 41020 48402 41076 48412
rect 41244 48402 41300 48414
rect 41356 48802 41412 48814
rect 41356 48750 41358 48802
rect 41410 48750 41412 48802
rect 41356 48356 41412 48750
rect 41356 48290 41412 48300
rect 40348 47516 40852 47572
rect 40908 48242 40964 48254
rect 40908 48190 40910 48242
rect 40962 48190 40964 48242
rect 40236 47406 40238 47458
rect 40290 47406 40292 47458
rect 40236 47394 40292 47406
rect 40460 47348 40516 47358
rect 40348 47292 40460 47348
rect 40012 46732 40180 46788
rect 40236 47236 40292 47246
rect 39900 46004 39956 46014
rect 39900 45910 39956 45948
rect 39900 45220 39956 45230
rect 39452 45164 39844 45220
rect 39340 45108 39396 45164
rect 39340 45052 39620 45108
rect 39564 44994 39620 45052
rect 39564 44942 39566 44994
rect 39618 44942 39620 44994
rect 39564 44930 39620 44942
rect 39676 44996 39732 45006
rect 39676 44324 39732 44940
rect 39452 44322 39732 44324
rect 39452 44270 39678 44322
rect 39730 44270 39732 44322
rect 39452 44268 39732 44270
rect 39340 44212 39396 44222
rect 38892 41122 38948 41132
rect 39004 41132 39172 41188
rect 39228 44210 39396 44212
rect 39228 44158 39342 44210
rect 39394 44158 39396 44210
rect 39228 44156 39396 44158
rect 38668 40574 38670 40626
rect 38722 40574 38724 40626
rect 38556 40402 38612 40414
rect 38556 40350 38558 40402
rect 38610 40350 38612 40402
rect 38556 40292 38612 40350
rect 38444 40236 38556 40292
rect 38444 39730 38500 40236
rect 38556 40226 38612 40236
rect 38444 39678 38446 39730
rect 38498 39678 38500 39730
rect 38444 39666 38500 39678
rect 38668 38836 38724 40574
rect 38892 40404 38948 40414
rect 38892 40310 38948 40348
rect 38892 39842 38948 39854
rect 38892 39790 38894 39842
rect 38946 39790 38948 39842
rect 38892 39730 38948 39790
rect 38892 39678 38894 39730
rect 38946 39678 38948 39730
rect 38892 39666 38948 39678
rect 38668 38770 38724 38780
rect 37884 36642 37940 36652
rect 37996 38612 38388 38668
rect 37772 34916 37828 35532
rect 37772 34822 37828 34860
rect 37884 36372 37940 36382
rect 37772 34132 37828 34142
rect 37884 34132 37940 36316
rect 37996 35924 38052 38612
rect 39004 38388 39060 41132
rect 39116 40964 39172 40974
rect 39116 40870 39172 40908
rect 39116 40628 39172 40638
rect 39116 40534 39172 40572
rect 39228 38668 39284 44156
rect 39340 44146 39396 44156
rect 39340 43764 39396 43774
rect 39452 43764 39508 44268
rect 39676 44258 39732 44268
rect 39340 43762 39508 43764
rect 39340 43710 39342 43762
rect 39394 43710 39508 43762
rect 39340 43708 39508 43710
rect 39340 43698 39396 43708
rect 39788 42756 39844 45164
rect 39900 45126 39956 45164
rect 40012 45108 40068 46732
rect 40124 46564 40180 46574
rect 40236 46564 40292 47180
rect 40124 46562 40292 46564
rect 40124 46510 40126 46562
rect 40178 46510 40292 46562
rect 40124 46508 40292 46510
rect 40124 45220 40180 46508
rect 40348 45332 40404 47292
rect 40460 47254 40516 47292
rect 40572 47236 40628 47246
rect 40572 47142 40628 47180
rect 40572 46004 40628 46014
rect 40460 45778 40516 45790
rect 40460 45726 40462 45778
rect 40514 45726 40516 45778
rect 40460 45556 40516 45726
rect 40572 45778 40628 45948
rect 40572 45726 40574 45778
rect 40626 45726 40628 45778
rect 40572 45714 40628 45726
rect 40460 45490 40516 45500
rect 40348 45266 40404 45276
rect 40124 45154 40180 45164
rect 40236 45218 40292 45230
rect 40236 45166 40238 45218
rect 40290 45166 40292 45218
rect 40236 45108 40292 45166
rect 40684 45108 40740 47516
rect 40908 47348 40964 48190
rect 40908 47282 40964 47292
rect 41020 48132 41076 48142
rect 40796 47236 40852 47246
rect 40796 47142 40852 47180
rect 41020 47124 41076 48076
rect 41020 47058 41076 47068
rect 41020 46004 41076 46014
rect 40796 45892 40852 45902
rect 40796 45798 40852 45836
rect 41020 45332 41076 45948
rect 41244 45666 41300 45678
rect 41244 45614 41246 45666
rect 41298 45614 41300 45666
rect 41244 45556 41300 45614
rect 41244 45490 41300 45500
rect 41468 45332 41524 51436
rect 41692 51266 41748 51278
rect 41692 51214 41694 51266
rect 41746 51214 41748 51266
rect 41692 50428 41748 51214
rect 41580 50372 41748 50428
rect 41580 50036 41636 50372
rect 41580 49942 41636 49980
rect 41580 48916 41636 48926
rect 41580 48822 41636 48860
rect 41020 45330 41188 45332
rect 41020 45278 41022 45330
rect 41074 45278 41188 45330
rect 41020 45276 41188 45278
rect 41020 45266 41076 45276
rect 40236 45052 40740 45108
rect 40012 44210 40068 45052
rect 40012 44158 40014 44210
rect 40066 44158 40068 44210
rect 39900 43988 39956 43998
rect 39900 43762 39956 43932
rect 39900 43710 39902 43762
rect 39954 43710 39956 43762
rect 39900 43698 39956 43710
rect 40012 43540 40068 44158
rect 40348 44098 40404 44110
rect 40348 44046 40350 44098
rect 40402 44046 40404 44098
rect 40348 43764 40404 44046
rect 40348 43698 40404 43708
rect 40124 43540 40180 43550
rect 40012 43538 40180 43540
rect 40012 43486 40126 43538
rect 40178 43486 40180 43538
rect 40012 43484 40180 43486
rect 40124 43474 40180 43484
rect 39564 42700 39844 42756
rect 39900 43428 39956 43438
rect 39340 42196 39396 42206
rect 39340 41186 39396 42140
rect 39340 41134 39342 41186
rect 39394 41134 39396 41186
rect 39340 40628 39396 41134
rect 39340 40562 39396 40572
rect 39452 41972 39508 41982
rect 39340 40404 39396 40414
rect 39452 40404 39508 41916
rect 39340 40402 39508 40404
rect 39340 40350 39342 40402
rect 39394 40350 39508 40402
rect 39340 40348 39508 40350
rect 39340 39842 39396 40348
rect 39340 39790 39342 39842
rect 39394 39790 39396 39842
rect 39340 39778 39396 39790
rect 39564 39620 39620 42700
rect 39676 42532 39732 42542
rect 39676 40292 39732 42476
rect 39900 41972 39956 43372
rect 40012 41972 40068 41982
rect 39900 41970 40068 41972
rect 39900 41918 40014 41970
rect 40066 41918 40068 41970
rect 39900 41916 40068 41918
rect 40012 41300 40068 41916
rect 39788 41188 39844 41198
rect 39788 41094 39844 41132
rect 40012 41186 40068 41244
rect 40012 41134 40014 41186
rect 40066 41134 40068 41186
rect 40012 41122 40068 41134
rect 40460 41860 40516 45052
rect 40684 44772 40740 44782
rect 40684 44212 40740 44716
rect 40684 44118 40740 44156
rect 41020 44212 41076 44222
rect 41020 44118 41076 44156
rect 41132 44210 41188 45276
rect 41132 44158 41134 44210
rect 41186 44158 41188 44210
rect 41132 44146 41188 44158
rect 41244 45330 41524 45332
rect 41244 45278 41470 45330
rect 41522 45278 41524 45330
rect 41244 45276 41524 45278
rect 40796 43988 40852 43998
rect 40852 43932 40964 43988
rect 40796 43922 40852 43932
rect 40684 43876 40740 43886
rect 40684 42530 40740 43820
rect 40684 42478 40686 42530
rect 40738 42478 40740 42530
rect 40684 42084 40740 42478
rect 40908 42196 40964 43932
rect 41020 43764 41076 43774
rect 41020 43670 41076 43708
rect 41244 43316 41300 45276
rect 41468 45266 41524 45276
rect 41580 48580 41636 48590
rect 41356 45108 41412 45118
rect 41356 45014 41412 45052
rect 41468 44882 41524 44894
rect 41468 44830 41470 44882
rect 41522 44830 41524 44882
rect 41468 44548 41524 44830
rect 41468 44482 41524 44492
rect 41580 44436 41636 48524
rect 41916 47908 41972 52220
rect 42028 51380 42084 52892
rect 42140 52882 42196 52892
rect 42028 51314 42084 51324
rect 42140 52050 42196 52062
rect 42140 51998 42142 52050
rect 42194 51998 42196 52050
rect 42028 51044 42084 51054
rect 42028 49140 42084 50988
rect 42140 50428 42196 51998
rect 42252 51938 42308 53228
rect 42364 53172 42420 53340
rect 42476 53172 42532 53182
rect 42364 53170 42532 53172
rect 42364 53118 42478 53170
rect 42530 53118 42532 53170
rect 42364 53116 42532 53118
rect 42476 53106 42532 53116
rect 42700 52836 42756 53678
rect 42924 53618 42980 54012
rect 43484 54068 43540 55132
rect 43596 54852 43652 56588
rect 44156 55300 44212 57484
rect 44268 57446 44324 57484
rect 44604 57428 44660 57438
rect 44604 56980 44660 57372
rect 44604 56914 44660 56924
rect 44828 56866 44884 57708
rect 45164 57698 45220 57708
rect 45276 58434 45332 58446
rect 45276 58382 45278 58434
rect 45330 58382 45332 58434
rect 45276 57428 45332 58382
rect 46172 58324 46228 59054
rect 46396 58324 46452 58334
rect 46172 58322 46452 58324
rect 46172 58270 46398 58322
rect 46450 58270 46452 58322
rect 46172 58268 46452 58270
rect 45612 57876 45668 57886
rect 45612 57782 45668 57820
rect 45836 57876 45892 57886
rect 46172 57876 46228 57886
rect 45836 57874 46228 57876
rect 45836 57822 45838 57874
rect 45890 57822 46174 57874
rect 46226 57822 46228 57874
rect 45836 57820 46228 57822
rect 45836 57810 45892 57820
rect 46172 57810 46228 57820
rect 45500 57650 45556 57662
rect 45500 57598 45502 57650
rect 45554 57598 45556 57650
rect 45500 57540 45556 57598
rect 45500 57474 45556 57484
rect 46060 57650 46116 57662
rect 46060 57598 46062 57650
rect 46114 57598 46116 57650
rect 44828 56814 44830 56866
rect 44882 56814 44884 56866
rect 44828 56802 44884 56814
rect 44940 57372 45332 57428
rect 44940 56642 44996 57372
rect 45164 57204 45220 57214
rect 44940 56590 44942 56642
rect 44994 56590 44996 56642
rect 44604 55972 44660 55982
rect 44156 55244 44324 55300
rect 43932 55188 43988 55198
rect 43932 55094 43988 55132
rect 44044 55076 44100 55086
rect 44044 54982 44100 55020
rect 44156 55074 44212 55086
rect 44156 55022 44158 55074
rect 44210 55022 44212 55074
rect 43596 54796 43764 54852
rect 43596 54628 43652 54638
rect 43596 54534 43652 54572
rect 43708 54404 43764 54796
rect 44156 54740 44212 55022
rect 44044 54738 44212 54740
rect 44044 54686 44158 54738
rect 44210 54686 44212 54738
rect 44044 54684 44212 54686
rect 43484 54002 43540 54012
rect 43596 54348 43764 54404
rect 43820 54404 43876 54414
rect 42924 53566 42926 53618
rect 42978 53566 42980 53618
rect 42924 53554 42980 53566
rect 43372 53730 43428 53742
rect 43372 53678 43374 53730
rect 43426 53678 43428 53730
rect 42924 52836 42980 52846
rect 43372 52836 43428 53678
rect 42700 52834 43428 52836
rect 42700 52782 42926 52834
rect 42978 52782 43374 52834
rect 43426 52782 43428 52834
rect 42700 52780 43428 52782
rect 42924 52770 42980 52780
rect 42252 51886 42254 51938
rect 42306 51886 42308 51938
rect 42252 51874 42308 51886
rect 42476 51940 42532 51950
rect 42476 51938 42756 51940
rect 42476 51886 42478 51938
rect 42530 51886 42756 51938
rect 42476 51884 42756 51886
rect 42476 51874 42532 51884
rect 42700 51492 42756 51884
rect 42588 51380 42644 51390
rect 42588 51286 42644 51324
rect 42700 51266 42756 51436
rect 42700 51214 42702 51266
rect 42754 51214 42756 51266
rect 42700 51202 42756 51214
rect 42812 51938 42868 51950
rect 42812 51886 42814 51938
rect 42866 51886 42868 51938
rect 42812 51044 42868 51886
rect 42700 50988 42868 51044
rect 42924 51154 42980 51166
rect 42924 51102 42926 51154
rect 42978 51102 42980 51154
rect 42700 50428 42756 50988
rect 42140 50372 42756 50428
rect 42812 50594 42868 50606
rect 42812 50542 42814 50594
rect 42866 50542 42868 50594
rect 42028 49084 42196 49140
rect 41692 47852 41972 47908
rect 41692 45444 41748 47852
rect 41804 47684 41860 47694
rect 41804 47458 41860 47628
rect 41804 47406 41806 47458
rect 41858 47406 41860 47458
rect 41804 47394 41860 47406
rect 41916 47570 41972 47582
rect 41916 47518 41918 47570
rect 41970 47518 41972 47570
rect 41804 47124 41860 47134
rect 41804 45556 41860 47068
rect 41916 46564 41972 47518
rect 42028 46564 42084 46574
rect 41916 46562 42084 46564
rect 41916 46510 42030 46562
rect 42082 46510 42084 46562
rect 41916 46508 42084 46510
rect 42028 45892 42084 46508
rect 42140 46452 42196 49084
rect 42252 47236 42308 47246
rect 42252 46676 42308 47180
rect 42476 46676 42532 50372
rect 42812 49588 42868 50542
rect 42924 50484 42980 51102
rect 43036 50708 43092 50718
rect 43036 50614 43092 50652
rect 43148 50484 43204 50494
rect 42924 50482 43316 50484
rect 42924 50430 43150 50482
rect 43202 50430 43316 50482
rect 42924 50428 43316 50430
rect 43148 50418 43204 50428
rect 43260 49810 43316 50428
rect 43260 49758 43262 49810
rect 43314 49758 43316 49810
rect 43260 49746 43316 49758
rect 42812 49522 42868 49532
rect 43260 49252 43316 49262
rect 43260 48468 43316 49196
rect 43260 48402 43316 48412
rect 43036 48356 43092 48366
rect 42924 48354 43092 48356
rect 42924 48302 43038 48354
rect 43090 48302 43092 48354
rect 42924 48300 43092 48302
rect 42588 48242 42644 48254
rect 42588 48190 42590 48242
rect 42642 48190 42644 48242
rect 42588 46898 42644 48190
rect 42812 48242 42868 48254
rect 42812 48190 42814 48242
rect 42866 48190 42868 48242
rect 42588 46846 42590 46898
rect 42642 46846 42644 46898
rect 42588 46834 42644 46846
rect 42700 48130 42756 48142
rect 42700 48078 42702 48130
rect 42754 48078 42756 48130
rect 42700 46676 42756 48078
rect 42812 47684 42868 48190
rect 42812 47618 42868 47628
rect 42812 47458 42868 47470
rect 42812 47406 42814 47458
rect 42866 47406 42868 47458
rect 42812 47236 42868 47406
rect 42812 47170 42868 47180
rect 42252 46674 42420 46676
rect 42252 46622 42254 46674
rect 42306 46622 42420 46674
rect 42252 46620 42420 46622
rect 42476 46620 42644 46676
rect 42252 46610 42308 46620
rect 42364 46564 42420 46620
rect 42364 46508 42532 46564
rect 42140 46396 42420 46452
rect 42252 45892 42308 45902
rect 42028 45836 42252 45892
rect 42252 45798 42308 45836
rect 41804 45500 41972 45556
rect 41692 45388 41860 45444
rect 41580 44370 41636 44380
rect 41692 45220 41748 45230
rect 41356 44324 41412 44334
rect 41412 44268 41524 44324
rect 41356 44258 41412 44268
rect 41468 44212 41524 44268
rect 41580 44212 41636 44222
rect 41468 44210 41636 44212
rect 41468 44158 41582 44210
rect 41634 44158 41636 44210
rect 41468 44156 41636 44158
rect 41580 44146 41636 44156
rect 41692 44210 41748 45164
rect 41692 44158 41694 44210
rect 41746 44158 41748 44210
rect 41692 44146 41748 44158
rect 41356 44100 41412 44110
rect 41356 44098 41524 44100
rect 41356 44046 41358 44098
rect 41410 44046 41524 44098
rect 41356 44044 41524 44046
rect 41356 44034 41412 44044
rect 41468 43540 41524 44044
rect 41692 43988 41748 43998
rect 41580 43540 41636 43550
rect 41468 43484 41580 43540
rect 41580 43446 41636 43484
rect 41244 43260 41524 43316
rect 41244 42868 41300 42878
rect 41244 42774 41300 42812
rect 40908 42140 41076 42196
rect 40684 42018 40740 42028
rect 40908 41970 40964 41982
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40908 41860 40964 41918
rect 40460 41804 40964 41860
rect 40460 41186 40516 41804
rect 40460 41134 40462 41186
rect 40514 41134 40516 41186
rect 40460 41122 40516 41134
rect 40572 41300 40628 41310
rect 41020 41300 41076 42140
rect 40572 41186 40628 41244
rect 40572 41134 40574 41186
rect 40626 41134 40628 41186
rect 40572 41122 40628 41134
rect 40908 41244 41076 41300
rect 41244 42082 41300 42094
rect 41244 42030 41246 42082
rect 41298 42030 41300 42082
rect 40684 41074 40740 41086
rect 40684 41022 40686 41074
rect 40738 41022 40740 41074
rect 39900 40962 39956 40974
rect 39900 40910 39902 40962
rect 39954 40910 39956 40962
rect 39788 40628 39844 40638
rect 39900 40628 39956 40910
rect 40684 40628 40740 41022
rect 39900 40572 40180 40628
rect 39788 40404 39844 40572
rect 39900 40404 39956 40414
rect 39788 40402 39956 40404
rect 39788 40350 39902 40402
rect 39954 40350 39956 40402
rect 39788 40348 39956 40350
rect 39900 40338 39956 40348
rect 39676 40236 39844 40292
rect 39564 39554 39620 39564
rect 39340 39508 39396 39518
rect 39340 38948 39396 39452
rect 39676 39508 39732 39518
rect 39676 39414 39732 39452
rect 39340 38882 39396 38892
rect 39788 38668 39844 40236
rect 39228 38612 39396 38668
rect 39788 38612 40068 38668
rect 38556 38332 39060 38388
rect 38444 38164 38500 38174
rect 38332 38162 38500 38164
rect 38332 38110 38446 38162
rect 38498 38110 38500 38162
rect 38332 38108 38500 38110
rect 38108 37380 38164 37390
rect 38108 37286 38164 37324
rect 38332 36484 38388 38108
rect 38444 38098 38500 38108
rect 38556 37828 38612 38332
rect 38780 38052 38836 38062
rect 38780 37958 38836 37996
rect 38444 37826 38612 37828
rect 38444 37774 38558 37826
rect 38610 37774 38612 37826
rect 38444 37772 38612 37774
rect 39004 37828 39060 38332
rect 39228 37828 39284 37838
rect 39004 37826 39284 37828
rect 39004 37774 39230 37826
rect 39282 37774 39284 37826
rect 39004 37772 39284 37774
rect 38444 37266 38500 37772
rect 38556 37762 38612 37772
rect 38444 37214 38446 37266
rect 38498 37214 38500 37266
rect 38444 37202 38500 37214
rect 38332 36418 38388 36428
rect 39116 36372 39172 36382
rect 39116 36278 39172 36316
rect 38444 36258 38500 36270
rect 38780 36260 38836 36270
rect 38444 36206 38446 36258
rect 38498 36206 38500 36258
rect 37996 35868 38276 35924
rect 38108 35700 38164 35710
rect 37772 34130 37940 34132
rect 37772 34078 37774 34130
rect 37826 34078 37940 34130
rect 37772 34076 37940 34078
rect 37996 35698 38164 35700
rect 37996 35646 38110 35698
rect 38162 35646 38164 35698
rect 37996 35644 38164 35646
rect 37772 34066 37828 34076
rect 37548 33964 37716 34020
rect 37436 33294 37438 33346
rect 37490 33294 37492 33346
rect 37436 33282 37492 33294
rect 37548 33684 37604 33694
rect 37212 33058 37268 33068
rect 37212 32676 37268 32686
rect 37212 32582 37268 32620
rect 37436 32564 37492 32574
rect 37436 32470 37492 32508
rect 36876 32340 36932 32350
rect 36876 26908 36932 32284
rect 37436 31668 37492 31678
rect 36988 30212 37044 30222
rect 36988 30118 37044 30156
rect 37100 30210 37156 30222
rect 37100 30158 37102 30210
rect 37154 30158 37156 30210
rect 37100 29988 37156 30158
rect 37436 30210 37492 31612
rect 37548 30994 37604 33628
rect 37548 30942 37550 30994
rect 37602 30942 37604 30994
rect 37548 30930 37604 30942
rect 37436 30158 37438 30210
rect 37490 30158 37492 30210
rect 37436 30146 37492 30158
rect 37660 29988 37716 33964
rect 37884 33460 37940 33470
rect 37884 30996 37940 33404
rect 37996 33458 38052 35644
rect 38108 35634 38164 35644
rect 38108 35476 38164 35486
rect 38108 34242 38164 35420
rect 38108 34190 38110 34242
rect 38162 34190 38164 34242
rect 38108 34178 38164 34190
rect 37996 33406 37998 33458
rect 38050 33406 38052 33458
rect 37996 33394 38052 33406
rect 38220 32674 38276 35868
rect 38444 35700 38500 36206
rect 38444 35634 38500 35644
rect 38556 36258 38836 36260
rect 38556 36206 38782 36258
rect 38834 36206 38836 36258
rect 38556 36204 38836 36206
rect 38556 35586 38612 36204
rect 38780 36194 38836 36204
rect 39228 36260 39284 37772
rect 39228 36194 39284 36204
rect 39004 35700 39060 35738
rect 39340 35700 39396 38612
rect 39564 38052 39620 38062
rect 39452 37996 39564 38052
rect 39452 36708 39508 37996
rect 39564 37986 39620 37996
rect 39900 38052 39956 38062
rect 39900 37958 39956 37996
rect 39676 37826 39732 37838
rect 39676 37774 39678 37826
rect 39730 37774 39732 37826
rect 39564 37380 39620 37390
rect 39676 37380 39732 37774
rect 39564 37378 39732 37380
rect 39564 37326 39566 37378
rect 39618 37326 39732 37378
rect 39564 37324 39732 37326
rect 39788 37380 39844 37390
rect 39564 37314 39620 37324
rect 39452 36652 39732 36708
rect 39452 36484 39508 36494
rect 39452 36390 39508 36428
rect 39004 35634 39060 35644
rect 39228 35644 39396 35700
rect 39676 35810 39732 36652
rect 39788 36482 39844 37324
rect 40012 36596 40068 38612
rect 40124 36820 40180 40572
rect 40684 40562 40740 40572
rect 40236 40516 40292 40526
rect 40236 39844 40292 40460
rect 40796 40516 40852 40526
rect 40796 40404 40852 40460
rect 40684 40348 40852 40404
rect 40236 39788 40404 39844
rect 40236 39620 40292 39630
rect 40236 39526 40292 39564
rect 40348 39396 40404 39788
rect 40236 39340 40404 39396
rect 40236 37380 40292 39340
rect 40460 38836 40516 38846
rect 40236 37324 40404 37380
rect 40124 36754 40180 36764
rect 40236 37154 40292 37166
rect 40236 37102 40238 37154
rect 40290 37102 40292 37154
rect 40236 36932 40292 37102
rect 40012 36540 40180 36596
rect 39788 36430 39790 36482
rect 39842 36430 39844 36482
rect 39788 36418 39844 36430
rect 39900 36372 39956 36382
rect 39900 36278 39956 36316
rect 40012 36370 40068 36382
rect 40012 36318 40014 36370
rect 40066 36318 40068 36370
rect 39676 35758 39678 35810
rect 39730 35758 39732 35810
rect 38556 35534 38558 35586
rect 38610 35534 38612 35586
rect 38556 35522 38612 35534
rect 39004 35476 39060 35486
rect 39004 35382 39060 35420
rect 38556 35252 38612 35262
rect 38332 34916 38388 34926
rect 38332 33684 38388 34860
rect 38444 34916 38500 34926
rect 38556 34916 38612 35196
rect 39228 34916 39284 35644
rect 39340 35474 39396 35486
rect 39340 35422 39342 35474
rect 39394 35422 39396 35474
rect 39340 35252 39396 35422
rect 39340 35186 39396 35196
rect 39676 35138 39732 35758
rect 39788 36260 39844 36270
rect 39788 35810 39844 36204
rect 39788 35758 39790 35810
rect 39842 35758 39844 35810
rect 39788 35700 39844 35758
rect 39788 35634 39844 35644
rect 39900 36148 39956 36158
rect 39676 35086 39678 35138
rect 39730 35086 39732 35138
rect 39676 35074 39732 35086
rect 38444 34914 38612 34916
rect 38444 34862 38446 34914
rect 38498 34862 38612 34914
rect 38444 34860 38612 34862
rect 38444 34850 38500 34860
rect 38388 33628 38500 33684
rect 38332 33618 38388 33628
rect 38444 33346 38500 33628
rect 38444 33294 38446 33346
rect 38498 33294 38500 33346
rect 38444 33282 38500 33294
rect 38556 33348 38612 34860
rect 38892 34914 39284 34916
rect 38892 34862 39230 34914
rect 39282 34862 39284 34914
rect 38892 34860 39284 34862
rect 38780 33348 38836 33358
rect 38556 33346 38836 33348
rect 38556 33294 38782 33346
rect 38834 33294 38836 33346
rect 38556 33292 38836 33294
rect 38220 32622 38222 32674
rect 38274 32622 38276 32674
rect 38220 32610 38276 32622
rect 38332 33234 38388 33246
rect 38332 33182 38334 33234
rect 38386 33182 38388 33234
rect 38332 32676 38388 33182
rect 38556 32786 38612 32798
rect 38556 32734 38558 32786
rect 38610 32734 38612 32786
rect 38444 32676 38500 32686
rect 38332 32674 38500 32676
rect 38332 32622 38446 32674
rect 38498 32622 38500 32674
rect 38332 32620 38500 32622
rect 38444 32610 38500 32620
rect 38556 32564 38612 32734
rect 38556 32498 38612 32508
rect 38780 31668 38836 33292
rect 38892 32562 38948 34860
rect 39228 34850 39284 34860
rect 39676 34804 39732 34814
rect 39900 34804 39956 36092
rect 40012 35922 40068 36318
rect 40012 35870 40014 35922
rect 40066 35870 40068 35922
rect 40012 35858 40068 35870
rect 39732 34748 39956 34804
rect 38892 32510 38894 32562
rect 38946 32510 38948 32562
rect 38892 32498 38948 32510
rect 39004 34020 39060 34030
rect 39004 32340 39060 33964
rect 39676 34020 39732 34748
rect 39676 33926 39732 33964
rect 40124 33348 40180 36540
rect 40236 35924 40292 36876
rect 40348 36148 40404 37324
rect 40348 36082 40404 36092
rect 40348 35924 40404 35934
rect 40236 35922 40404 35924
rect 40236 35870 40350 35922
rect 40402 35870 40404 35922
rect 40236 35868 40404 35870
rect 40348 35858 40404 35868
rect 40236 35700 40292 35710
rect 40236 34354 40292 35644
rect 40236 34302 40238 34354
rect 40290 34302 40292 34354
rect 40236 34290 40292 34302
rect 40348 34690 40404 34702
rect 40348 34638 40350 34690
rect 40402 34638 40404 34690
rect 40348 34244 40404 34638
rect 40348 34178 40404 34188
rect 40460 33908 40516 38780
rect 40572 36258 40628 36270
rect 40572 36206 40574 36258
rect 40626 36206 40628 36258
rect 40572 35700 40628 36206
rect 40572 35634 40628 35644
rect 40684 35140 40740 40348
rect 40908 39620 40964 41244
rect 41244 41188 41300 42030
rect 41020 41132 41244 41188
rect 41020 40628 41076 41132
rect 41244 41122 41300 41132
rect 41132 40964 41188 40974
rect 41132 40962 41412 40964
rect 41132 40910 41134 40962
rect 41186 40910 41412 40962
rect 41132 40908 41412 40910
rect 41132 40898 41188 40908
rect 41244 40740 41300 40750
rect 41132 40628 41188 40638
rect 41020 40626 41188 40628
rect 41020 40574 41134 40626
rect 41186 40574 41188 40626
rect 41020 40572 41188 40574
rect 41132 40562 41188 40572
rect 41132 39620 41188 39630
rect 40908 39618 41132 39620
rect 40908 39566 40910 39618
rect 40962 39566 41132 39618
rect 40908 39564 41132 39566
rect 40908 39554 40964 39564
rect 40796 39060 40852 39070
rect 40796 35252 40852 39004
rect 41020 38948 41076 38958
rect 40908 38892 41020 38948
rect 40908 37266 40964 38892
rect 41020 38882 41076 38892
rect 41020 38724 41076 38734
rect 41132 38724 41188 39564
rect 41244 39508 41300 40684
rect 41244 39414 41300 39452
rect 41020 38722 41188 38724
rect 41020 38670 41022 38722
rect 41074 38670 41188 38722
rect 41020 38668 41188 38670
rect 41020 38658 41076 38668
rect 41132 37268 41188 37278
rect 40908 37214 40910 37266
rect 40962 37214 40964 37266
rect 40908 37202 40964 37214
rect 41020 37212 41132 37268
rect 40908 36372 40964 36382
rect 41020 36372 41076 37212
rect 41132 37174 41188 37212
rect 40908 36370 41076 36372
rect 40908 36318 40910 36370
rect 40962 36318 41076 36370
rect 40908 36316 41076 36318
rect 41132 36820 41188 36830
rect 40908 36306 40964 36316
rect 41132 35812 41188 36764
rect 41244 36484 41300 36494
rect 41244 36390 41300 36428
rect 41132 35718 41188 35756
rect 41356 35698 41412 40908
rect 41468 39058 41524 43260
rect 41580 41300 41636 41310
rect 41580 41206 41636 41244
rect 41580 41076 41636 41086
rect 41580 40514 41636 41020
rect 41692 40628 41748 43932
rect 41692 40534 41748 40572
rect 41580 40462 41582 40514
rect 41634 40462 41636 40514
rect 41580 40180 41636 40462
rect 41804 40292 41860 45388
rect 41916 44324 41972 45500
rect 42028 45220 42084 45230
rect 42028 45126 42084 45164
rect 41916 44268 42196 44324
rect 41916 44098 41972 44110
rect 41916 44046 41918 44098
rect 41970 44046 41972 44098
rect 41916 43708 41972 44046
rect 42028 43764 42084 43784
rect 41916 43652 42084 43708
rect 42028 43538 42084 43652
rect 42028 43486 42030 43538
rect 42082 43486 42084 43538
rect 42028 43474 42084 43486
rect 41916 42868 41972 42878
rect 41916 42532 41972 42812
rect 42140 42644 42196 44268
rect 41916 40740 41972 42476
rect 42028 42588 42196 42644
rect 42028 41076 42084 42588
rect 42252 42532 42308 42542
rect 42028 41010 42084 41020
rect 42140 42530 42308 42532
rect 42140 42478 42254 42530
rect 42306 42478 42308 42530
rect 42140 42476 42308 42478
rect 41916 40674 41972 40684
rect 41916 40404 41972 40414
rect 41916 40402 42084 40404
rect 41916 40350 41918 40402
rect 41970 40350 42084 40402
rect 41916 40348 42084 40350
rect 41916 40338 41972 40348
rect 41580 40114 41636 40124
rect 41692 40236 41860 40292
rect 41580 39620 41636 39630
rect 41580 39526 41636 39564
rect 41468 39006 41470 39058
rect 41522 39006 41524 39058
rect 41468 38668 41524 39006
rect 41692 39506 41748 40236
rect 42028 40178 42084 40348
rect 42028 40126 42030 40178
rect 42082 40126 42084 40178
rect 42028 40114 42084 40126
rect 42140 39956 42196 42476
rect 42252 42466 42308 42476
rect 42252 40628 42308 40638
rect 42252 40534 42308 40572
rect 41692 39454 41694 39506
rect 41746 39454 41748 39506
rect 41692 38948 41748 39454
rect 41804 39900 42196 39956
rect 41804 39060 41860 39900
rect 41916 39620 41972 39630
rect 41916 39526 41972 39564
rect 41804 38966 41860 39004
rect 42252 39508 42308 39518
rect 42252 39058 42308 39452
rect 42252 39006 42254 39058
rect 42306 39006 42308 39058
rect 41692 38882 41748 38892
rect 41468 38612 41972 38668
rect 41916 37490 41972 38612
rect 41916 37438 41918 37490
rect 41970 37438 41972 37490
rect 41916 37426 41972 37438
rect 41804 37268 41860 37278
rect 41804 37174 41860 37212
rect 42140 37268 42196 37278
rect 42140 37174 42196 37212
rect 41468 37044 41524 37054
rect 41468 37042 41860 37044
rect 41468 36990 41470 37042
rect 41522 36990 41860 37042
rect 41468 36988 41860 36990
rect 41468 36978 41524 36988
rect 41692 36484 41748 36494
rect 41692 36390 41748 36428
rect 41356 35646 41358 35698
rect 41410 35646 41412 35698
rect 40796 35196 41076 35252
rect 40460 33842 40516 33852
rect 40572 35084 40740 35140
rect 40572 33460 40628 35084
rect 40908 34804 40964 34814
rect 40908 34710 40964 34748
rect 41020 34802 41076 35196
rect 41244 34916 41300 34926
rect 41356 34916 41412 35646
rect 41692 35476 41748 35486
rect 41692 35382 41748 35420
rect 41692 35140 41748 35150
rect 41468 34916 41524 34926
rect 41356 34914 41524 34916
rect 41356 34862 41470 34914
rect 41522 34862 41524 34914
rect 41356 34860 41524 34862
rect 41244 34822 41300 34860
rect 41468 34850 41524 34860
rect 41020 34750 41022 34802
rect 41074 34750 41076 34802
rect 41020 34130 41076 34750
rect 41020 34078 41022 34130
rect 41074 34078 41076 34130
rect 39900 33292 40180 33348
rect 40236 33404 40628 33460
rect 40908 33908 40964 33918
rect 39788 33236 39844 33246
rect 39788 33142 39844 33180
rect 39564 33124 39620 33134
rect 39564 32786 39620 33068
rect 39564 32734 39566 32786
rect 39618 32734 39620 32786
rect 39564 32722 39620 32734
rect 39788 32900 39844 32910
rect 39788 32674 39844 32844
rect 39788 32622 39790 32674
rect 39842 32622 39844 32674
rect 39788 32610 39844 32622
rect 38780 31602 38836 31612
rect 38892 32284 39060 32340
rect 38556 31556 38612 31566
rect 37884 30994 38388 30996
rect 37884 30942 37886 30994
rect 37938 30942 38388 30994
rect 37884 30940 38388 30942
rect 37884 30930 37940 30940
rect 37156 29932 37380 29988
rect 37100 29922 37156 29932
rect 37324 29426 37380 29932
rect 37324 29374 37326 29426
rect 37378 29374 37380 29426
rect 37324 29362 37380 29374
rect 37436 29932 37716 29988
rect 37324 28530 37380 28542
rect 37324 28478 37326 28530
rect 37378 28478 37380 28530
rect 36988 27748 37044 27758
rect 37324 27748 37380 28478
rect 36988 27746 37380 27748
rect 36988 27694 36990 27746
rect 37042 27694 37380 27746
rect 36988 27692 37380 27694
rect 37436 27748 37492 29932
rect 38332 29538 38388 30940
rect 38556 30994 38612 31500
rect 38556 30942 38558 30994
rect 38610 30942 38612 30994
rect 38556 30930 38612 30942
rect 38444 29986 38500 29998
rect 38444 29934 38446 29986
rect 38498 29934 38500 29986
rect 38444 29876 38500 29934
rect 38500 29820 38612 29876
rect 38444 29810 38500 29820
rect 38332 29486 38334 29538
rect 38386 29486 38388 29538
rect 38332 29474 38388 29486
rect 38108 28756 38164 28766
rect 37660 28532 37716 28542
rect 37660 28438 37716 28476
rect 37548 28084 37604 28094
rect 37548 27970 37604 28028
rect 37548 27918 37550 27970
rect 37602 27918 37604 27970
rect 37548 27906 37604 27918
rect 37436 27692 37604 27748
rect 36988 27188 37044 27692
rect 36988 27122 37044 27132
rect 37436 27074 37492 27086
rect 37436 27022 37438 27074
rect 37490 27022 37492 27074
rect 36876 26852 37268 26908
rect 37212 25618 37268 26852
rect 37212 25566 37214 25618
rect 37266 25566 37268 25618
rect 36876 24948 36932 24958
rect 37212 24948 37268 25566
rect 36876 24946 37212 24948
rect 36876 24894 36878 24946
rect 36930 24894 37212 24946
rect 36876 24892 37212 24894
rect 36876 24882 36932 24892
rect 37212 24722 37268 24892
rect 37212 24670 37214 24722
rect 37266 24670 37268 24722
rect 37212 24658 37268 24670
rect 37436 24834 37492 27022
rect 37436 24782 37438 24834
rect 37490 24782 37492 24834
rect 37324 23940 37380 23950
rect 37100 23938 37380 23940
rect 37100 23886 37326 23938
rect 37378 23886 37380 23938
rect 37100 23884 37380 23886
rect 37100 23156 37156 23884
rect 37324 23874 37380 23884
rect 37436 23492 37492 24782
rect 37436 23426 37492 23436
rect 37548 23268 37604 27692
rect 37660 27300 37716 27310
rect 37660 27206 37716 27244
rect 37996 27300 38052 27310
rect 37996 27206 38052 27244
rect 37996 25060 38052 25070
rect 37884 24948 37940 24958
rect 37884 24854 37940 24892
rect 37996 24834 38052 25004
rect 37996 24782 37998 24834
rect 38050 24782 38052 24834
rect 37996 24724 38052 24782
rect 37772 24668 38052 24724
rect 37660 24612 37716 24622
rect 37660 23938 37716 24556
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 37660 23874 37716 23886
rect 37660 23716 37716 23726
rect 37660 23622 37716 23660
rect 36988 23154 37156 23156
rect 36988 23102 37102 23154
rect 37154 23102 37156 23154
rect 36988 23100 37156 23102
rect 36988 22482 37044 23100
rect 37100 23090 37156 23100
rect 37212 23212 37604 23268
rect 36988 22430 36990 22482
rect 37042 22430 37044 22482
rect 36988 22418 37044 22430
rect 36876 20018 36932 20030
rect 36876 19966 36878 20018
rect 36930 19966 36932 20018
rect 36876 19572 36932 19966
rect 37100 20020 37156 20030
rect 37212 20020 37268 23212
rect 37772 22596 37828 24668
rect 37548 22540 37828 22596
rect 37884 24498 37940 24510
rect 37884 24446 37886 24498
rect 37938 24446 37940 24498
rect 37436 22482 37492 22494
rect 37436 22430 37438 22482
rect 37490 22430 37492 22482
rect 37436 22260 37492 22430
rect 37436 22194 37492 22204
rect 37436 21924 37492 21934
rect 37100 20018 37268 20020
rect 37100 19966 37102 20018
rect 37154 19966 37268 20018
rect 37100 19964 37268 19966
rect 37324 20132 37380 20142
rect 37100 19796 37156 19964
rect 37100 19730 37156 19740
rect 36876 19506 36932 19516
rect 37212 19348 37268 19358
rect 37212 19254 37268 19292
rect 36988 19236 37044 19246
rect 36988 19142 37044 19180
rect 37100 18564 37156 18574
rect 37100 17780 37156 18508
rect 37212 18338 37268 18350
rect 37212 18286 37214 18338
rect 37266 18286 37268 18338
rect 37212 18228 37268 18286
rect 37212 18162 37268 18172
rect 37212 17780 37268 17790
rect 37100 17778 37268 17780
rect 37100 17726 37214 17778
rect 37266 17726 37268 17778
rect 37100 17724 37268 17726
rect 37212 17714 37268 17724
rect 37100 16212 37156 16222
rect 36204 16210 36596 16212
rect 36204 16158 36206 16210
rect 36258 16158 36596 16210
rect 36204 16156 36596 16158
rect 36204 16146 36260 16156
rect 35980 15374 35982 15426
rect 36034 15374 36036 15426
rect 35868 15316 35924 15326
rect 35980 15316 36036 15374
rect 36540 15426 36596 16156
rect 36540 15374 36542 15426
rect 36594 15374 36596 15426
rect 36540 15362 36596 15374
rect 36764 16210 37156 16212
rect 36764 16158 37102 16210
rect 37154 16158 37156 16210
rect 36764 16156 37156 16158
rect 35084 15092 35364 15148
rect 35420 15260 35700 15316
rect 35420 15202 35476 15260
rect 35420 15150 35422 15202
rect 35474 15150 35476 15202
rect 35420 15138 35476 15150
rect 35084 14756 35140 15092
rect 35532 15090 35588 15102
rect 35532 15038 35534 15090
rect 35586 15038 35588 15090
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14700 35252 14756
rect 34972 14588 35140 14644
rect 34412 14420 34468 14430
rect 34412 14418 34804 14420
rect 34412 14366 34414 14418
rect 34466 14366 34804 14418
rect 34412 14364 34804 14366
rect 34412 14354 34468 14364
rect 34300 14308 34356 14318
rect 33740 14306 34356 14308
rect 33740 14254 34302 14306
rect 34354 14254 34356 14306
rect 33740 14252 34356 14254
rect 34300 14242 34356 14252
rect 34748 13858 34804 14364
rect 34748 13806 34750 13858
rect 34802 13806 34804 13858
rect 34748 12962 34804 13806
rect 34748 12910 34750 12962
rect 34802 12910 34804 12962
rect 34748 12898 34804 12910
rect 34972 14418 35028 14430
rect 34972 14366 34974 14418
rect 35026 14366 35028 14418
rect 34972 12962 35028 14366
rect 34972 12910 34974 12962
rect 35026 12910 35028 12962
rect 34972 12898 35028 12910
rect 34972 12738 35028 12750
rect 34972 12686 34974 12738
rect 35026 12686 35028 12738
rect 34188 11508 34244 11518
rect 33740 11396 33796 11406
rect 33740 11302 33796 11340
rect 34188 11394 34244 11452
rect 34188 11342 34190 11394
rect 34242 11342 34244 11394
rect 34188 10834 34244 11342
rect 34188 10782 34190 10834
rect 34242 10782 34244 10834
rect 34188 10770 34244 10782
rect 34972 10724 35028 12686
rect 35084 11508 35140 14588
rect 35196 13746 35252 14700
rect 35420 14530 35476 14542
rect 35420 14478 35422 14530
rect 35474 14478 35476 14530
rect 35420 14420 35476 14478
rect 35420 14354 35476 14364
rect 35196 13694 35198 13746
rect 35250 13694 35252 13746
rect 35196 13682 35252 13694
rect 35532 14308 35588 15038
rect 35532 13634 35588 14252
rect 35532 13582 35534 13634
rect 35586 13582 35588 13634
rect 35532 13570 35588 13582
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35644 13076 35700 15260
rect 35924 15260 36036 15316
rect 36092 15316 36148 15326
rect 35868 15250 35924 15260
rect 36092 15222 36148 15260
rect 36764 15316 36820 16156
rect 37100 16146 37156 16156
rect 36764 15148 36820 15260
rect 36652 15092 36820 15148
rect 36876 15426 36932 15438
rect 36876 15374 36878 15426
rect 36930 15374 36932 15426
rect 35868 14644 35924 14654
rect 35868 14550 35924 14588
rect 36540 14644 36596 14654
rect 36652 14644 36708 15092
rect 36540 14642 36708 14644
rect 36540 14590 36542 14642
rect 36594 14590 36708 14642
rect 36540 14588 36708 14590
rect 36540 14578 36596 14588
rect 36876 14532 36932 15374
rect 37324 15316 37380 20076
rect 37436 18676 37492 21868
rect 37548 19908 37604 22540
rect 37660 22372 37716 22382
rect 37884 22372 37940 24446
rect 37996 23826 38052 23838
rect 37996 23774 37998 23826
rect 38050 23774 38052 23826
rect 37996 22932 38052 23774
rect 38108 23266 38164 28700
rect 38556 28642 38612 29820
rect 38556 28590 38558 28642
rect 38610 28590 38612 28642
rect 38556 28578 38612 28590
rect 38668 28754 38724 28766
rect 38668 28702 38670 28754
rect 38722 28702 38724 28754
rect 38668 28532 38724 28702
rect 38556 27860 38612 27870
rect 38444 27804 38556 27860
rect 38332 27412 38388 27422
rect 38332 26514 38388 27356
rect 38444 26908 38500 27804
rect 38556 27766 38612 27804
rect 38668 27076 38724 28476
rect 38668 27010 38724 27020
rect 38780 28420 38836 28430
rect 38780 27300 38836 28364
rect 38780 26962 38836 27244
rect 38780 26910 38782 26962
rect 38834 26910 38836 26962
rect 38444 26852 38612 26908
rect 38780 26898 38836 26910
rect 38332 26462 38334 26514
rect 38386 26462 38388 26514
rect 38332 26450 38388 26462
rect 38444 25060 38500 25070
rect 38444 24946 38500 25004
rect 38444 24894 38446 24946
rect 38498 24894 38500 24946
rect 38444 24882 38500 24894
rect 38108 23214 38110 23266
rect 38162 23214 38164 23266
rect 38108 23202 38164 23214
rect 38332 23938 38388 23950
rect 38332 23886 38334 23938
rect 38386 23886 38388 23938
rect 38332 23268 38388 23886
rect 38332 23202 38388 23212
rect 37996 22876 38500 22932
rect 38444 22482 38500 22876
rect 38556 22596 38612 26852
rect 38780 25172 38836 25182
rect 38668 25116 38780 25172
rect 38668 22820 38724 25116
rect 38780 25106 38836 25116
rect 38892 23938 38948 32284
rect 39788 31668 39844 31678
rect 39116 29876 39172 29886
rect 39116 29538 39172 29820
rect 39564 29876 39620 29886
rect 39564 29650 39620 29820
rect 39564 29598 39566 29650
rect 39618 29598 39620 29650
rect 39564 29586 39620 29598
rect 39116 29486 39118 29538
rect 39170 29486 39172 29538
rect 39116 29474 39172 29486
rect 39564 29316 39620 29326
rect 39004 29204 39060 29214
rect 39004 29110 39060 29148
rect 39452 28868 39508 28878
rect 39452 28774 39508 28812
rect 39116 28644 39172 28654
rect 39004 28532 39060 28542
rect 39004 28438 39060 28476
rect 39004 28084 39060 28094
rect 39004 27074 39060 28028
rect 39004 27022 39006 27074
rect 39058 27022 39060 27074
rect 39004 27010 39060 27022
rect 38892 23886 38894 23938
rect 38946 23886 38948 23938
rect 38780 23380 38836 23390
rect 38892 23380 38948 23886
rect 38780 23378 38948 23380
rect 38780 23326 38782 23378
rect 38834 23326 38948 23378
rect 38780 23324 38948 23326
rect 39004 26516 39060 26526
rect 39004 24164 39060 26460
rect 39116 24948 39172 28588
rect 39340 28532 39396 28542
rect 39340 28084 39396 28476
rect 39452 28420 39508 28430
rect 39452 28326 39508 28364
rect 39564 28196 39620 29260
rect 39340 28018 39396 28028
rect 39452 28140 39620 28196
rect 39452 25060 39508 28140
rect 39564 27972 39620 27982
rect 39564 25172 39620 27916
rect 39788 27970 39844 31612
rect 39900 29316 39956 33292
rect 40124 33124 40180 33134
rect 40236 33124 40292 33404
rect 40180 33068 40292 33124
rect 40124 33030 40180 33068
rect 40012 32900 40068 32910
rect 40068 32844 40180 32900
rect 40012 32834 40068 32844
rect 40012 29986 40068 29998
rect 40012 29934 40014 29986
rect 40066 29934 40068 29986
rect 40012 29764 40068 29934
rect 40012 29698 40068 29708
rect 39900 29250 39956 29260
rect 39788 27918 39790 27970
rect 39842 27918 39844 27970
rect 39788 27906 39844 27918
rect 40124 27972 40180 32844
rect 40460 32788 40516 32798
rect 40348 32676 40404 32686
rect 40348 30210 40404 32620
rect 40348 30158 40350 30210
rect 40402 30158 40404 30210
rect 40348 30100 40404 30158
rect 40348 29876 40404 30044
rect 40236 29820 40404 29876
rect 40236 28754 40292 29820
rect 40348 29652 40404 29662
rect 40348 29558 40404 29596
rect 40460 29540 40516 32732
rect 40908 32788 40964 33852
rect 41020 33234 41076 34078
rect 41692 34018 41748 35084
rect 41692 33966 41694 34018
rect 41746 33966 41748 34018
rect 41244 33684 41300 33694
rect 41244 33346 41300 33628
rect 41244 33294 41246 33346
rect 41298 33294 41300 33346
rect 41020 33182 41022 33234
rect 41074 33182 41076 33234
rect 41020 33170 41076 33182
rect 41132 33236 41188 33246
rect 40908 32674 40964 32732
rect 40908 32622 40910 32674
rect 40962 32622 40964 32674
rect 40908 32610 40964 32622
rect 41132 31892 41188 33180
rect 41244 32900 41300 33294
rect 41356 33234 41412 33246
rect 41356 33182 41358 33234
rect 41410 33182 41412 33234
rect 41356 33124 41412 33182
rect 41356 33058 41412 33068
rect 41692 33012 41748 33966
rect 41692 32946 41748 32956
rect 41244 32844 41412 32900
rect 41356 32788 41412 32844
rect 41692 32788 41748 32798
rect 41356 32732 41524 32788
rect 41244 32676 41300 32686
rect 41244 32582 41300 32620
rect 41020 31890 41188 31892
rect 41020 31838 41134 31890
rect 41186 31838 41188 31890
rect 41020 31836 41188 31838
rect 40684 31556 40740 31566
rect 40684 31462 40740 31500
rect 40908 30882 40964 30894
rect 40908 30830 40910 30882
rect 40962 30830 40964 30882
rect 40572 30098 40628 30110
rect 40572 30046 40574 30098
rect 40626 30046 40628 30098
rect 40572 29764 40628 30046
rect 40572 29698 40628 29708
rect 40684 30100 40740 30110
rect 40908 30100 40964 30830
rect 40684 30098 40964 30100
rect 40684 30046 40686 30098
rect 40738 30046 40964 30098
rect 40684 30044 40964 30046
rect 40460 29484 40628 29540
rect 40236 28702 40238 28754
rect 40290 28702 40292 28754
rect 40236 28690 40292 28702
rect 40460 29316 40516 29326
rect 40460 28980 40516 29260
rect 40460 28866 40516 28924
rect 40460 28814 40462 28866
rect 40514 28814 40516 28866
rect 40236 28084 40292 28094
rect 40236 27990 40292 28028
rect 40124 27906 40180 27916
rect 40348 27860 40404 27870
rect 40348 27766 40404 27804
rect 40236 27636 40292 27646
rect 40236 27542 40292 27580
rect 39788 27412 39844 27422
rect 40460 27412 40516 28814
rect 39564 25106 39620 25116
rect 39676 27356 39788 27412
rect 39452 24994 39508 25004
rect 39564 24948 39620 24958
rect 39676 24948 39732 27356
rect 39788 27346 39844 27356
rect 40124 27356 40516 27412
rect 39900 27076 39956 27086
rect 39900 26982 39956 27020
rect 39116 24946 39396 24948
rect 39116 24894 39118 24946
rect 39170 24894 39396 24946
rect 39116 24892 39396 24894
rect 39116 24882 39172 24892
rect 39340 24836 39396 24892
rect 39564 24946 39732 24948
rect 39564 24894 39566 24946
rect 39618 24894 39732 24946
rect 39564 24892 39732 24894
rect 39564 24882 39620 24892
rect 39452 24836 39508 24846
rect 39340 24834 39508 24836
rect 39340 24782 39454 24834
rect 39506 24782 39508 24834
rect 39340 24780 39508 24782
rect 39004 24108 39284 24164
rect 38780 23314 38836 23324
rect 38668 22754 38724 22764
rect 38556 22540 38724 22596
rect 38444 22430 38446 22482
rect 38498 22430 38500 22482
rect 38444 22418 38500 22430
rect 37660 22370 37884 22372
rect 37660 22318 37662 22370
rect 37714 22318 37884 22370
rect 37660 22316 37884 22318
rect 37660 22306 37716 22316
rect 37884 22278 37940 22316
rect 38556 22372 38612 22382
rect 38332 22260 38388 22270
rect 38388 22204 38500 22260
rect 38332 22166 38388 22204
rect 37772 21028 37828 21038
rect 37996 21028 38052 21038
rect 37772 21026 38052 21028
rect 37772 20974 37774 21026
rect 37826 20974 37998 21026
rect 38050 20974 38052 21026
rect 37772 20972 38052 20974
rect 37772 20962 37828 20972
rect 37996 20962 38052 20972
rect 37660 20690 37716 20702
rect 37660 20638 37662 20690
rect 37714 20638 37716 20690
rect 37660 20244 37716 20638
rect 38220 20578 38276 20590
rect 38220 20526 38222 20578
rect 38274 20526 38276 20578
rect 38220 20468 38276 20526
rect 37996 20412 38276 20468
rect 37884 20244 37940 20254
rect 37660 20242 37940 20244
rect 37660 20190 37886 20242
rect 37938 20190 37940 20242
rect 37660 20188 37940 20190
rect 37884 20178 37940 20188
rect 37548 19814 37604 19852
rect 37884 20020 37940 20030
rect 37548 19572 37604 19582
rect 37548 19458 37604 19516
rect 37548 19406 37550 19458
rect 37602 19406 37604 19458
rect 37548 19394 37604 19406
rect 37436 18610 37492 18620
rect 37548 18788 37604 18798
rect 37548 15540 37604 18732
rect 37660 18676 37716 18686
rect 37660 18450 37716 18620
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 37660 18386 37716 18398
rect 37884 18676 37940 19964
rect 37996 19796 38052 20412
rect 38108 20132 38164 20142
rect 38108 20038 38164 20076
rect 38220 20020 38276 20030
rect 38220 19926 38276 19964
rect 37996 19730 38052 19740
rect 38332 19236 38388 19246
rect 38332 19142 38388 19180
rect 37884 17556 37940 18620
rect 38108 19010 38164 19022
rect 38108 18958 38110 19010
rect 38162 18958 38164 19010
rect 38108 18452 38164 18958
rect 38220 19012 38276 19050
rect 38220 18946 38276 18956
rect 38220 18788 38276 18798
rect 38220 18674 38276 18732
rect 38220 18622 38222 18674
rect 38274 18622 38276 18674
rect 38220 18610 38276 18622
rect 38332 18676 38388 18686
rect 38332 18618 38388 18620
rect 38332 18566 38334 18618
rect 38386 18566 38388 18618
rect 38332 18554 38388 18566
rect 38444 18452 38500 22204
rect 38556 22258 38612 22316
rect 38556 22206 38558 22258
rect 38610 22206 38612 22258
rect 38556 22194 38612 22206
rect 38668 22036 38724 22540
rect 38612 21980 38724 22036
rect 38612 21924 38668 21980
rect 38556 21868 38668 21924
rect 38556 21026 38612 21868
rect 38556 20974 38558 21026
rect 38610 20974 38612 21026
rect 38556 20962 38612 20974
rect 39004 20916 39060 24108
rect 39228 24050 39284 24108
rect 39228 23998 39230 24050
rect 39282 23998 39284 24050
rect 39228 23986 39284 23998
rect 39340 23156 39396 23166
rect 39340 22372 39396 23100
rect 39452 22596 39508 24780
rect 39676 23938 39732 24892
rect 39900 25060 39956 25070
rect 39788 24724 39844 24734
rect 39788 24630 39844 24668
rect 39676 23886 39678 23938
rect 39730 23886 39732 23938
rect 39676 23154 39732 23886
rect 39676 23102 39678 23154
rect 39730 23102 39732 23154
rect 39676 23090 39732 23102
rect 39788 23492 39844 23502
rect 39452 22530 39508 22540
rect 39564 22930 39620 22942
rect 39564 22878 39566 22930
rect 39618 22878 39620 22930
rect 39452 22372 39508 22382
rect 39340 22370 39508 22372
rect 39340 22318 39454 22370
rect 39506 22318 39508 22370
rect 39340 22316 39508 22318
rect 39340 21924 39396 22316
rect 39452 22306 39508 22316
rect 39340 21858 39396 21868
rect 39116 20916 39172 20926
rect 39004 20860 39116 20916
rect 38668 20578 38724 20590
rect 38668 20526 38670 20578
rect 38722 20526 38724 20578
rect 38668 20356 38724 20526
rect 38556 20300 38724 20356
rect 38556 20020 38612 20300
rect 39004 20244 39060 20860
rect 39116 20822 39172 20860
rect 38668 20188 39060 20244
rect 38668 20186 38724 20188
rect 38668 20134 38670 20186
rect 38722 20134 38724 20186
rect 38668 20122 38724 20134
rect 38556 19954 38612 19964
rect 38780 20020 38836 20030
rect 38780 19926 38836 19964
rect 39340 20020 39396 20030
rect 39564 20020 39620 22878
rect 39788 22258 39844 23436
rect 39788 22206 39790 22258
rect 39842 22206 39844 22258
rect 39788 22194 39844 22206
rect 39788 20916 39844 20926
rect 39788 20356 39844 20860
rect 39788 20130 39844 20300
rect 39788 20078 39790 20130
rect 39842 20078 39844 20130
rect 39788 20066 39844 20078
rect 39900 20132 39956 25004
rect 40012 24836 40068 24846
rect 40012 22484 40068 24780
rect 40012 22390 40068 22428
rect 39900 20066 39956 20076
rect 39340 20018 39732 20020
rect 39340 19966 39342 20018
rect 39394 19966 39732 20018
rect 39340 19964 39732 19966
rect 39340 19954 39396 19964
rect 38668 19794 38724 19806
rect 38668 19742 38670 19794
rect 38722 19742 38724 19794
rect 38668 19236 38724 19742
rect 39564 19348 39620 19358
rect 39004 19236 39060 19246
rect 38668 19234 39060 19236
rect 38668 19182 38670 19234
rect 38722 19182 39006 19234
rect 39058 19182 39060 19234
rect 38668 19180 39060 19182
rect 38668 19170 38724 19180
rect 39004 19170 39060 19180
rect 38668 18676 38724 18686
rect 39228 18676 39284 18686
rect 38724 18620 38836 18676
rect 38668 18610 38724 18620
rect 38780 18562 38836 18620
rect 38780 18510 38782 18562
rect 38834 18510 38836 18562
rect 38780 18498 38836 18510
rect 38108 18386 38164 18396
rect 38332 18396 38500 18452
rect 38668 18450 38724 18462
rect 38668 18398 38670 18450
rect 38722 18398 38724 18450
rect 38220 18228 38276 18238
rect 38332 18228 38388 18396
rect 38220 18226 38388 18228
rect 38220 18174 38222 18226
rect 38274 18174 38388 18226
rect 38220 18172 38388 18174
rect 38668 18228 38724 18398
rect 39004 18452 39060 18462
rect 39004 18358 39060 18396
rect 38220 18162 38276 18172
rect 38668 18162 38724 18172
rect 38780 18340 38836 18350
rect 37884 17462 37940 17500
rect 38556 18004 38612 18014
rect 38780 18004 38836 18284
rect 38332 17444 38388 17454
rect 38332 17350 38388 17388
rect 38556 17444 38612 17948
rect 37100 15260 37380 15316
rect 37436 15316 37492 15326
rect 36876 14466 36932 14476
rect 36988 15204 37044 15214
rect 36876 14308 36932 14318
rect 36876 14214 36932 14252
rect 35308 13020 35700 13076
rect 36092 14196 36148 14206
rect 35308 12962 35364 13020
rect 35308 12910 35310 12962
rect 35362 12910 35364 12962
rect 35308 12898 35364 12910
rect 36092 12850 36148 14140
rect 36988 13972 37044 15148
rect 37100 14418 37156 15260
rect 37436 15222 37492 15260
rect 37548 15148 37604 15484
rect 37996 15540 38052 15550
rect 37772 15316 37828 15326
rect 37772 15222 37828 15260
rect 37548 15092 37716 15148
rect 37100 14366 37102 14418
rect 37154 14366 37156 14418
rect 37100 14196 37156 14366
rect 37100 14130 37156 14140
rect 37212 14532 37268 14542
rect 37100 13972 37156 13982
rect 36988 13970 37156 13972
rect 36988 13918 37102 13970
rect 37154 13918 37156 13970
rect 36988 13916 37156 13918
rect 37100 13906 37156 13916
rect 36316 13858 36372 13870
rect 36316 13806 36318 13858
rect 36370 13806 36372 13858
rect 36204 13412 36260 13422
rect 36204 12962 36260 13356
rect 36204 12910 36206 12962
rect 36258 12910 36260 12962
rect 36204 12898 36260 12910
rect 36092 12798 36094 12850
rect 36146 12798 36148 12850
rect 36092 12786 36148 12798
rect 35868 12738 35924 12750
rect 35868 12686 35870 12738
rect 35922 12686 35924 12738
rect 35532 12292 35588 12302
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11452 35476 11508
rect 35028 10668 35140 10724
rect 34972 10658 35028 10668
rect 34748 10610 34804 10622
rect 34748 10558 34750 10610
rect 34802 10558 34804 10610
rect 33628 9874 33684 9884
rect 34188 10500 34244 10510
rect 34188 9938 34244 10444
rect 34188 9886 34190 9938
rect 34242 9886 34244 9938
rect 33516 9044 33572 9054
rect 33180 6514 33236 6524
rect 33404 8036 33460 8046
rect 33404 7698 33460 7980
rect 33404 7646 33406 7698
rect 33458 7646 33460 7698
rect 33404 6578 33460 7646
rect 33516 7698 33572 8988
rect 34188 8260 34244 9886
rect 34748 9940 34804 10558
rect 34972 10500 35028 10510
rect 34860 9940 34916 9950
rect 34748 9938 34916 9940
rect 34748 9886 34862 9938
rect 34914 9886 34916 9938
rect 34748 9884 34916 9886
rect 34524 9714 34580 9726
rect 34524 9662 34526 9714
rect 34578 9662 34580 9714
rect 34524 9156 34580 9662
rect 34860 9604 34916 9884
rect 34972 9826 35028 10444
rect 34972 9774 34974 9826
rect 35026 9774 35028 9826
rect 34972 9762 35028 9774
rect 34860 9548 35028 9604
rect 34748 9156 34804 9166
rect 34524 9154 34804 9156
rect 34524 9102 34750 9154
rect 34802 9102 34804 9154
rect 34524 9100 34804 9102
rect 34748 9090 34804 9100
rect 34860 8930 34916 8942
rect 34860 8878 34862 8930
rect 34914 8878 34916 8930
rect 34524 8484 34580 8494
rect 34412 8260 34468 8270
rect 34188 8258 34412 8260
rect 34188 8206 34190 8258
rect 34242 8206 34412 8258
rect 34188 8204 34412 8206
rect 34188 8166 34244 8204
rect 34412 8194 34468 8204
rect 34524 8146 34580 8428
rect 34748 8260 34804 8270
rect 34860 8260 34916 8878
rect 34748 8258 34916 8260
rect 34748 8206 34750 8258
rect 34802 8206 34916 8258
rect 34748 8204 34916 8206
rect 34748 8194 34804 8204
rect 34524 8094 34526 8146
rect 34578 8094 34580 8146
rect 34524 8082 34580 8094
rect 34636 8036 34692 8046
rect 34636 7942 34692 7980
rect 33516 7646 33518 7698
rect 33570 7646 33572 7698
rect 33516 7634 33572 7646
rect 33628 7476 33684 7486
rect 34972 7476 35028 9548
rect 35084 9042 35140 10668
rect 35420 10610 35476 11452
rect 35420 10558 35422 10610
rect 35474 10558 35476 10610
rect 35420 10500 35476 10558
rect 35532 10612 35588 12236
rect 35644 10724 35700 10734
rect 35644 10630 35700 10668
rect 35532 10546 35588 10556
rect 35420 10434 35476 10444
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35084 8990 35086 9042
rect 35138 8990 35140 9042
rect 35084 8978 35140 8990
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35084 8484 35140 8522
rect 35084 8418 35140 8428
rect 35868 8428 35924 12686
rect 36316 12292 36372 13806
rect 37212 13860 37268 14476
rect 37660 13970 37716 15092
rect 37660 13918 37662 13970
rect 37714 13918 37716 13970
rect 37660 13906 37716 13918
rect 37548 13860 37604 13870
rect 37212 13858 37548 13860
rect 37212 13806 37214 13858
rect 37266 13806 37548 13858
rect 37212 13804 37548 13806
rect 37212 13794 37268 13804
rect 37548 13766 37604 13804
rect 36652 13746 36708 13758
rect 36652 13694 36654 13746
rect 36706 13694 36708 13746
rect 36652 13412 36708 13694
rect 36540 12404 36596 12414
rect 36652 12404 36708 13356
rect 36540 12402 36708 12404
rect 36540 12350 36542 12402
rect 36594 12350 36708 12402
rect 36540 12348 36708 12350
rect 36876 13746 36932 13758
rect 36876 13694 36878 13746
rect 36930 13694 36932 13746
rect 36540 12338 36596 12348
rect 36204 12236 36372 12292
rect 36204 11284 36260 12236
rect 36204 11190 36260 11228
rect 36316 11396 36372 11406
rect 36316 11282 36372 11340
rect 36316 11230 36318 11282
rect 36370 11230 36372 11282
rect 36316 11218 36372 11230
rect 36540 11170 36596 11182
rect 36540 11118 36542 11170
rect 36594 11118 36596 11170
rect 36540 9044 36596 11118
rect 36764 10500 36820 10510
rect 36764 10406 36820 10444
rect 36540 8978 36596 8988
rect 36876 8428 36932 13694
rect 37660 13522 37716 13534
rect 37660 13470 37662 13522
rect 37714 13470 37716 13522
rect 37100 13412 37156 13422
rect 37100 13074 37156 13356
rect 37100 13022 37102 13074
rect 37154 13022 37156 13074
rect 37100 13010 37156 13022
rect 37324 11396 37380 11406
rect 37324 11302 37380 11340
rect 37548 10612 37604 10622
rect 37548 10518 37604 10556
rect 37436 9716 37492 9726
rect 37436 9622 37492 9660
rect 37660 9268 37716 13470
rect 37772 11394 37828 11406
rect 37772 11342 37774 11394
rect 37826 11342 37828 11394
rect 37772 9716 37828 11342
rect 37996 10498 38052 15484
rect 38444 15428 38500 15438
rect 38220 15426 38500 15428
rect 38220 15374 38446 15426
rect 38498 15374 38500 15426
rect 38220 15372 38500 15374
rect 38220 14530 38276 15372
rect 38444 15362 38500 15372
rect 38556 15428 38612 17388
rect 38332 15202 38388 15214
rect 38332 15150 38334 15202
rect 38386 15150 38388 15202
rect 38332 14644 38388 15150
rect 38332 14550 38388 14588
rect 38220 14478 38222 14530
rect 38274 14478 38276 14530
rect 38220 14420 38276 14478
rect 38220 14354 38276 14364
rect 38220 13972 38276 13982
rect 38108 13860 38164 13870
rect 38108 13766 38164 13804
rect 38220 11396 38276 13916
rect 38444 13746 38500 13758
rect 38444 13694 38446 13746
rect 38498 13694 38500 13746
rect 38444 13636 38500 13694
rect 38444 13570 38500 13580
rect 38220 11330 38276 11340
rect 37996 10446 37998 10498
rect 38050 10446 38052 10498
rect 37996 10434 38052 10446
rect 37996 9828 38052 9838
rect 38556 9828 38612 15372
rect 38668 17948 38836 18004
rect 38668 13412 38724 17948
rect 38892 17892 38948 17902
rect 38780 17668 38836 17678
rect 38780 17108 38836 17612
rect 38780 17014 38836 17052
rect 38780 15316 38836 15326
rect 38780 13748 38836 15260
rect 38780 13654 38836 13692
rect 38668 13346 38724 13356
rect 38780 11956 38836 11966
rect 38780 10724 38836 11900
rect 38892 10836 38948 17836
rect 39228 17780 39284 18620
rect 39452 18452 39508 18462
rect 39452 18358 39508 18396
rect 39564 18228 39620 19292
rect 39676 19236 39732 19964
rect 39676 19142 39732 19180
rect 39900 19906 39956 19918
rect 39900 19854 39902 19906
rect 39954 19854 39956 19906
rect 39900 19236 39956 19854
rect 39004 17668 39060 17678
rect 39004 17574 39060 17612
rect 39116 17556 39172 17566
rect 39228 17556 39284 17724
rect 39340 18172 39620 18228
rect 39788 19122 39844 19134
rect 39788 19070 39790 19122
rect 39842 19070 39844 19122
rect 39340 17666 39396 18172
rect 39676 17780 39732 17790
rect 39676 17686 39732 17724
rect 39340 17614 39342 17666
rect 39394 17614 39396 17666
rect 39340 17602 39396 17614
rect 39116 17554 39284 17556
rect 39116 17502 39118 17554
rect 39170 17502 39284 17554
rect 39116 17500 39284 17502
rect 39788 17556 39844 19070
rect 39900 18450 39956 19180
rect 39900 18398 39902 18450
rect 39954 18398 39956 18450
rect 39900 18386 39956 18398
rect 40124 18340 40180 27356
rect 40572 26908 40628 29484
rect 40684 29428 40740 30044
rect 40684 29362 40740 29372
rect 40908 29764 40964 29774
rect 40908 29426 40964 29708
rect 40908 29374 40910 29426
rect 40962 29374 40964 29426
rect 40908 29362 40964 29374
rect 40460 26852 40628 26908
rect 40796 28418 40852 28430
rect 40796 28366 40798 28418
rect 40850 28366 40852 28418
rect 40796 26908 40852 28366
rect 41020 27412 41076 31836
rect 41132 31826 41188 31836
rect 41356 31892 41412 31902
rect 41356 31798 41412 31836
rect 41244 30772 41300 30782
rect 41132 30212 41188 30222
rect 41132 30118 41188 30156
rect 41244 29650 41300 30716
rect 41244 29598 41246 29650
rect 41298 29598 41300 29650
rect 41244 29586 41300 29598
rect 41356 30100 41412 30110
rect 41356 29538 41412 30044
rect 41468 29876 41524 32732
rect 41692 32694 41748 32732
rect 41692 31556 41748 31566
rect 41580 31554 41748 31556
rect 41580 31502 41694 31554
rect 41746 31502 41748 31554
rect 41580 31500 41748 31502
rect 41580 30994 41636 31500
rect 41692 31490 41748 31500
rect 41580 30942 41582 30994
rect 41634 30942 41636 30994
rect 41580 30098 41636 30942
rect 41804 30994 41860 36988
rect 42252 35308 42308 39006
rect 42364 38612 42420 46396
rect 42476 46114 42532 46508
rect 42476 46062 42478 46114
rect 42530 46062 42532 46114
rect 42476 46050 42532 46062
rect 42588 44772 42644 46620
rect 42700 46610 42756 46620
rect 42812 46116 42868 46126
rect 42924 46116 42980 48300
rect 43036 48290 43092 48300
rect 42812 46114 42980 46116
rect 42812 46062 42814 46114
rect 42866 46062 42980 46114
rect 42812 46060 42980 46062
rect 42812 46050 42868 46060
rect 42588 44706 42644 44716
rect 43260 45892 43316 45902
rect 42588 44548 42644 44558
rect 42588 44322 42644 44492
rect 43260 44546 43316 45836
rect 43260 44494 43262 44546
rect 43314 44494 43316 44546
rect 43260 44482 43316 44494
rect 43372 44548 43428 52780
rect 43484 50708 43540 50718
rect 43484 50594 43540 50652
rect 43484 50542 43486 50594
rect 43538 50542 43540 50594
rect 43484 50530 43540 50542
rect 43596 49252 43652 54348
rect 43820 54310 43876 54348
rect 43820 53732 43876 53742
rect 44044 53732 44100 54684
rect 44156 54674 44212 54684
rect 44268 54516 44324 55244
rect 43820 53730 44100 53732
rect 43820 53678 43822 53730
rect 43874 53678 44100 53730
rect 43820 53676 44100 53678
rect 44156 54460 44324 54516
rect 43820 53666 43876 53676
rect 43820 51492 43876 51502
rect 43820 51398 43876 51436
rect 44044 51490 44100 51502
rect 44044 51438 44046 51490
rect 44098 51438 44100 51490
rect 44044 51380 44100 51438
rect 44044 51314 44100 51324
rect 43820 51268 43876 51278
rect 43820 50428 43876 51212
rect 43932 51266 43988 51278
rect 43932 51214 43934 51266
rect 43986 51214 43988 51266
rect 43932 50594 43988 51214
rect 43932 50542 43934 50594
rect 43986 50542 43988 50594
rect 43932 50530 43988 50542
rect 43820 50372 43988 50428
rect 43708 49810 43764 49822
rect 43708 49758 43710 49810
rect 43762 49758 43764 49810
rect 43708 49588 43764 49758
rect 43708 49522 43764 49532
rect 43484 49196 43652 49252
rect 43484 47682 43540 49196
rect 43820 49026 43876 49038
rect 43820 48974 43822 49026
rect 43874 48974 43876 49026
rect 43820 48356 43876 48974
rect 43820 48290 43876 48300
rect 43484 47630 43486 47682
rect 43538 47630 43540 47682
rect 43484 47618 43540 47630
rect 43820 46676 43876 46686
rect 43820 46582 43876 46620
rect 43708 46004 43764 46014
rect 43708 45910 43764 45948
rect 43372 44492 43540 44548
rect 42588 44270 42590 44322
rect 42642 44270 42644 44322
rect 42588 44258 42644 44270
rect 42700 44434 42756 44446
rect 42700 44382 42702 44434
rect 42754 44382 42756 44434
rect 42476 43652 42532 43662
rect 42700 43652 42756 44382
rect 42476 43650 42756 43652
rect 42476 43598 42478 43650
rect 42530 43598 42756 43650
rect 42476 43596 42756 43598
rect 42812 43764 42868 43774
rect 42812 43650 42868 43708
rect 42812 43598 42814 43650
rect 42866 43598 42868 43650
rect 42476 42756 42532 43596
rect 42812 43586 42868 43598
rect 43036 43540 43092 43550
rect 43036 43446 43092 43484
rect 43372 43316 43428 43326
rect 43148 43314 43428 43316
rect 43148 43262 43374 43314
rect 43426 43262 43428 43314
rect 43148 43260 43428 43262
rect 42588 42980 42644 42990
rect 42588 42978 42868 42980
rect 42588 42926 42590 42978
rect 42642 42926 42868 42978
rect 42588 42924 42868 42926
rect 42588 42914 42644 42924
rect 42476 42700 42756 42756
rect 42700 42642 42756 42700
rect 42700 42590 42702 42642
rect 42754 42590 42756 42642
rect 42700 42578 42756 42590
rect 42812 42644 42868 42924
rect 43036 42868 43092 42878
rect 43148 42868 43204 43260
rect 43372 43250 43428 43260
rect 43484 43092 43540 44492
rect 43036 42866 43204 42868
rect 43036 42814 43038 42866
rect 43090 42814 43204 42866
rect 43036 42812 43204 42814
rect 43372 43036 43540 43092
rect 43036 42802 43092 42812
rect 43260 42756 43316 42766
rect 43148 42754 43316 42756
rect 43148 42702 43262 42754
rect 43314 42702 43316 42754
rect 43148 42700 43316 42702
rect 43148 42644 43204 42700
rect 43260 42690 43316 42700
rect 42812 42588 43204 42644
rect 42476 42532 42532 42542
rect 42476 42438 42532 42476
rect 42700 41076 42756 41086
rect 42700 40626 42756 41020
rect 42700 40574 42702 40626
rect 42754 40574 42756 40626
rect 42700 40562 42756 40574
rect 42588 40178 42644 40190
rect 42588 40126 42590 40178
rect 42642 40126 42644 40178
rect 42476 39620 42532 39630
rect 42476 39284 42532 39564
rect 42588 39620 42644 40126
rect 43036 39730 43092 39742
rect 43036 39678 43038 39730
rect 43090 39678 43092 39730
rect 43036 39620 43092 39678
rect 42588 39618 42980 39620
rect 42588 39566 42590 39618
rect 42642 39566 42980 39618
rect 42588 39564 42980 39566
rect 42588 39554 42644 39564
rect 42476 39228 42756 39284
rect 42700 38946 42756 39228
rect 42924 39058 42980 39564
rect 43036 39554 43092 39564
rect 43372 39396 43428 43036
rect 43596 42530 43652 42542
rect 43596 42478 43598 42530
rect 43650 42478 43652 42530
rect 43596 40852 43652 42478
rect 43932 41188 43988 50372
rect 44156 49924 44212 54460
rect 44268 53844 44324 53854
rect 44268 53750 44324 53788
rect 44268 50484 44324 50522
rect 44268 50418 44324 50428
rect 44156 49868 44324 49924
rect 44156 49698 44212 49710
rect 44156 49646 44158 49698
rect 44210 49646 44212 49698
rect 44156 49026 44212 49646
rect 44268 49138 44324 49868
rect 44268 49086 44270 49138
rect 44322 49086 44324 49138
rect 44268 49074 44324 49086
rect 44156 48974 44158 49026
rect 44210 48974 44212 49026
rect 44156 48916 44212 48974
rect 44156 48860 44436 48916
rect 44380 48354 44436 48860
rect 44380 48302 44382 48354
rect 44434 48302 44436 48354
rect 44380 48290 44436 48302
rect 44492 48356 44548 48366
rect 44492 46786 44548 48300
rect 44492 46734 44494 46786
rect 44546 46734 44548 46786
rect 44492 46722 44548 46734
rect 44156 46676 44212 46686
rect 44044 46562 44100 46574
rect 44044 46510 44046 46562
rect 44098 46510 44100 46562
rect 44044 45892 44100 46510
rect 44044 45798 44100 45836
rect 44156 45778 44212 46620
rect 44604 45892 44660 55916
rect 44940 53844 44996 56590
rect 44940 53778 44996 53788
rect 45052 56980 45108 56990
rect 45052 50428 45108 56924
rect 45164 56866 45220 57148
rect 46060 57204 46116 57598
rect 46060 57138 46116 57148
rect 46172 57426 46228 57438
rect 46172 57374 46174 57426
rect 46226 57374 46228 57426
rect 45164 56814 45166 56866
rect 45218 56814 45220 56866
rect 45164 56802 45220 56814
rect 45500 57092 45556 57102
rect 45276 55076 45332 55086
rect 45276 54514 45332 55020
rect 45276 54462 45278 54514
rect 45330 54462 45332 54514
rect 44940 50372 45108 50428
rect 45164 53956 45220 53966
rect 44156 45726 44158 45778
rect 44210 45726 44212 45778
rect 44156 45714 44212 45726
rect 44268 45836 44660 45892
rect 44716 48242 44772 48254
rect 44716 48190 44718 48242
rect 44770 48190 44772 48242
rect 43596 40786 43652 40796
rect 43820 41132 43988 41188
rect 43708 40404 43764 40414
rect 43708 40310 43764 40348
rect 43596 40290 43652 40302
rect 43596 40238 43598 40290
rect 43650 40238 43652 40290
rect 43596 39956 43652 40238
rect 43484 39620 43540 39630
rect 43596 39620 43652 39900
rect 43484 39618 43652 39620
rect 43484 39566 43486 39618
rect 43538 39566 43652 39618
rect 43484 39564 43652 39566
rect 43484 39554 43540 39564
rect 43372 39340 43540 39396
rect 42924 39006 42926 39058
rect 42978 39006 42980 39058
rect 42924 38994 42980 39006
rect 42700 38894 42702 38946
rect 42754 38894 42756 38946
rect 42700 38882 42756 38894
rect 43372 38836 43428 38846
rect 43260 38834 43428 38836
rect 43260 38782 43374 38834
rect 43426 38782 43428 38834
rect 43260 38780 43428 38782
rect 43036 38724 43092 38734
rect 43260 38724 43316 38780
rect 43372 38770 43428 38780
rect 43036 38722 43316 38724
rect 43036 38670 43038 38722
rect 43090 38670 43316 38722
rect 43036 38668 43316 38670
rect 43484 38668 43540 39340
rect 43820 39172 43876 41132
rect 43932 40404 43988 40414
rect 43988 40348 44100 40404
rect 43932 40338 43988 40348
rect 44044 39620 44100 40348
rect 44156 39956 44212 39966
rect 44156 39842 44212 39900
rect 44156 39790 44158 39842
rect 44210 39790 44212 39842
rect 44156 39778 44212 39790
rect 43932 39564 44100 39620
rect 44156 39620 44212 39630
rect 43932 39506 43988 39564
rect 43932 39454 43934 39506
rect 43986 39454 43988 39506
rect 43932 39442 43988 39454
rect 44044 39394 44100 39406
rect 44044 39342 44046 39394
rect 44098 39342 44100 39394
rect 43820 39116 43988 39172
rect 43708 38948 43764 38958
rect 43708 38854 43764 38892
rect 43036 38658 43092 38668
rect 43372 38612 43428 38622
rect 43484 38612 43652 38668
rect 42364 38546 42420 38556
rect 43148 38610 43428 38612
rect 43148 38558 43374 38610
rect 43426 38558 43428 38610
rect 43148 38556 43428 38558
rect 43148 37492 43204 38556
rect 43372 38546 43428 38556
rect 42812 37436 43204 37492
rect 42364 35812 42420 35850
rect 42364 35746 42420 35756
rect 42476 35698 42532 35710
rect 42476 35646 42478 35698
rect 42530 35646 42532 35698
rect 41916 35252 42308 35308
rect 42364 35586 42420 35598
rect 42364 35534 42366 35586
rect 42418 35534 42420 35586
rect 41916 31892 41972 35252
rect 42028 34914 42084 34926
rect 42028 34862 42030 34914
rect 42082 34862 42084 34914
rect 42028 33684 42084 34862
rect 42028 33618 42084 33628
rect 42252 31892 42308 31902
rect 41972 31890 42308 31892
rect 41972 31838 42254 31890
rect 42306 31838 42308 31890
rect 41972 31836 42308 31838
rect 41916 31798 41972 31836
rect 42252 31826 42308 31836
rect 42364 31668 42420 35534
rect 42476 34916 42532 35646
rect 42476 34822 42532 34860
rect 42812 34356 42868 37436
rect 43036 37268 43092 37278
rect 43036 35810 43092 37212
rect 43372 37266 43428 37278
rect 43372 37214 43374 37266
rect 43426 37214 43428 37266
rect 43372 35812 43428 37214
rect 43484 37268 43540 37278
rect 43484 37154 43540 37212
rect 43484 37102 43486 37154
rect 43538 37102 43540 37154
rect 43484 37090 43540 37102
rect 43596 36596 43652 38612
rect 43596 36530 43652 36540
rect 43036 35758 43038 35810
rect 43090 35758 43092 35810
rect 43036 35746 43092 35758
rect 43148 35756 43428 35812
rect 43148 35476 43204 35756
rect 43372 35698 43428 35756
rect 43372 35646 43374 35698
rect 43426 35646 43428 35698
rect 43372 35634 43428 35646
rect 42924 34916 42980 34926
rect 43148 34916 43204 35420
rect 42924 34914 43204 34916
rect 42924 34862 42926 34914
rect 42978 34862 43204 34914
rect 42924 34860 43204 34862
rect 43260 35586 43316 35598
rect 43260 35534 43262 35586
rect 43314 35534 43316 35586
rect 42924 34850 42980 34860
rect 42812 34300 43204 34356
rect 42924 34130 42980 34142
rect 42924 34078 42926 34130
rect 42978 34078 42980 34130
rect 42700 33908 42756 33918
rect 42140 31612 42420 31668
rect 42476 33906 42756 33908
rect 42476 33854 42702 33906
rect 42754 33854 42756 33906
rect 42476 33852 42756 33854
rect 42476 33124 42532 33852
rect 42700 33842 42756 33852
rect 42924 33684 42980 34078
rect 42924 33618 42980 33628
rect 43148 33572 43204 34300
rect 43260 34130 43316 35534
rect 43932 35308 43988 39116
rect 44044 38948 44100 39342
rect 44044 38882 44100 38892
rect 44156 38668 44212 39564
rect 43820 35252 43988 35308
rect 44044 38612 44212 38668
rect 43260 34078 43262 34130
rect 43314 34078 43316 34130
rect 43260 34066 43316 34078
rect 43372 34802 43428 34814
rect 43372 34750 43374 34802
rect 43426 34750 43428 34802
rect 43372 34132 43428 34750
rect 43596 34354 43652 34366
rect 43596 34302 43598 34354
rect 43650 34302 43652 34354
rect 43484 34132 43540 34142
rect 43372 34130 43540 34132
rect 43372 34078 43486 34130
rect 43538 34078 43540 34130
rect 43372 34076 43540 34078
rect 43484 34066 43540 34076
rect 43148 33516 43540 33572
rect 42700 33348 42756 33358
rect 42700 33254 42756 33292
rect 43372 33346 43428 33358
rect 43372 33294 43374 33346
rect 43426 33294 43428 33346
rect 43372 33236 43428 33294
rect 42924 33180 43428 33236
rect 42812 33124 42868 33134
rect 41804 30942 41806 30994
rect 41858 30942 41860 30994
rect 41804 30210 41860 30942
rect 41804 30158 41806 30210
rect 41858 30158 41860 30210
rect 41804 30146 41860 30158
rect 42028 31444 42084 31454
rect 41580 30046 41582 30098
rect 41634 30046 41636 30098
rect 41580 30034 41636 30046
rect 41468 29820 41636 29876
rect 41356 29486 41358 29538
rect 41410 29486 41412 29538
rect 41356 29474 41412 29486
rect 41468 29428 41524 29438
rect 41468 29334 41524 29372
rect 41244 28980 41300 28990
rect 41244 28754 41300 28924
rect 41244 28702 41246 28754
rect 41298 28702 41300 28754
rect 41244 28690 41300 28702
rect 41020 27346 41076 27356
rect 41244 27300 41300 27310
rect 41244 27206 41300 27244
rect 40796 26852 40964 26908
rect 40460 25172 40516 26852
rect 40572 25394 40628 25406
rect 40572 25342 40574 25394
rect 40626 25342 40628 25394
rect 40572 25284 40628 25342
rect 40908 25284 40964 26852
rect 40572 25228 40964 25284
rect 40460 25116 40740 25172
rect 40348 24724 40404 24762
rect 40348 24658 40404 24668
rect 40348 24498 40404 24510
rect 40348 24446 40350 24498
rect 40402 24446 40404 24498
rect 40348 23938 40404 24446
rect 40348 23886 40350 23938
rect 40402 23886 40404 23938
rect 40348 23874 40404 23886
rect 40236 23492 40292 23502
rect 40236 23154 40292 23436
rect 40236 23102 40238 23154
rect 40290 23102 40292 23154
rect 40236 23090 40292 23102
rect 40572 22484 40628 22494
rect 40572 22390 40628 22428
rect 40460 22148 40516 22158
rect 40236 22146 40516 22148
rect 40236 22094 40462 22146
rect 40514 22094 40516 22146
rect 40236 22092 40516 22094
rect 40236 20020 40292 22092
rect 40460 22082 40516 22092
rect 40236 19926 40292 19964
rect 40236 19348 40292 19358
rect 40236 19234 40292 19292
rect 40236 19182 40238 19234
rect 40290 19182 40292 19234
rect 40236 19170 40292 19182
rect 40348 18564 40404 18574
rect 40348 18470 40404 18508
rect 40124 18274 40180 18284
rect 40348 18340 40404 18350
rect 40124 17780 40180 17790
rect 40124 17686 40180 17724
rect 39788 17500 39956 17556
rect 39116 17490 39172 17500
rect 39116 14532 39172 14542
rect 39788 14532 39844 14542
rect 39116 14438 39172 14476
rect 39676 14530 39844 14532
rect 39676 14478 39790 14530
rect 39842 14478 39844 14530
rect 39676 14476 39844 14478
rect 39452 13748 39508 13758
rect 39676 13748 39732 14476
rect 39788 14466 39844 14476
rect 39900 13860 39956 17500
rect 40124 15426 40180 15438
rect 40124 15374 40126 15426
rect 40178 15374 40180 15426
rect 40124 15148 40180 15374
rect 40348 15426 40404 18284
rect 40348 15374 40350 15426
rect 40402 15374 40404 15426
rect 40348 15362 40404 15374
rect 40124 15092 40516 15148
rect 39508 13746 39732 13748
rect 39508 13694 39678 13746
rect 39730 13694 39732 13746
rect 39508 13692 39732 13694
rect 39452 13682 39508 13692
rect 39676 13682 39732 13692
rect 39788 13804 39956 13860
rect 40012 14642 40068 14654
rect 40012 14590 40014 14642
rect 40066 14590 40068 14642
rect 39004 13524 39060 13534
rect 39004 13430 39060 13468
rect 39340 13522 39396 13534
rect 39340 13470 39342 13522
rect 39394 13470 39396 13522
rect 39340 12964 39396 13470
rect 39788 13412 39844 13804
rect 39900 13524 39956 13534
rect 40012 13524 40068 14590
rect 40460 14644 40516 15092
rect 40460 14550 40516 14588
rect 39956 13468 40068 13524
rect 40124 14532 40180 14542
rect 39900 13430 39956 13468
rect 39340 12898 39396 12908
rect 39452 13356 39844 13412
rect 38892 10780 39172 10836
rect 38780 10668 38948 10724
rect 38668 9828 38724 9838
rect 38556 9772 38668 9828
rect 37996 9734 38052 9772
rect 38668 9734 38724 9772
rect 37772 9650 37828 9660
rect 38108 9716 38164 9726
rect 38108 9622 38164 9660
rect 38332 9716 38388 9726
rect 38332 9622 38388 9660
rect 37212 9044 37268 9054
rect 37212 8950 37268 8988
rect 37660 9042 37716 9212
rect 38668 9268 38724 9278
rect 38668 9174 38724 9212
rect 37660 8990 37662 9042
rect 37714 8990 37716 9042
rect 37660 8978 37716 8990
rect 38444 9044 38500 9054
rect 38444 8950 38500 8988
rect 35868 8372 36148 8428
rect 35084 8260 35140 8270
rect 35084 8166 35140 8204
rect 33628 7474 34580 7476
rect 33628 7422 33630 7474
rect 33682 7422 34580 7474
rect 33628 7420 34580 7422
rect 33628 7410 33684 7420
rect 33404 6526 33406 6578
rect 33458 6526 33460 6578
rect 33404 6514 33460 6526
rect 33852 6802 33908 6814
rect 33852 6750 33854 6802
rect 33906 6750 33908 6802
rect 33852 6580 33908 6750
rect 34524 6802 34580 7420
rect 34972 7410 35028 7420
rect 35420 8146 35476 8158
rect 35420 8094 35422 8146
rect 35474 8094 35476 8146
rect 35420 7252 35476 8094
rect 34524 6750 34526 6802
rect 34578 6750 34580 6802
rect 34524 6738 34580 6750
rect 34972 7196 35476 7252
rect 35532 7476 35588 7486
rect 34412 6692 34468 6702
rect 34412 6598 34468 6636
rect 33852 6514 33908 6524
rect 34636 6580 34692 6590
rect 34636 6486 34692 6524
rect 33180 6132 33236 6142
rect 33180 6038 33236 6076
rect 33852 6132 33908 6142
rect 32508 6020 32564 6030
rect 32396 6018 32564 6020
rect 32396 5966 32510 6018
rect 32562 5966 32564 6018
rect 32396 5964 32564 5966
rect 32508 5954 32564 5964
rect 33852 6018 33908 6076
rect 33852 5966 33854 6018
rect 33906 5966 33908 6018
rect 33852 5954 33908 5966
rect 32172 5742 32174 5794
rect 32226 5742 32228 5794
rect 32172 5730 32228 5742
rect 33628 5908 33684 5918
rect 33628 5794 33684 5852
rect 33628 5742 33630 5794
rect 33682 5742 33684 5794
rect 33628 5730 33684 5742
rect 34972 5346 35028 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35308 6578 35364 6590
rect 35308 6526 35310 6578
rect 35362 6526 35364 6578
rect 35308 5908 35364 6526
rect 35420 6468 35476 6478
rect 35420 6374 35476 6412
rect 35532 6130 35588 7420
rect 36092 6804 36148 8372
rect 36092 6738 36148 6748
rect 36652 8372 36932 8428
rect 38108 8930 38164 8942
rect 38108 8878 38110 8930
rect 38162 8878 38164 8930
rect 38108 8428 38164 8878
rect 38780 8818 38836 8830
rect 38780 8766 38782 8818
rect 38834 8766 38836 8818
rect 38108 8372 38612 8428
rect 35532 6078 35534 6130
rect 35586 6078 35588 6130
rect 35532 6066 35588 6078
rect 35644 6578 35700 6590
rect 35644 6526 35646 6578
rect 35698 6526 35700 6578
rect 35532 5908 35588 5918
rect 35308 5906 35532 5908
rect 35308 5854 35310 5906
rect 35362 5854 35532 5906
rect 35308 5852 35532 5854
rect 35308 5842 35364 5852
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34972 5294 34974 5346
rect 35026 5294 35028 5346
rect 34972 5282 35028 5294
rect 35532 5234 35588 5852
rect 35532 5182 35534 5234
rect 35586 5182 35588 5234
rect 35532 5170 35588 5182
rect 35644 5796 35700 6526
rect 35868 6580 35924 6590
rect 35868 6578 36036 6580
rect 35868 6526 35870 6578
rect 35922 6526 36036 6578
rect 35868 6524 36036 6526
rect 35868 6514 35924 6524
rect 35644 5122 35700 5740
rect 35644 5070 35646 5122
rect 35698 5070 35700 5122
rect 35644 5058 35700 5070
rect 31948 4846 31950 4898
rect 32002 4846 32004 4898
rect 31948 4834 32004 4846
rect 35980 4562 36036 6524
rect 36428 6466 36484 6478
rect 36428 6414 36430 6466
rect 36482 6414 36484 6466
rect 36428 6132 36484 6414
rect 36428 6066 36484 6076
rect 36092 5908 36148 5918
rect 36652 5908 36708 8372
rect 36764 6804 36820 6814
rect 37772 6804 37828 6814
rect 36820 6748 36932 6804
rect 36764 6738 36820 6748
rect 36092 5814 36148 5852
rect 36204 5906 36708 5908
rect 36204 5854 36654 5906
rect 36706 5854 36708 5906
rect 36204 5852 36708 5854
rect 35980 4510 35982 4562
rect 36034 4510 36036 4562
rect 35980 4498 36036 4510
rect 35868 4450 35924 4462
rect 35868 4398 35870 4450
rect 35922 4398 35924 4450
rect 35868 4340 35924 4398
rect 36204 4340 36260 5852
rect 36652 5842 36708 5852
rect 36876 5796 36932 6748
rect 37660 6692 37716 6702
rect 37548 6690 37716 6692
rect 37548 6638 37662 6690
rect 37714 6638 37716 6690
rect 37548 6636 37716 6638
rect 36764 5794 36932 5796
rect 36764 5742 36878 5794
rect 36930 5742 36932 5794
rect 36764 5740 36932 5742
rect 36764 4452 36820 5740
rect 36876 5730 36932 5740
rect 37324 6578 37380 6590
rect 37324 6526 37326 6578
rect 37378 6526 37380 6578
rect 37324 6132 37380 6526
rect 37212 5236 37268 5246
rect 37324 5236 37380 6076
rect 37548 6020 37604 6636
rect 37660 6626 37716 6636
rect 37548 5906 37604 5964
rect 37548 5854 37550 5906
rect 37602 5854 37604 5906
rect 37548 5842 37604 5854
rect 37436 5796 37492 5806
rect 37436 5702 37492 5740
rect 37212 5234 37380 5236
rect 37212 5182 37214 5234
rect 37266 5182 37380 5234
rect 37212 5180 37380 5182
rect 37212 5170 37268 5180
rect 37772 5122 37828 6748
rect 38556 6690 38612 8372
rect 38780 6804 38836 8766
rect 38780 6738 38836 6748
rect 38556 6638 38558 6690
rect 38610 6638 38612 6690
rect 37884 6132 37940 6142
rect 37884 5906 37940 6076
rect 37884 5854 37886 5906
rect 37938 5854 37940 5906
rect 37884 5842 37940 5854
rect 37772 5070 37774 5122
rect 37826 5070 37828 5122
rect 37772 5058 37828 5070
rect 37996 5796 38052 5806
rect 37996 5122 38052 5740
rect 37996 5070 37998 5122
rect 38050 5070 38052 5122
rect 37996 5058 38052 5070
rect 38332 5124 38388 5134
rect 38556 5124 38612 6638
rect 38892 6466 38948 10668
rect 38892 6414 38894 6466
rect 38946 6414 38948 6466
rect 38892 6402 38948 6414
rect 39004 10610 39060 10622
rect 39004 10558 39006 10610
rect 39058 10558 39060 10610
rect 38892 6132 38948 6142
rect 38332 5122 38612 5124
rect 38332 5070 38334 5122
rect 38386 5070 38612 5122
rect 38332 5068 38612 5070
rect 38780 5682 38836 5694
rect 38780 5630 38782 5682
rect 38834 5630 38836 5682
rect 38332 5058 38388 5068
rect 38108 5012 38164 5022
rect 38108 4918 38164 4956
rect 38668 4564 38724 4574
rect 38780 4564 38836 5630
rect 38892 5234 38948 6076
rect 38892 5182 38894 5234
rect 38946 5182 38948 5234
rect 38892 5170 38948 5182
rect 39004 5236 39060 10558
rect 39116 6804 39172 10780
rect 39228 10386 39284 10398
rect 39228 10334 39230 10386
rect 39282 10334 39284 10386
rect 39228 9938 39284 10334
rect 39228 9886 39230 9938
rect 39282 9886 39284 9938
rect 39228 9874 39284 9886
rect 39340 9716 39396 9726
rect 39340 9622 39396 9660
rect 39452 8036 39508 13356
rect 39788 12964 39844 12974
rect 39788 12870 39844 12908
rect 40012 12964 40068 12974
rect 40124 12964 40180 14476
rect 40012 12962 40180 12964
rect 40012 12910 40014 12962
rect 40066 12910 40180 12962
rect 40012 12908 40180 12910
rect 40236 13522 40292 13534
rect 40236 13470 40238 13522
rect 40290 13470 40292 13522
rect 40236 12964 40292 13470
rect 40348 12964 40404 12974
rect 40236 12962 40404 12964
rect 40236 12910 40350 12962
rect 40402 12910 40404 12962
rect 40236 12908 40404 12910
rect 40012 12898 40068 12908
rect 40348 12898 40404 12908
rect 39900 12852 39956 12862
rect 39900 12758 39956 12796
rect 40124 9604 40180 9614
rect 40124 8258 40180 9548
rect 40124 8206 40126 8258
rect 40178 8206 40180 8258
rect 40124 8194 40180 8206
rect 39452 7980 39732 8036
rect 39564 6804 39620 6814
rect 39116 6802 39620 6804
rect 39116 6750 39566 6802
rect 39618 6750 39620 6802
rect 39116 6748 39620 6750
rect 39564 6738 39620 6748
rect 39564 6132 39620 6142
rect 39676 6132 39732 7980
rect 39900 8034 39956 8046
rect 39900 7982 39902 8034
rect 39954 7982 39956 8034
rect 39900 6578 39956 7982
rect 39900 6526 39902 6578
rect 39954 6526 39956 6578
rect 39900 6514 39956 6526
rect 39116 6076 39508 6132
rect 39116 6018 39172 6076
rect 39116 5966 39118 6018
rect 39170 5966 39172 6018
rect 39116 5954 39172 5966
rect 39340 5908 39396 5918
rect 39228 5906 39396 5908
rect 39228 5854 39342 5906
rect 39394 5854 39396 5906
rect 39228 5852 39396 5854
rect 39004 5180 39172 5236
rect 39004 5012 39060 5022
rect 38668 4562 38836 4564
rect 38668 4510 38670 4562
rect 38722 4510 38836 4562
rect 38668 4508 38836 4510
rect 38892 4956 39004 5012
rect 38892 4562 38948 4956
rect 39004 4918 39060 4956
rect 38892 4510 38894 4562
rect 38946 4510 38948 4562
rect 38668 4498 38724 4508
rect 38892 4498 38948 4510
rect 35868 4284 36260 4340
rect 36316 4396 36820 4452
rect 31500 4274 31556 4284
rect 36316 4228 36372 4396
rect 38780 4340 38836 4350
rect 39116 4340 39172 5180
rect 38780 4338 39172 4340
rect 38780 4286 38782 4338
rect 38834 4286 39172 4338
rect 38780 4284 39172 4286
rect 39228 4338 39284 5852
rect 39340 5842 39396 5852
rect 39452 5796 39508 6076
rect 39620 6076 39732 6132
rect 39564 6038 39620 6076
rect 39676 5906 39732 5918
rect 39676 5854 39678 5906
rect 39730 5854 39732 5906
rect 39676 5796 39732 5854
rect 39452 5740 39732 5796
rect 39228 4286 39230 4338
rect 39282 4286 39284 4338
rect 38780 4274 38836 4284
rect 39228 4274 39284 4286
rect 39452 4900 39508 4910
rect 39452 4340 39508 4844
rect 39564 4564 39620 4574
rect 39676 4564 39732 5740
rect 40460 5122 40516 5134
rect 40460 5070 40462 5122
rect 40514 5070 40516 5122
rect 40460 4900 40516 5070
rect 40460 4834 40516 4844
rect 39564 4562 39732 4564
rect 39564 4510 39566 4562
rect 39618 4510 39732 4562
rect 39564 4508 39732 4510
rect 40236 4788 40292 4798
rect 39564 4498 39620 4508
rect 39676 4340 39732 4350
rect 39452 4338 39732 4340
rect 39452 4286 39678 4338
rect 39730 4286 39732 4338
rect 39452 4284 39732 4286
rect 39676 4274 39732 4284
rect 30044 4114 30212 4116
rect 30044 4062 30046 4114
rect 30098 4062 30212 4114
rect 30044 4060 30212 4062
rect 36092 4172 36372 4228
rect 36092 4114 36148 4172
rect 36092 4062 36094 4114
rect 36146 4062 36148 4114
rect 30044 4050 30100 4060
rect 36092 4050 36148 4062
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 24892 3602 24948 3612
rect 40236 3666 40292 4732
rect 40236 3614 40238 3666
rect 40290 3614 40292 3666
rect 40236 3602 40292 3614
rect 40684 3668 40740 25116
rect 40796 23938 40852 23950
rect 40796 23886 40798 23938
rect 40850 23886 40852 23938
rect 40796 23378 40852 23886
rect 40908 23826 40964 25228
rect 40908 23774 40910 23826
rect 40962 23774 40964 23826
rect 40908 23762 40964 23774
rect 41020 25506 41076 25518
rect 41020 25454 41022 25506
rect 41074 25454 41076 25506
rect 41020 24724 41076 25454
rect 40796 23326 40798 23378
rect 40850 23326 40852 23378
rect 40796 23314 40852 23326
rect 40908 23492 40964 23502
rect 40908 22484 40964 23436
rect 41020 23378 41076 24668
rect 41020 23326 41022 23378
rect 41074 23326 41076 23378
rect 41020 23314 41076 23326
rect 41132 24836 41188 24846
rect 41132 23266 41188 24780
rect 41580 24724 41636 29820
rect 42028 25620 42084 31388
rect 42140 25844 42196 31612
rect 42476 31556 42532 33068
rect 42588 33122 42868 33124
rect 42588 33070 42814 33122
rect 42866 33070 42868 33122
rect 42588 33068 42868 33070
rect 42588 31892 42644 33068
rect 42812 33058 42868 33068
rect 42924 33122 42980 33180
rect 42924 33070 42926 33122
rect 42978 33070 42980 33122
rect 42700 32004 42756 32014
rect 42924 32004 42980 33070
rect 42700 32002 42980 32004
rect 42700 31950 42702 32002
rect 42754 31950 42980 32002
rect 42700 31948 42980 31950
rect 43036 33012 43092 33022
rect 42700 31938 42756 31948
rect 42588 31826 42644 31836
rect 42476 31490 42532 31500
rect 42588 31666 42644 31678
rect 42588 31614 42590 31666
rect 42642 31614 42644 31666
rect 42476 31106 42532 31118
rect 42476 31054 42478 31106
rect 42530 31054 42532 31106
rect 42252 30772 42308 30782
rect 42252 30678 42308 30716
rect 42364 30212 42420 30222
rect 42476 30212 42532 31054
rect 42588 30882 42644 31614
rect 42588 30830 42590 30882
rect 42642 30830 42644 30882
rect 42588 30818 42644 30830
rect 42420 30156 42532 30212
rect 42588 30212 42644 30222
rect 42364 30118 42420 30156
rect 42476 29986 42532 29998
rect 42476 29934 42478 29986
rect 42530 29934 42532 29986
rect 42476 26908 42532 29934
rect 42588 29538 42644 30156
rect 42588 29486 42590 29538
rect 42642 29486 42644 29538
rect 42588 29474 42644 29486
rect 42700 29428 42756 29438
rect 42700 29334 42756 29372
rect 42476 26852 42980 26908
rect 42140 25788 42420 25844
rect 42028 25564 42308 25620
rect 41692 25506 41748 25518
rect 41692 25454 41694 25506
rect 41746 25454 41748 25506
rect 41692 24836 41748 25454
rect 42140 25284 42196 25294
rect 42140 25190 42196 25228
rect 42252 25060 42308 25564
rect 42140 25004 42308 25060
rect 41692 24770 41748 24780
rect 41916 24836 41972 24846
rect 41580 24658 41636 24668
rect 41132 23214 41134 23266
rect 41186 23214 41188 23266
rect 41132 23202 41188 23214
rect 41244 24050 41300 24062
rect 41244 23998 41246 24050
rect 41298 23998 41300 24050
rect 41020 22484 41076 22494
rect 40908 22482 41076 22484
rect 40908 22430 41022 22482
rect 41074 22430 41076 22482
rect 40908 22428 41076 22430
rect 41020 22418 41076 22428
rect 41132 20578 41188 20590
rect 41132 20526 41134 20578
rect 41186 20526 41188 20578
rect 41020 20356 41076 20366
rect 41020 20242 41076 20300
rect 41020 20190 41022 20242
rect 41074 20190 41076 20242
rect 41020 20178 41076 20190
rect 41020 19348 41076 19358
rect 41020 19254 41076 19292
rect 40908 19236 40964 19246
rect 40908 19142 40964 19180
rect 41132 15148 41188 20526
rect 40796 15092 41188 15148
rect 40796 9826 40852 15092
rect 40908 14644 40964 14654
rect 40908 14550 40964 14588
rect 41132 14532 41188 14542
rect 41132 14438 41188 14476
rect 41244 13076 41300 23998
rect 41692 23938 41748 23950
rect 41692 23886 41694 23938
rect 41746 23886 41748 23938
rect 41580 23492 41636 23502
rect 41580 23378 41636 23436
rect 41580 23326 41582 23378
rect 41634 23326 41636 23378
rect 41580 23314 41636 23326
rect 41468 22484 41524 22494
rect 41468 21026 41524 22428
rect 41692 21812 41748 23886
rect 41916 23828 41972 24780
rect 41916 23826 42084 23828
rect 41916 23774 41918 23826
rect 41970 23774 42084 23826
rect 41916 23772 42084 23774
rect 41916 23762 41972 23772
rect 42028 22596 42084 23772
rect 41916 22540 42084 22596
rect 41916 22148 41972 22540
rect 42028 22372 42084 22382
rect 42140 22372 42196 25004
rect 42252 24836 42308 24846
rect 42364 24836 42420 25788
rect 42812 25508 42868 25518
rect 42252 24834 42420 24836
rect 42252 24782 42254 24834
rect 42306 24782 42420 24834
rect 42252 24780 42420 24782
rect 42476 25506 42868 25508
rect 42476 25454 42814 25506
rect 42866 25454 42868 25506
rect 42476 25452 42868 25454
rect 42476 25284 42532 25452
rect 42812 25442 42868 25452
rect 42252 22484 42308 24780
rect 42476 24722 42532 25228
rect 42924 24948 42980 26852
rect 42812 24892 42980 24948
rect 42476 24670 42478 24722
rect 42530 24670 42532 24722
rect 42476 24658 42532 24670
rect 42588 24836 42644 24846
rect 42588 22594 42644 24780
rect 42700 24612 42756 24622
rect 42700 23826 42756 24556
rect 42700 23774 42702 23826
rect 42754 23774 42756 23826
rect 42700 23762 42756 23774
rect 42588 22542 42590 22594
rect 42642 22542 42644 22594
rect 42588 22530 42644 22542
rect 42700 23604 42756 23614
rect 42252 22418 42308 22428
rect 42028 22370 42196 22372
rect 42028 22318 42030 22370
rect 42082 22318 42196 22370
rect 42028 22316 42196 22318
rect 42028 22306 42084 22316
rect 41916 22092 42084 22148
rect 41468 20974 41470 21026
rect 41522 20974 41524 21026
rect 41468 20962 41524 20974
rect 41580 21756 41748 21812
rect 41580 19458 41636 21756
rect 41580 19406 41582 19458
rect 41634 19406 41636 19458
rect 41580 19348 41636 19406
rect 41580 19282 41636 19292
rect 41692 20690 41748 20702
rect 41692 20638 41694 20690
rect 41746 20638 41748 20690
rect 41692 18564 41748 20638
rect 41580 17668 41636 17678
rect 41580 16882 41636 17612
rect 41580 16830 41582 16882
rect 41634 16830 41636 16882
rect 41580 16818 41636 16830
rect 41692 16770 41748 18508
rect 41804 19906 41860 19918
rect 41804 19854 41806 19906
rect 41858 19854 41860 19906
rect 41804 18340 41860 19854
rect 41804 18274 41860 18284
rect 42028 17668 42084 22092
rect 42140 20690 42196 22316
rect 42700 21812 42756 23548
rect 42252 21756 42700 21812
rect 42252 21698 42308 21756
rect 42700 21718 42756 21756
rect 42252 21646 42254 21698
rect 42306 21646 42308 21698
rect 42252 21634 42308 21646
rect 42700 21588 42756 21598
rect 42812 21588 42868 24892
rect 43036 24834 43092 32956
rect 43484 30212 43540 33516
rect 43596 33348 43652 34302
rect 43596 33254 43652 33292
rect 43484 30146 43540 30156
rect 43708 31892 43764 31902
rect 43484 29652 43540 29662
rect 43372 29538 43428 29550
rect 43372 29486 43374 29538
rect 43426 29486 43428 29538
rect 43372 28868 43428 29486
rect 43372 28802 43428 28812
rect 43484 28756 43540 29596
rect 43484 28662 43540 28700
rect 43596 29428 43652 29438
rect 43596 28420 43652 29372
rect 43708 28980 43764 31836
rect 43820 29204 43876 35252
rect 44044 32900 44100 38612
rect 44268 37604 44324 45836
rect 44380 45668 44436 45678
rect 44380 45666 44660 45668
rect 44380 45614 44382 45666
rect 44434 45614 44660 45666
rect 44380 45612 44660 45614
rect 44380 45602 44436 45612
rect 44604 44996 44660 45612
rect 44716 45218 44772 48190
rect 44716 45166 44718 45218
rect 44770 45166 44772 45218
rect 44716 45154 44772 45166
rect 44828 45218 44884 45230
rect 44828 45166 44830 45218
rect 44882 45166 44884 45218
rect 44828 44996 44884 45166
rect 44604 44940 44884 44996
rect 44380 42308 44436 42318
rect 44380 40292 44436 42252
rect 44940 41972 44996 50372
rect 45164 47908 45220 53900
rect 45276 53620 45332 54462
rect 45500 54292 45556 57036
rect 46172 55636 46228 57374
rect 45612 55580 46228 55636
rect 45612 55410 45668 55580
rect 45612 55358 45614 55410
rect 45666 55358 45668 55410
rect 45612 54514 45668 55358
rect 45836 55298 45892 55310
rect 45836 55246 45838 55298
rect 45890 55246 45892 55298
rect 45836 54852 45892 55246
rect 46172 55300 46228 55580
rect 46172 55234 46228 55244
rect 46172 55074 46228 55086
rect 46172 55022 46174 55074
rect 46226 55022 46228 55074
rect 46060 54852 46116 54862
rect 45836 54796 46060 54852
rect 46060 54786 46116 54796
rect 45612 54462 45614 54514
rect 45666 54462 45668 54514
rect 45612 54450 45668 54462
rect 45500 54236 45668 54292
rect 45500 53620 45556 53630
rect 45276 53618 45556 53620
rect 45276 53566 45502 53618
rect 45554 53566 45556 53618
rect 45276 53564 45556 53566
rect 45500 53554 45556 53564
rect 45612 50428 45668 54236
rect 45948 53842 46004 53854
rect 45948 53790 45950 53842
rect 46002 53790 46004 53842
rect 45500 50372 45668 50428
rect 45836 53620 45892 53630
rect 45500 49028 45556 50372
rect 45500 48962 45556 48972
rect 45612 50260 45668 50270
rect 45388 48132 45444 48142
rect 45164 47842 45220 47852
rect 45276 48076 45388 48132
rect 45164 46004 45220 46014
rect 45276 46004 45332 48076
rect 45388 48038 45444 48076
rect 45612 48130 45668 50204
rect 45836 48244 45892 53564
rect 45948 50594 46004 53790
rect 46060 53732 46116 53742
rect 46172 53732 46228 55022
rect 46060 53730 46228 53732
rect 46060 53678 46062 53730
rect 46114 53678 46228 53730
rect 46060 53676 46228 53678
rect 46284 54852 46340 54862
rect 46284 54514 46340 54796
rect 46284 54462 46286 54514
rect 46338 54462 46340 54514
rect 46060 53666 46116 53676
rect 46284 53620 46340 54462
rect 46172 53564 46340 53620
rect 46172 51380 46228 53564
rect 46284 51380 46340 51390
rect 46172 51324 46284 51380
rect 46284 51314 46340 51324
rect 45948 50542 45950 50594
rect 46002 50542 46004 50594
rect 45948 49698 46004 50542
rect 45948 49646 45950 49698
rect 46002 49646 46004 49698
rect 45948 49634 46004 49646
rect 46060 50706 46116 50718
rect 46060 50654 46062 50706
rect 46114 50654 46116 50706
rect 46060 49250 46116 50654
rect 46396 50428 46452 58268
rect 46508 58322 46564 59164
rect 46732 58772 46788 62132
rect 46508 58270 46510 58322
rect 46562 58270 46564 58322
rect 46508 58258 46564 58270
rect 46620 58716 46788 58772
rect 46508 55074 46564 55086
rect 46508 55022 46510 55074
rect 46562 55022 46564 55074
rect 46508 53730 46564 55022
rect 46620 54628 46676 58716
rect 46956 58434 47012 58446
rect 46956 58382 46958 58434
rect 47010 58382 47012 58434
rect 46732 58210 46788 58222
rect 46732 58158 46734 58210
rect 46786 58158 46788 58210
rect 46732 56196 46788 58158
rect 46844 57764 46900 57774
rect 46956 57764 47012 58382
rect 46900 57708 47012 57764
rect 46844 57670 46900 57708
rect 46732 56140 46900 56196
rect 46732 55972 46788 55982
rect 46732 55412 46788 55916
rect 46844 55860 46900 56140
rect 47068 56082 47124 56094
rect 47068 56030 47070 56082
rect 47122 56030 47124 56082
rect 47068 55972 47124 56030
rect 47068 55906 47124 55916
rect 46844 55804 47012 55860
rect 46732 55346 46788 55356
rect 46844 55298 46900 55310
rect 46844 55246 46846 55298
rect 46898 55246 46900 55298
rect 46732 54852 46788 54862
rect 46844 54852 46900 55246
rect 46788 54796 46900 54852
rect 46732 54786 46788 54796
rect 46844 54628 46900 54638
rect 46620 54626 46900 54628
rect 46620 54574 46846 54626
rect 46898 54574 46900 54626
rect 46620 54572 46900 54574
rect 46844 54562 46900 54572
rect 46508 53678 46510 53730
rect 46562 53678 46564 53730
rect 46508 53666 46564 53678
rect 46620 54180 46676 54190
rect 46620 51604 46676 54124
rect 46956 53956 47012 55804
rect 47068 55300 47124 55310
rect 47068 55206 47124 55244
rect 46956 53900 47124 53956
rect 46956 53730 47012 53742
rect 46956 53678 46958 53730
rect 47010 53678 47012 53730
rect 46956 53508 47012 53678
rect 47068 53732 47124 53900
rect 47068 53666 47124 53676
rect 46732 53452 46956 53508
rect 46732 53170 46788 53452
rect 46956 53442 47012 53452
rect 46732 53118 46734 53170
rect 46786 53118 46788 53170
rect 46732 53106 46788 53118
rect 46620 51602 47012 51604
rect 46620 51550 46622 51602
rect 46674 51550 47012 51602
rect 46620 51548 47012 51550
rect 46620 51538 46676 51548
rect 46284 50372 46452 50428
rect 46844 51380 46900 51390
rect 46284 49924 46340 50372
rect 46284 49858 46340 49868
rect 46060 49198 46062 49250
rect 46114 49198 46116 49250
rect 46060 49186 46116 49198
rect 46172 49810 46228 49822
rect 46172 49758 46174 49810
rect 46226 49758 46228 49810
rect 46172 49026 46228 49758
rect 46396 49812 46452 49822
rect 46396 49138 46452 49756
rect 46396 49086 46398 49138
rect 46450 49086 46452 49138
rect 46396 49074 46452 49086
rect 46172 48974 46174 49026
rect 46226 48974 46228 49026
rect 46172 48466 46228 48974
rect 46172 48414 46174 48466
rect 46226 48414 46228 48466
rect 46172 48402 46228 48414
rect 46732 49028 46788 49038
rect 46732 48466 46788 48972
rect 46732 48414 46734 48466
rect 46786 48414 46788 48466
rect 46732 48402 46788 48414
rect 45836 48188 46004 48244
rect 45612 48078 45614 48130
rect 45666 48078 45668 48130
rect 45220 45948 45332 46004
rect 45164 45910 45220 45948
rect 45052 45106 45108 45118
rect 45052 45054 45054 45106
rect 45106 45054 45108 45106
rect 45052 44996 45108 45054
rect 45052 44930 45108 44940
rect 45276 43428 45332 45948
rect 45612 45778 45668 48078
rect 45724 48132 45780 48142
rect 45780 48076 45892 48132
rect 45724 48066 45780 48076
rect 45836 48018 45892 48076
rect 45836 47966 45838 48018
rect 45890 47966 45892 48018
rect 45836 47954 45892 47966
rect 45612 45726 45614 45778
rect 45666 45726 45668 45778
rect 45612 43540 45668 45726
rect 45724 44996 45780 45006
rect 45724 44902 45780 44940
rect 45836 44884 45892 44894
rect 45836 43876 45892 44828
rect 45948 44436 46004 48188
rect 46620 47908 46676 47918
rect 46620 46900 46676 47852
rect 46620 46806 46676 46844
rect 46844 45666 46900 51324
rect 46956 51378 47012 51548
rect 46956 51326 46958 51378
rect 47010 51326 47012 51378
rect 46956 51314 47012 51326
rect 46956 49028 47012 49038
rect 46956 48934 47012 48972
rect 47180 48468 47236 48478
rect 47180 48374 47236 48412
rect 47292 48244 47348 79200
rect 48188 78036 48244 78046
rect 48188 76690 48244 77980
rect 48188 76638 48190 76690
rect 48242 76638 48244 76690
rect 48188 76626 48244 76638
rect 48188 75572 48244 75582
rect 48188 75478 48244 75516
rect 48188 73442 48244 73454
rect 48188 73390 48190 73442
rect 48242 73390 48244 73442
rect 48188 73108 48244 73390
rect 48188 73042 48244 73052
rect 48188 70754 48244 70766
rect 48188 70702 48190 70754
rect 48242 70702 48244 70754
rect 48188 70644 48244 70702
rect 48188 70578 48244 70588
rect 48188 68738 48244 68750
rect 48188 68686 48190 68738
rect 48242 68686 48244 68738
rect 48188 68180 48244 68686
rect 48188 68114 48244 68124
rect 48188 66050 48244 66062
rect 48188 65998 48190 66050
rect 48242 65998 48244 66050
rect 48188 65716 48244 65998
rect 48188 65650 48244 65660
rect 48188 64034 48244 64046
rect 48188 63982 48190 64034
rect 48242 63982 48244 64034
rect 48188 63252 48244 63982
rect 48188 63186 48244 63196
rect 48188 61346 48244 61358
rect 48188 61294 48190 61346
rect 48242 61294 48244 61346
rect 48188 60788 48244 61294
rect 48188 60722 48244 60732
rect 48076 58324 48132 58334
rect 48076 58230 48132 58268
rect 48076 55970 48132 55982
rect 48076 55918 48078 55970
rect 48130 55918 48132 55970
rect 48076 55860 48132 55918
rect 48076 55794 48132 55804
rect 47404 53732 47460 53742
rect 47404 50594 47460 53676
rect 48076 53620 48132 53630
rect 48076 53526 48132 53564
rect 48076 51266 48132 51278
rect 48076 51214 48078 51266
rect 48130 51214 48132 51266
rect 48076 50932 48132 51214
rect 48076 50866 48132 50876
rect 47404 50542 47406 50594
rect 47458 50542 47460 50594
rect 47404 50530 47460 50542
rect 47628 50706 47684 50718
rect 47628 50654 47630 50706
rect 47682 50654 47684 50706
rect 47516 49812 47572 49822
rect 47516 49718 47572 49756
rect 47292 48178 47348 48188
rect 47404 48354 47460 48366
rect 47404 48302 47406 48354
rect 47458 48302 47460 48354
rect 46956 46900 47012 46910
rect 46956 46674 47012 46844
rect 46956 46622 46958 46674
rect 47010 46622 47012 46674
rect 46956 46610 47012 46622
rect 46844 45614 46846 45666
rect 46898 45614 46900 45666
rect 46844 45602 46900 45614
rect 46956 45778 47012 45790
rect 46956 45726 46958 45778
rect 47010 45726 47012 45778
rect 45948 44342 46004 44380
rect 46508 44884 46564 44894
rect 46284 44212 46340 44222
rect 46284 44210 46452 44212
rect 46284 44158 46286 44210
rect 46338 44158 46452 44210
rect 46284 44156 46452 44158
rect 46284 44146 46340 44156
rect 45836 43820 46228 43876
rect 45948 43540 46004 43550
rect 45612 43538 46004 43540
rect 45612 43486 45950 43538
rect 46002 43486 46004 43538
rect 45612 43484 46004 43486
rect 45276 43334 45332 43372
rect 45836 42196 45892 43484
rect 45948 43474 46004 43484
rect 46172 42754 46228 43820
rect 46396 42868 46452 44156
rect 46508 44210 46564 44828
rect 46508 44158 46510 44210
rect 46562 44158 46564 44210
rect 46508 44146 46564 44158
rect 46620 44546 46676 44558
rect 46620 44494 46622 44546
rect 46674 44494 46676 44546
rect 46620 43764 46676 44494
rect 46956 44324 47012 45726
rect 46620 43698 46676 43708
rect 46844 44268 47012 44324
rect 47068 44436 47124 44446
rect 47068 44322 47124 44380
rect 47068 44270 47070 44322
rect 47122 44270 47124 44322
rect 46172 42702 46174 42754
rect 46226 42702 46228 42754
rect 46172 42690 46228 42702
rect 46284 42866 46452 42868
rect 46284 42814 46398 42866
rect 46450 42814 46452 42866
rect 46284 42812 46452 42814
rect 46284 42308 46340 42812
rect 46396 42802 46452 42812
rect 46508 43538 46564 43550
rect 46508 43486 46510 43538
rect 46562 43486 46564 43538
rect 46508 43428 46564 43486
rect 46620 43540 46676 43550
rect 46620 43446 46676 43484
rect 46844 43538 46900 44268
rect 47068 44258 47124 44270
rect 47404 43876 47460 48302
rect 47292 43820 47460 43876
rect 46844 43486 46846 43538
rect 46898 43486 46900 43538
rect 45836 42130 45892 42140
rect 46172 42252 46340 42308
rect 45724 42084 45780 42094
rect 44940 41906 44996 41916
rect 45388 42082 45780 42084
rect 45388 42030 45726 42082
rect 45778 42030 45780 42082
rect 45388 42028 45780 42030
rect 45388 41524 45444 42028
rect 45724 42018 45780 42028
rect 45836 41970 45892 41982
rect 45836 41918 45838 41970
rect 45890 41918 45892 41970
rect 45724 41748 45780 41758
rect 45724 41654 45780 41692
rect 45052 41468 45556 41524
rect 45052 41410 45108 41468
rect 45052 41358 45054 41410
rect 45106 41358 45108 41410
rect 45052 41346 45108 41358
rect 45388 41186 45444 41198
rect 45388 41134 45390 41186
rect 45442 41134 45444 41186
rect 45388 41076 45444 41134
rect 45164 40852 45220 40862
rect 45220 40796 45332 40852
rect 45164 40786 45220 40796
rect 44492 40516 44548 40526
rect 44492 40422 44548 40460
rect 45276 40402 45332 40796
rect 45388 40516 45444 41020
rect 45388 40450 45444 40460
rect 45276 40350 45278 40402
rect 45330 40350 45332 40402
rect 45052 40292 45108 40302
rect 44380 40236 44548 40292
rect 44380 39844 44436 39854
rect 44380 39172 44436 39788
rect 44492 39620 44548 40236
rect 44492 39554 44548 39564
rect 44828 40290 45108 40292
rect 44828 40238 45054 40290
rect 45106 40238 45108 40290
rect 44828 40236 45108 40238
rect 44828 39394 44884 40236
rect 45052 40226 45108 40236
rect 45052 39620 45108 39630
rect 45276 39620 45332 40350
rect 45052 39618 45332 39620
rect 45052 39566 45054 39618
rect 45106 39566 45332 39618
rect 45052 39564 45332 39566
rect 45500 39618 45556 41468
rect 45836 41186 45892 41918
rect 46172 41748 46228 42252
rect 46508 42196 46564 43372
rect 46844 42866 46900 43486
rect 47180 43540 47236 43550
rect 47180 43446 47236 43484
rect 46844 42814 46846 42866
rect 46898 42814 46900 42866
rect 46844 42802 46900 42814
rect 47068 43426 47124 43438
rect 47068 43374 47070 43426
rect 47122 43374 47124 43426
rect 46508 42140 46676 42196
rect 46172 41682 46228 41692
rect 46396 42084 46452 42094
rect 45836 41134 45838 41186
rect 45890 41134 45892 41186
rect 45836 41122 45892 41134
rect 45612 41074 45668 41086
rect 45612 41022 45614 41074
rect 45666 41022 45668 41074
rect 45612 40964 45668 41022
rect 46060 41074 46116 41086
rect 46060 41022 46062 41074
rect 46114 41022 46116 41074
rect 46060 40964 46116 41022
rect 46172 41076 46228 41086
rect 46172 40982 46228 41020
rect 45612 40908 46116 40964
rect 45948 40516 46004 40526
rect 46060 40516 46116 40908
rect 45948 40514 46116 40516
rect 45948 40462 45950 40514
rect 46002 40462 46116 40514
rect 45948 40460 46116 40462
rect 45948 40450 46004 40460
rect 45500 39566 45502 39618
rect 45554 39566 45556 39618
rect 45052 39554 45108 39564
rect 45500 39554 45556 39566
rect 44828 39342 44830 39394
rect 44882 39342 44884 39394
rect 44380 39116 44548 39172
rect 44044 32834 44100 32844
rect 44156 37548 44324 37604
rect 43932 30098 43988 30110
rect 43932 30046 43934 30098
rect 43986 30046 43988 30098
rect 43932 29652 43988 30046
rect 43932 29586 43988 29596
rect 44044 29986 44100 29998
rect 44044 29934 44046 29986
rect 44098 29934 44100 29986
rect 43932 29428 43988 29438
rect 44044 29428 44100 29934
rect 43988 29372 44100 29428
rect 43932 29334 43988 29372
rect 43820 29148 44100 29204
rect 43708 28924 43988 28980
rect 43708 28754 43764 28766
rect 43708 28702 43710 28754
rect 43762 28702 43764 28754
rect 43708 28644 43764 28702
rect 43708 28578 43764 28588
rect 43708 28420 43764 28430
rect 43596 28418 43764 28420
rect 43596 28366 43710 28418
rect 43762 28366 43764 28418
rect 43596 28364 43764 28366
rect 43708 28354 43764 28364
rect 43932 28196 43988 28924
rect 43708 28140 43988 28196
rect 43708 26292 43764 28140
rect 44044 28084 44100 29148
rect 43932 28028 44100 28084
rect 43708 26290 43876 26292
rect 43708 26238 43710 26290
rect 43762 26238 43876 26290
rect 43708 26236 43876 26238
rect 43708 26226 43764 26236
rect 43372 26180 43428 26190
rect 43372 26178 43652 26180
rect 43372 26126 43374 26178
rect 43426 26126 43652 26178
rect 43372 26124 43652 26126
rect 43372 26114 43428 26124
rect 43596 25620 43652 26124
rect 43708 25620 43764 25630
rect 43596 25618 43764 25620
rect 43596 25566 43710 25618
rect 43762 25566 43764 25618
rect 43596 25564 43764 25566
rect 43036 24782 43038 24834
rect 43090 24782 43092 24834
rect 42924 24724 42980 24734
rect 42924 23938 42980 24668
rect 43036 24612 43092 24782
rect 43148 25506 43204 25518
rect 43148 25454 43150 25506
rect 43202 25454 43204 25506
rect 43148 24836 43204 25454
rect 43148 24770 43204 24780
rect 43596 24724 43652 25564
rect 43708 25554 43764 25564
rect 43596 24658 43652 24668
rect 43820 24722 43876 26236
rect 43820 24670 43822 24722
rect 43874 24670 43876 24722
rect 43820 24658 43876 24670
rect 43036 24546 43092 24556
rect 43148 24610 43204 24622
rect 43148 24558 43150 24610
rect 43202 24558 43204 24610
rect 42924 23886 42926 23938
rect 42978 23886 42980 23938
rect 42924 23874 42980 23886
rect 43036 24050 43092 24062
rect 43036 23998 43038 24050
rect 43090 23998 43092 24050
rect 42140 20638 42142 20690
rect 42194 20638 42196 20690
rect 42140 20626 42196 20638
rect 42476 21586 42868 21588
rect 42476 21534 42702 21586
rect 42754 21534 42868 21586
rect 42476 21532 42868 21534
rect 42252 20020 42308 20030
rect 42476 20020 42532 21532
rect 42700 21522 42756 21532
rect 43036 20132 43092 23998
rect 42252 20018 42532 20020
rect 42252 19966 42254 20018
rect 42306 19966 42532 20018
rect 42252 19964 42532 19966
rect 42588 20076 43092 20132
rect 42140 19348 42196 19358
rect 42140 17778 42196 19292
rect 42140 17726 42142 17778
rect 42194 17726 42196 17778
rect 42140 17714 42196 17726
rect 42028 17574 42084 17612
rect 42140 16772 42196 16782
rect 41692 16718 41694 16770
rect 41746 16718 41748 16770
rect 41692 16706 41748 16718
rect 42028 16770 42196 16772
rect 42028 16718 42142 16770
rect 42194 16718 42196 16770
rect 42028 16716 42196 16718
rect 41916 15986 41972 15998
rect 41916 15934 41918 15986
rect 41970 15934 41972 15986
rect 41804 14644 41860 14654
rect 41916 14644 41972 15934
rect 42028 15148 42084 16716
rect 42140 16706 42196 16716
rect 42252 16548 42308 19964
rect 42140 16492 42308 16548
rect 42140 15986 42196 16492
rect 42252 16212 42308 16222
rect 42252 16210 42420 16212
rect 42252 16158 42254 16210
rect 42306 16158 42420 16210
rect 42252 16156 42420 16158
rect 42252 16146 42308 16156
rect 42140 15934 42142 15986
rect 42194 15934 42196 15986
rect 42140 15922 42196 15934
rect 42364 15986 42420 16156
rect 42364 15934 42366 15986
rect 42418 15934 42420 15986
rect 42364 15922 42420 15934
rect 42588 15148 42644 20076
rect 42700 19908 42756 19918
rect 43036 19908 43092 19918
rect 42700 19906 43092 19908
rect 42700 19854 42702 19906
rect 42754 19854 43038 19906
rect 43090 19854 43092 19906
rect 42700 19852 43092 19854
rect 42700 19842 42756 19852
rect 43036 19842 43092 19852
rect 43148 19684 43204 24558
rect 43708 24612 43764 24622
rect 43708 24162 43764 24556
rect 43708 24110 43710 24162
rect 43762 24110 43764 24162
rect 43708 24050 43764 24110
rect 43708 23998 43710 24050
rect 43762 23998 43764 24050
rect 43708 23986 43764 23998
rect 43820 24500 43876 24510
rect 43260 21812 43316 21822
rect 43260 20242 43316 21756
rect 43260 20190 43262 20242
rect 43314 20190 43316 20242
rect 43260 20178 43316 20190
rect 43484 21586 43540 21598
rect 43484 21534 43486 21586
rect 43538 21534 43540 21586
rect 43372 19794 43428 19806
rect 43372 19742 43374 19794
rect 43426 19742 43428 19794
rect 43148 19628 43316 19684
rect 42700 17556 42756 17566
rect 43036 17556 43092 17566
rect 42700 17554 43092 17556
rect 42700 17502 42702 17554
rect 42754 17502 43038 17554
rect 43090 17502 43092 17554
rect 42700 17500 43092 17502
rect 42700 17490 42756 17500
rect 43036 16770 43092 17500
rect 43260 17554 43316 19628
rect 43260 17502 43262 17554
rect 43314 17502 43316 17554
rect 43036 16718 43038 16770
rect 43090 16718 43092 16770
rect 43036 16706 43092 16718
rect 43148 17442 43204 17454
rect 43148 17390 43150 17442
rect 43202 17390 43204 17442
rect 43036 16212 43092 16222
rect 43036 16118 43092 16156
rect 42924 16098 42980 16110
rect 42924 16046 42926 16098
rect 42978 16046 42980 16098
rect 42812 15988 42868 15998
rect 42924 15988 42980 16046
rect 43148 16100 43204 17390
rect 43260 16882 43316 17502
rect 43260 16830 43262 16882
rect 43314 16830 43316 16882
rect 43260 16818 43316 16830
rect 43260 16324 43316 16334
rect 43372 16324 43428 19742
rect 43484 18340 43540 21534
rect 43484 18274 43540 18284
rect 43260 16322 43428 16324
rect 43260 16270 43262 16322
rect 43314 16270 43428 16322
rect 43260 16268 43428 16270
rect 43596 16658 43652 16670
rect 43596 16606 43598 16658
rect 43650 16606 43652 16658
rect 43260 16258 43316 16268
rect 43148 16044 43428 16100
rect 42812 15986 42980 15988
rect 42812 15934 42814 15986
rect 42866 15934 42980 15986
rect 42812 15932 42980 15934
rect 42812 15922 42868 15932
rect 43372 15148 43428 16044
rect 42028 15092 42196 15148
rect 41804 14642 41972 14644
rect 41804 14590 41806 14642
rect 41858 14590 41972 14642
rect 41804 14588 41972 14590
rect 41804 14578 41860 14588
rect 41020 13074 41300 13076
rect 41020 13022 41246 13074
rect 41298 13022 41300 13074
rect 41020 13020 41300 13022
rect 41020 12290 41076 13020
rect 41244 13010 41300 13020
rect 41692 12852 41748 12862
rect 41692 12758 41748 12796
rect 41020 12238 41022 12290
rect 41074 12238 41076 12290
rect 41020 12226 41076 12238
rect 41132 12068 41188 12078
rect 41468 12068 41524 12078
rect 41132 12066 41468 12068
rect 41132 12014 41134 12066
rect 41186 12014 41468 12066
rect 41132 12012 41468 12014
rect 41132 12002 41188 12012
rect 41468 11974 41524 12012
rect 41692 11956 41748 11966
rect 42028 11956 42084 11966
rect 41692 11862 41748 11900
rect 41916 11954 42084 11956
rect 41916 11902 42030 11954
rect 42082 11902 42084 11954
rect 41916 11900 42084 11902
rect 41916 11394 41972 11900
rect 42028 11890 42084 11900
rect 42140 11396 42196 15092
rect 42476 15092 42644 15148
rect 43148 15092 43428 15148
rect 41916 11342 41918 11394
rect 41970 11342 41972 11394
rect 41916 11330 41972 11342
rect 42028 11340 42196 11396
rect 42252 12852 42308 12862
rect 42252 11394 42308 12796
rect 42364 12068 42420 12078
rect 42364 11974 42420 12012
rect 42476 11732 42532 15092
rect 42588 12962 42644 12974
rect 42588 12910 42590 12962
rect 42642 12910 42644 12962
rect 42588 11956 42644 12910
rect 42924 11956 42980 11966
rect 42588 11862 42644 11900
rect 42700 11954 42980 11956
rect 42700 11902 42926 11954
rect 42978 11902 42980 11954
rect 42700 11900 42980 11902
rect 42252 11342 42254 11394
rect 42306 11342 42308 11394
rect 40796 9774 40798 9826
rect 40850 9774 40852 9826
rect 40796 9762 40852 9774
rect 40908 9604 40964 9614
rect 42028 9604 42084 11340
rect 42252 11330 42308 11342
rect 42364 11676 42532 11732
rect 42140 11170 42196 11182
rect 42140 11118 42142 11170
rect 42194 11118 42196 11170
rect 42140 9828 42196 11118
rect 42364 9940 42420 11676
rect 42700 11620 42756 11900
rect 42924 11890 42980 11900
rect 42476 11564 42756 11620
rect 42476 11394 42532 11564
rect 42476 11342 42478 11394
rect 42530 11342 42532 11394
rect 42476 11330 42532 11342
rect 43148 10612 43204 15092
rect 43596 14644 43652 16606
rect 43708 15876 43764 15886
rect 43708 14754 43764 15820
rect 43708 14702 43710 14754
rect 43762 14702 43764 14754
rect 43708 14690 43764 14702
rect 43484 14532 43540 14542
rect 43260 13076 43316 13086
rect 43260 12180 43316 13020
rect 43372 12180 43428 12190
rect 43260 12178 43428 12180
rect 43260 12126 43374 12178
rect 43426 12126 43428 12178
rect 43260 12124 43428 12126
rect 43372 12114 43428 12124
rect 43372 11956 43428 11966
rect 43484 11956 43540 14476
rect 43596 13636 43652 14588
rect 43820 14530 43876 24444
rect 43820 14478 43822 14530
rect 43874 14478 43876 14530
rect 43820 13858 43876 14478
rect 43820 13806 43822 13858
rect 43874 13806 43876 13858
rect 43820 13794 43876 13806
rect 43932 13860 43988 28028
rect 44156 26908 44212 37548
rect 44268 37380 44324 37390
rect 44268 37286 44324 37324
rect 44492 35308 44548 39116
rect 44828 37380 44884 39342
rect 44940 39394 44996 39406
rect 44940 39342 44942 39394
rect 44994 39342 44996 39394
rect 44940 38668 44996 39342
rect 45836 39396 45892 39406
rect 44940 38612 45220 38668
rect 44828 37314 44884 37324
rect 44380 35252 44548 35308
rect 44268 34130 44324 34142
rect 44268 34078 44270 34130
rect 44322 34078 44324 34130
rect 44268 33458 44324 34078
rect 44268 33406 44270 33458
rect 44322 33406 44324 33458
rect 44268 33394 44324 33406
rect 44380 30436 44436 35252
rect 45164 34916 45220 38612
rect 45388 37154 45444 37166
rect 45388 37102 45390 37154
rect 45442 37102 45444 37154
rect 45388 35812 45444 37102
rect 45612 36484 45668 36494
rect 45612 36390 45668 36428
rect 45388 35810 45780 35812
rect 45388 35758 45390 35810
rect 45442 35758 45780 35810
rect 45388 35756 45780 35758
rect 45388 35746 45444 35756
rect 45612 35588 45668 35598
rect 45500 35532 45612 35588
rect 45500 35474 45556 35532
rect 45612 35522 45668 35532
rect 45500 35422 45502 35474
rect 45554 35422 45556 35474
rect 45388 35028 45444 35038
rect 44828 34914 45220 34916
rect 44828 34862 45166 34914
rect 45218 34862 45220 34914
rect 44828 34860 45220 34862
rect 44828 34354 44884 34860
rect 45164 34850 45220 34860
rect 45276 35026 45444 35028
rect 45276 34974 45390 35026
rect 45442 34974 45444 35026
rect 45276 34972 45444 34974
rect 45276 34468 45332 34972
rect 45388 34962 45444 34972
rect 44828 34302 44830 34354
rect 44882 34302 44884 34354
rect 44828 34290 44884 34302
rect 44940 34412 45332 34468
rect 44492 34132 44548 34142
rect 44716 34132 44772 34142
rect 44940 34132 44996 34412
rect 45500 34354 45556 35422
rect 45724 34804 45780 35756
rect 45836 35028 45892 39340
rect 46060 37604 46116 37614
rect 45948 37548 46060 37604
rect 45948 37378 46004 37548
rect 46060 37538 46116 37548
rect 45948 37326 45950 37378
rect 46002 37326 46004 37378
rect 45948 37314 46004 37326
rect 46060 37268 46116 37278
rect 45948 37044 46004 37054
rect 45948 36706 46004 36988
rect 45948 36654 45950 36706
rect 46002 36654 46004 36706
rect 45948 36642 46004 36654
rect 46060 35586 46116 37212
rect 46396 36594 46452 42028
rect 46396 36542 46398 36594
rect 46450 36542 46452 36594
rect 46396 36530 46452 36542
rect 46508 41972 46564 41982
rect 46172 36484 46228 36494
rect 46228 36428 46340 36484
rect 46172 36390 46228 36428
rect 46060 35534 46062 35586
rect 46114 35534 46116 35586
rect 45836 34972 46004 35028
rect 45836 34804 45892 34814
rect 45724 34802 45892 34804
rect 45724 34750 45838 34802
rect 45890 34750 45892 34802
rect 45724 34748 45892 34750
rect 45836 34738 45892 34748
rect 45500 34302 45502 34354
rect 45554 34302 45556 34354
rect 45500 34290 45556 34302
rect 45052 34244 45108 34254
rect 45052 34150 45108 34188
rect 45724 34244 45780 34254
rect 45724 34150 45780 34188
rect 44492 34130 44996 34132
rect 44492 34078 44494 34130
rect 44546 34078 44718 34130
rect 44770 34078 44996 34130
rect 44492 34076 44996 34078
rect 45276 34130 45332 34142
rect 45276 34078 45278 34130
rect 45330 34078 45332 34130
rect 44492 34066 44548 34076
rect 44716 34066 44772 34076
rect 44380 30370 44436 30380
rect 44268 29988 44324 29998
rect 44268 29986 44772 29988
rect 44268 29934 44270 29986
rect 44322 29934 44772 29986
rect 44268 29932 44772 29934
rect 44268 29922 44324 29932
rect 44604 29652 44660 29662
rect 44604 29426 44660 29596
rect 44604 29374 44606 29426
rect 44658 29374 44660 29426
rect 44604 29362 44660 29374
rect 44716 28642 44772 29932
rect 45276 29538 45332 34078
rect 45276 29486 45278 29538
rect 45330 29486 45332 29538
rect 45276 29474 45332 29486
rect 45388 34018 45444 34030
rect 45388 33966 45390 34018
rect 45442 33966 45444 34018
rect 45388 29092 45444 33966
rect 45724 33124 45780 33134
rect 44716 28590 44718 28642
rect 44770 28590 44772 28642
rect 44716 28578 44772 28590
rect 45052 29036 45444 29092
rect 45612 33122 45780 33124
rect 45612 33070 45726 33122
rect 45778 33070 45780 33122
rect 45612 33068 45780 33070
rect 44044 26852 44212 26908
rect 45052 26908 45108 29036
rect 45164 28868 45220 28878
rect 45612 28868 45668 33068
rect 45724 33058 45780 33068
rect 45948 32788 46004 34972
rect 46060 33124 46116 35534
rect 46172 35698 46228 35710
rect 46172 35646 46174 35698
rect 46226 35646 46228 35698
rect 46172 35588 46228 35646
rect 46172 35522 46228 35532
rect 46284 34580 46340 36428
rect 46284 34514 46340 34524
rect 46508 34132 46564 41916
rect 46620 36484 46676 42140
rect 47068 42084 47124 43374
rect 46844 42028 47124 42084
rect 46844 37604 46900 42028
rect 47180 41188 47236 41198
rect 47292 41188 47348 43820
rect 47404 43652 47460 43662
rect 47404 43538 47460 43596
rect 47404 43486 47406 43538
rect 47458 43486 47460 43538
rect 47404 43474 47460 43486
rect 47180 41186 47348 41188
rect 47180 41134 47182 41186
rect 47234 41134 47348 41186
rect 47180 41132 47348 41134
rect 47180 41122 47236 41132
rect 46732 37548 46844 37604
rect 46732 36484 46788 37548
rect 46844 37538 46900 37548
rect 46844 37268 46900 37278
rect 46844 37174 46900 37212
rect 46844 36484 46900 36494
rect 46732 36482 46900 36484
rect 46732 36430 46846 36482
rect 46898 36430 46900 36482
rect 46732 36428 46900 36430
rect 46620 36418 46676 36428
rect 46844 36418 46900 36428
rect 46620 36258 46676 36270
rect 46620 36206 46622 36258
rect 46674 36206 46676 36258
rect 46620 35812 46676 36206
rect 46732 36258 46788 36270
rect 46732 36206 46734 36258
rect 46786 36206 46788 36258
rect 46732 36036 46788 36206
rect 46732 35980 47012 36036
rect 46844 35812 46900 35822
rect 46620 35810 46900 35812
rect 46620 35758 46846 35810
rect 46898 35758 46900 35810
rect 46620 35756 46900 35758
rect 46844 35746 46900 35756
rect 46956 35140 47012 35980
rect 46956 35084 47236 35140
rect 46620 34468 46676 34478
rect 46676 34412 46788 34468
rect 46620 34402 46676 34412
rect 46508 34066 46564 34076
rect 46620 34242 46676 34254
rect 46620 34190 46622 34242
rect 46674 34190 46676 34242
rect 46508 33906 46564 33918
rect 46508 33854 46510 33906
rect 46562 33854 46564 33906
rect 46172 33348 46228 33358
rect 46172 33254 46228 33292
rect 46508 33348 46564 33854
rect 46620 33908 46676 34190
rect 46620 33842 46676 33852
rect 46508 33282 46564 33292
rect 46732 33346 46788 34412
rect 47068 34356 47124 34366
rect 46732 33294 46734 33346
rect 46786 33294 46788 33346
rect 46060 33068 46228 33124
rect 45836 32732 46004 32788
rect 45724 30212 45780 30222
rect 45724 29314 45780 30156
rect 45724 29262 45726 29314
rect 45778 29262 45780 29314
rect 45724 29250 45780 29262
rect 45164 28530 45220 28812
rect 45500 28812 45668 28868
rect 45276 28756 45332 28766
rect 45276 28662 45332 28700
rect 45164 28478 45166 28530
rect 45218 28478 45220 28530
rect 45164 28466 45220 28478
rect 45388 28532 45444 28542
rect 45388 28438 45444 28476
rect 45164 26964 45220 26974
rect 45052 26852 45220 26908
rect 44044 26068 44100 26852
rect 45164 26402 45220 26852
rect 45164 26350 45166 26402
rect 45218 26350 45220 26402
rect 45164 26338 45220 26350
rect 44156 26180 44212 26190
rect 44156 26086 44212 26124
rect 44828 26180 44884 26190
rect 44828 26086 44884 26124
rect 45164 26180 45220 26190
rect 44044 26002 44100 26012
rect 45164 25508 45220 26124
rect 45052 25506 45220 25508
rect 45052 25454 45166 25506
rect 45218 25454 45220 25506
rect 45052 25452 45220 25454
rect 44044 24724 44100 24734
rect 44044 24630 44100 24668
rect 44380 24724 44436 24734
rect 44716 24724 44772 24734
rect 44380 24722 44772 24724
rect 44380 24670 44382 24722
rect 44434 24670 44718 24722
rect 44770 24670 44772 24722
rect 44380 24668 44772 24670
rect 44380 24658 44436 24668
rect 44716 24658 44772 24668
rect 44828 24724 44884 24734
rect 44156 24162 44212 24174
rect 44156 24110 44158 24162
rect 44210 24110 44212 24162
rect 44156 24050 44212 24110
rect 44156 23998 44158 24050
rect 44210 23998 44212 24050
rect 44156 23986 44212 23998
rect 44828 21698 44884 24668
rect 45052 24722 45108 25452
rect 45164 25442 45220 25452
rect 45388 25620 45444 25630
rect 45052 24670 45054 24722
rect 45106 24670 45108 24722
rect 45052 24658 45108 24670
rect 45388 24724 45444 25564
rect 45388 24630 45444 24668
rect 45164 24610 45220 24622
rect 45164 24558 45166 24610
rect 45218 24558 45220 24610
rect 45052 24500 45108 24510
rect 45164 24500 45220 24558
rect 45108 24444 45220 24500
rect 45052 24434 45108 24444
rect 44828 21646 44830 21698
rect 44882 21646 44884 21698
rect 44828 21634 44884 21646
rect 44940 24052 44996 24062
rect 44828 20692 44884 20702
rect 44828 20598 44884 20636
rect 44380 20018 44436 20030
rect 44380 19966 44382 20018
rect 44434 19966 44436 20018
rect 44380 18340 44436 19966
rect 44604 20018 44660 20030
rect 44604 19966 44606 20018
rect 44658 19966 44660 20018
rect 44492 19906 44548 19918
rect 44492 19854 44494 19906
rect 44546 19854 44548 19906
rect 44492 19460 44548 19854
rect 44492 19394 44548 19404
rect 44604 19236 44660 19966
rect 44940 19460 44996 23996
rect 45500 23604 45556 28812
rect 45612 26962 45668 26974
rect 45612 26910 45614 26962
rect 45666 26910 45668 26962
rect 45612 25732 45668 26910
rect 45724 26964 45780 27002
rect 45724 26898 45780 26908
rect 45836 25844 45892 32732
rect 46060 32676 46116 32686
rect 46060 32582 46116 32620
rect 46172 31892 46228 33068
rect 46732 32676 46788 33294
rect 46732 32610 46788 32620
rect 46844 33906 46900 33918
rect 46844 33854 46846 33906
rect 46898 33854 46900 33906
rect 46844 32452 46900 33854
rect 47068 33796 47124 34300
rect 47180 34242 47236 35084
rect 47180 34190 47182 34242
rect 47234 34190 47236 34242
rect 47180 34178 47236 34190
rect 47068 33346 47124 33740
rect 47068 33294 47070 33346
rect 47122 33294 47124 33346
rect 47068 33282 47124 33294
rect 47292 33908 47348 33918
rect 47292 32562 47348 33852
rect 47628 33796 47684 50654
rect 47740 49924 47796 49934
rect 47740 49830 47796 49868
rect 47964 49812 48020 49822
rect 47740 48804 47796 48814
rect 47740 48710 47796 48748
rect 47740 48356 47796 48366
rect 47740 48262 47796 48300
rect 47740 44098 47796 44110
rect 47740 44046 47742 44098
rect 47794 44046 47796 44098
rect 47740 43764 47796 44046
rect 47740 43698 47796 43708
rect 47964 38668 48020 49756
rect 48076 46562 48132 46574
rect 48076 46510 48078 46562
rect 48130 46510 48132 46562
rect 48076 46004 48132 46510
rect 48076 45938 48132 45948
rect 48076 41076 48132 41086
rect 48076 40982 48132 41020
rect 47852 38612 48020 38668
rect 48188 38946 48244 38958
rect 48188 38894 48190 38946
rect 48242 38894 48244 38946
rect 48188 38724 48244 38894
rect 48188 38658 48244 38668
rect 47852 37154 47908 38612
rect 47852 37102 47854 37154
rect 47906 37102 47908 37154
rect 47852 37044 47908 37102
rect 47852 36978 47908 36988
rect 48188 36258 48244 36270
rect 48188 36206 48190 36258
rect 48242 36206 48244 36258
rect 48188 36148 48244 36206
rect 48188 36082 48244 36092
rect 47740 34468 47796 34478
rect 47740 34354 47796 34412
rect 47740 34302 47742 34354
rect 47794 34302 47796 34354
rect 47740 34290 47796 34302
rect 47628 33730 47684 33740
rect 48188 34242 48244 34254
rect 48188 34190 48190 34242
rect 48242 34190 48244 34242
rect 48188 33684 48244 34190
rect 48188 33618 48244 33628
rect 48300 33796 48356 33806
rect 48188 32676 48244 32686
rect 48300 32676 48356 33740
rect 48188 32674 48356 32676
rect 48188 32622 48190 32674
rect 48242 32622 48356 32674
rect 48188 32620 48356 32622
rect 48188 32610 48244 32620
rect 47292 32510 47294 32562
rect 47346 32510 47348 32562
rect 47292 32498 47348 32510
rect 47068 32452 47124 32462
rect 46844 32450 47124 32452
rect 46844 32398 47070 32450
rect 47122 32398 47124 32450
rect 46844 32396 47124 32398
rect 46284 31892 46340 31902
rect 46172 31836 46284 31892
rect 46284 31826 46340 31836
rect 45948 29538 46004 29550
rect 45948 29486 45950 29538
rect 46002 29486 46004 29538
rect 45948 28868 46004 29486
rect 45948 28802 46004 28812
rect 47068 28866 47124 32396
rect 47516 31892 47572 31902
rect 47180 29652 47236 29662
rect 47180 29426 47236 29596
rect 47516 29650 47572 31836
rect 48188 31554 48244 31566
rect 48188 31502 48190 31554
rect 48242 31502 48244 31554
rect 48188 31220 48244 31502
rect 48188 31154 48244 31164
rect 47516 29598 47518 29650
rect 47570 29598 47572 29650
rect 47516 29586 47572 29598
rect 47180 29374 47182 29426
rect 47234 29374 47236 29426
rect 47180 29362 47236 29374
rect 47068 28814 47070 28866
rect 47122 28814 47124 28866
rect 47068 28802 47124 28814
rect 46620 28756 46676 28766
rect 46508 28084 46564 28094
rect 46620 28084 46676 28700
rect 46508 28082 46676 28084
rect 46508 28030 46510 28082
rect 46562 28030 46676 28082
rect 46508 28028 46676 28030
rect 46732 28642 46788 28654
rect 46732 28590 46734 28642
rect 46786 28590 46788 28642
rect 46508 28018 46564 28028
rect 46620 27860 46676 27870
rect 46732 27860 46788 28590
rect 48188 28532 48244 28542
rect 48188 28438 48244 28476
rect 46620 27858 46788 27860
rect 46620 27806 46622 27858
rect 46674 27806 46788 27858
rect 46620 27804 46788 27806
rect 46508 27634 46564 27646
rect 46508 27582 46510 27634
rect 46562 27582 46564 27634
rect 45948 26850 46004 26862
rect 45948 26798 45950 26850
rect 46002 26798 46004 26850
rect 45948 26068 46004 26798
rect 46284 26290 46340 26302
rect 46284 26238 46286 26290
rect 46338 26238 46340 26290
rect 45948 26012 46228 26068
rect 45836 25788 46004 25844
rect 45612 25676 45892 25732
rect 45836 25618 45892 25676
rect 45836 25566 45838 25618
rect 45890 25566 45892 25618
rect 45836 25554 45892 25566
rect 45948 25060 46004 25788
rect 46172 25396 46228 26012
rect 46284 25620 46340 26238
rect 46508 26180 46564 27582
rect 46620 26516 46676 27804
rect 48188 26850 48244 26862
rect 48188 26798 48190 26850
rect 48242 26798 48244 26850
rect 46620 26450 46676 26460
rect 47404 26516 47460 26526
rect 47404 26402 47460 26460
rect 47404 26350 47406 26402
rect 47458 26350 47460 26402
rect 47404 26338 47460 26350
rect 46732 26292 46788 26302
rect 46508 26124 46676 26180
rect 46284 25554 46340 25564
rect 46396 25508 46452 25518
rect 46396 25414 46452 25452
rect 46620 25508 46676 26124
rect 46620 25442 46676 25452
rect 46284 25396 46340 25406
rect 46172 25394 46340 25396
rect 46172 25342 46286 25394
rect 46338 25342 46340 25394
rect 46172 25340 46340 25342
rect 46284 25330 46340 25340
rect 46508 25396 46564 25406
rect 46060 25284 46116 25294
rect 46060 25282 46228 25284
rect 46060 25230 46062 25282
rect 46114 25230 46228 25282
rect 46060 25228 46228 25230
rect 46060 25218 46116 25228
rect 45948 25004 46116 25060
rect 45388 23548 45556 23604
rect 45388 23044 45444 23548
rect 45276 22148 45332 22158
rect 45276 21810 45332 22092
rect 45276 21758 45278 21810
rect 45330 21758 45332 21810
rect 45276 21746 45332 21758
rect 45388 21924 45444 22988
rect 45500 23380 45556 23390
rect 45500 22482 45556 23324
rect 45836 23380 45892 23390
rect 45836 23286 45892 23324
rect 45724 23156 45780 23166
rect 45724 23154 46004 23156
rect 45724 23102 45726 23154
rect 45778 23102 46004 23154
rect 45724 23100 46004 23102
rect 45724 23090 45780 23100
rect 45500 22430 45502 22482
rect 45554 22430 45556 22482
rect 45500 22418 45556 22430
rect 45836 22930 45892 22942
rect 45836 22878 45838 22930
rect 45890 22878 45892 22930
rect 45388 21812 45444 21868
rect 45500 21812 45556 21822
rect 45388 21810 45556 21812
rect 45388 21758 45502 21810
rect 45554 21758 45556 21810
rect 45388 21756 45556 21758
rect 45500 21746 45556 21756
rect 45836 21586 45892 22878
rect 45836 21534 45838 21586
rect 45890 21534 45892 21586
rect 45836 21522 45892 21534
rect 45948 22482 46004 23100
rect 45948 22430 45950 22482
rect 46002 22430 46004 22482
rect 45948 22260 46004 22430
rect 45388 21474 45444 21486
rect 45388 21422 45390 21474
rect 45442 21422 45444 21474
rect 45388 20802 45444 21422
rect 45388 20750 45390 20802
rect 45442 20750 45444 20802
rect 45388 20242 45444 20750
rect 45388 20190 45390 20242
rect 45442 20190 45444 20242
rect 45388 20178 45444 20190
rect 45612 20914 45668 20926
rect 45612 20862 45614 20914
rect 45666 20862 45668 20914
rect 45164 20130 45220 20142
rect 45164 20078 45166 20130
rect 45218 20078 45220 20130
rect 45052 20020 45108 20030
rect 45164 20020 45220 20078
rect 45500 20132 45556 20142
rect 45612 20132 45668 20862
rect 45500 20130 45892 20132
rect 45500 20078 45502 20130
rect 45554 20078 45892 20130
rect 45500 20076 45892 20078
rect 45500 20066 45556 20076
rect 45052 20018 45220 20020
rect 45052 19966 45054 20018
rect 45106 19966 45220 20018
rect 45052 19964 45220 19966
rect 45052 19954 45108 19964
rect 44940 19404 45108 19460
rect 44604 19170 44660 19180
rect 44940 19234 44996 19246
rect 44940 19182 44942 19234
rect 44994 19182 44996 19234
rect 44940 18340 44996 19182
rect 44380 18284 44996 18340
rect 44044 14532 44100 14542
rect 44044 14438 44100 14476
rect 44268 14532 44324 14542
rect 44268 14438 44324 14476
rect 43932 13794 43988 13804
rect 44044 13746 44100 13758
rect 44044 13694 44046 13746
rect 44098 13694 44100 13746
rect 44044 13636 44100 13694
rect 43596 13580 44100 13636
rect 43820 12180 43876 12190
rect 44044 12180 44100 13580
rect 43820 12178 44100 12180
rect 43820 12126 43822 12178
rect 43874 12126 44100 12178
rect 43820 12124 44100 12126
rect 43820 12114 43876 12124
rect 43372 11954 43540 11956
rect 43372 11902 43374 11954
rect 43426 11902 43540 11954
rect 43372 11900 43540 11902
rect 43372 11890 43428 11900
rect 43484 10724 43540 11900
rect 43260 10612 43316 10622
rect 43148 10556 43260 10612
rect 43260 10518 43316 10556
rect 43484 10610 43540 10668
rect 44380 10724 44436 10734
rect 44044 10612 44100 10650
rect 43484 10558 43486 10610
rect 43538 10558 43540 10610
rect 43484 10546 43540 10558
rect 43932 10556 44044 10612
rect 43148 10388 43204 10398
rect 42588 10386 43204 10388
rect 42588 10334 43150 10386
rect 43202 10334 43204 10386
rect 42588 10332 43204 10334
rect 42364 9884 42532 9940
rect 42140 9734 42196 9772
rect 42028 9548 42196 9604
rect 40908 9510 40964 9548
rect 41692 8372 41748 8382
rect 41692 8370 41972 8372
rect 41692 8318 41694 8370
rect 41746 8318 41972 8370
rect 41692 8316 41972 8318
rect 41692 8306 41748 8316
rect 41132 8148 41188 8158
rect 41132 8054 41188 8092
rect 41916 7700 41972 8316
rect 42028 7700 42084 7710
rect 41916 7698 42084 7700
rect 41916 7646 42030 7698
rect 42082 7646 42084 7698
rect 41916 7644 42084 7646
rect 42028 7634 42084 7644
rect 42140 7700 42196 9548
rect 42140 7698 42308 7700
rect 42140 7646 42142 7698
rect 42194 7646 42308 7698
rect 42140 7644 42308 7646
rect 42140 7634 42196 7644
rect 41468 7476 41524 7486
rect 41356 7474 41524 7476
rect 41356 7422 41470 7474
rect 41522 7422 41524 7474
rect 41356 7420 41524 7422
rect 41132 6690 41188 6702
rect 41132 6638 41134 6690
rect 41186 6638 41188 6690
rect 40908 6020 40964 6030
rect 40908 5234 40964 5964
rect 40908 5182 40910 5234
rect 40962 5182 40964 5234
rect 40908 5170 40964 5182
rect 41132 5012 41188 6638
rect 41356 6130 41412 7420
rect 41468 7410 41524 7420
rect 41916 7476 41972 7486
rect 41916 7382 41972 7420
rect 41468 7252 41524 7262
rect 41468 6578 41524 7196
rect 42252 6690 42308 7644
rect 42252 6638 42254 6690
rect 42306 6638 42308 6690
rect 42252 6626 42308 6638
rect 42476 7476 42532 9884
rect 42588 9044 42644 10332
rect 43148 10322 43204 10332
rect 43596 10386 43652 10398
rect 43596 10334 43598 10386
rect 43650 10334 43652 10386
rect 42812 10164 42868 10174
rect 42812 9826 42868 10108
rect 42812 9774 42814 9826
rect 42866 9774 42868 9826
rect 42812 9762 42868 9774
rect 42924 9828 42980 9838
rect 42924 9266 42980 9772
rect 42924 9214 42926 9266
rect 42978 9214 42980 9266
rect 42924 9202 42980 9214
rect 43484 9828 43540 9838
rect 43596 9828 43652 10334
rect 43484 9826 43652 9828
rect 43484 9774 43486 9826
rect 43538 9774 43652 9826
rect 43484 9772 43652 9774
rect 42700 9044 42756 9054
rect 42588 9042 42756 9044
rect 42588 8990 42702 9042
rect 42754 8990 42756 9042
rect 42588 8988 42756 8990
rect 42700 8978 42756 8988
rect 43372 9044 43428 9054
rect 43372 8950 43428 8988
rect 43484 9042 43540 9772
rect 43932 9266 43988 10556
rect 44044 10546 44100 10556
rect 44044 10386 44100 10398
rect 44044 10334 44046 10386
rect 44098 10334 44100 10386
rect 44044 10164 44100 10334
rect 44380 10164 44436 10668
rect 44044 10098 44100 10108
rect 44156 10108 44436 10164
rect 43932 9214 43934 9266
rect 43986 9214 43988 9266
rect 43932 9202 43988 9214
rect 44156 9266 44212 10108
rect 44268 9940 44324 9950
rect 44492 9940 44548 18284
rect 45052 18004 45108 19404
rect 45836 19346 45892 20076
rect 45836 19294 45838 19346
rect 45890 19294 45892 19346
rect 45836 19282 45892 19294
rect 45388 19236 45444 19246
rect 45388 18900 45444 19180
rect 45388 18844 45668 18900
rect 44268 9938 44548 9940
rect 44268 9886 44270 9938
rect 44322 9886 44548 9938
rect 44268 9884 44548 9886
rect 44604 17948 45108 18004
rect 44268 9874 44324 9884
rect 44156 9214 44158 9266
rect 44210 9214 44212 9266
rect 44156 9202 44212 9214
rect 43484 8990 43486 9042
rect 43538 8990 43540 9042
rect 42476 6692 42532 7420
rect 42812 8930 42868 8942
rect 42812 8878 42814 8930
rect 42866 8878 42868 8930
rect 42812 7252 42868 8878
rect 42812 7186 42868 7196
rect 42588 6692 42644 6702
rect 42476 6690 42644 6692
rect 42476 6638 42590 6690
rect 42642 6638 42644 6690
rect 42476 6636 42644 6638
rect 42588 6626 42644 6636
rect 41468 6526 41470 6578
rect 41522 6526 41524 6578
rect 41468 6514 41524 6526
rect 42140 6578 42196 6590
rect 42140 6526 42142 6578
rect 42194 6526 42196 6578
rect 41356 6078 41358 6130
rect 41410 6078 41412 6130
rect 41356 6066 41412 6078
rect 41580 6020 41636 6030
rect 41580 5926 41636 5964
rect 41692 5908 41748 5918
rect 42140 5908 42196 6526
rect 41692 5906 42196 5908
rect 41692 5854 41694 5906
rect 41746 5854 42142 5906
rect 42194 5854 42196 5906
rect 41692 5852 42196 5854
rect 41692 5842 41748 5852
rect 42140 5842 42196 5852
rect 42364 6020 42420 6030
rect 42364 5906 42420 5964
rect 43036 6020 43092 6030
rect 43484 6020 43540 8990
rect 44044 9044 44100 9054
rect 44044 8950 44100 8988
rect 43036 6018 43540 6020
rect 43036 5966 43038 6018
rect 43090 5966 43540 6018
rect 43036 5964 43540 5966
rect 43036 5954 43092 5964
rect 42364 5854 42366 5906
rect 42418 5854 42420 5906
rect 42364 5842 42420 5854
rect 41132 4946 41188 4956
rect 44604 4788 44660 17948
rect 44828 16940 45108 16996
rect 44828 16212 44884 16940
rect 45052 16882 45108 16940
rect 45052 16830 45054 16882
rect 45106 16830 45108 16882
rect 45052 16818 45108 16830
rect 44828 16098 44884 16156
rect 44828 16046 44830 16098
rect 44882 16046 44884 16098
rect 44828 16034 44884 16046
rect 44940 16770 44996 16782
rect 44940 16718 44942 16770
rect 44994 16718 44996 16770
rect 44940 16100 44996 16718
rect 45612 16210 45668 18844
rect 45724 16996 45780 17006
rect 45948 16996 46004 22204
rect 45724 16994 46004 16996
rect 45724 16942 45726 16994
rect 45778 16942 46004 16994
rect 45724 16940 46004 16942
rect 45724 16930 45780 16940
rect 45612 16158 45614 16210
rect 45666 16158 45668 16210
rect 45612 16146 45668 16158
rect 44940 16044 45220 16100
rect 45164 15986 45220 16044
rect 45164 15934 45166 15986
rect 45218 15934 45220 15986
rect 45052 15874 45108 15886
rect 45052 15822 45054 15874
rect 45106 15822 45108 15874
rect 45052 15764 45108 15822
rect 45052 15698 45108 15708
rect 45164 15148 45220 15934
rect 45500 15986 45556 15998
rect 45500 15934 45502 15986
rect 45554 15934 45556 15986
rect 45500 15764 45556 15934
rect 45724 15876 45780 15886
rect 45724 15782 45780 15820
rect 45500 15698 45556 15708
rect 45164 15092 45332 15148
rect 44828 14644 44884 14654
rect 44828 14550 44884 14588
rect 45052 14530 45108 14542
rect 45052 14478 45054 14530
rect 45106 14478 45108 14530
rect 45052 13746 45108 14478
rect 45276 13972 45332 15092
rect 45388 14532 45444 14542
rect 45388 14438 45444 14476
rect 45388 13972 45444 13982
rect 45276 13970 45444 13972
rect 45276 13918 45390 13970
rect 45442 13918 45444 13970
rect 45276 13916 45444 13918
rect 45388 13906 45444 13916
rect 45052 13694 45054 13746
rect 45106 13694 45108 13746
rect 45052 13076 45108 13694
rect 45052 13010 45108 13020
rect 44604 4722 44660 4732
rect 45276 4116 45332 4126
rect 40684 3602 40740 3612
rect 44044 3668 44100 3678
rect 44044 3574 44100 3612
rect 45276 3668 45332 4060
rect 45276 3666 45668 3668
rect 45276 3614 45278 3666
rect 45330 3614 45668 3666
rect 45276 3612 45668 3614
rect 45276 3602 45332 3612
rect 26908 3556 26964 3566
rect 26908 3462 26964 3500
rect 27356 3554 27412 3566
rect 31388 3556 31444 3566
rect 27356 3502 27358 3554
rect 27410 3502 27412 3554
rect 21532 3444 21588 3454
rect 23436 3444 23492 3454
rect 23884 3444 23940 3454
rect 21420 3388 21532 3444
rect 18844 800 18900 3388
rect 19068 3378 19124 3388
rect 19404 3378 19460 3388
rect 21532 3378 21588 3388
rect 23324 3442 23940 3444
rect 23324 3390 23438 3442
rect 23490 3390 23886 3442
rect 23938 3390 23940 3442
rect 23324 3388 23940 3390
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 23324 2212 23380 3388
rect 23436 3378 23492 3388
rect 23884 3378 23940 3388
rect 27356 3444 27412 3502
rect 30940 3554 31444 3556
rect 30940 3502 31390 3554
rect 31442 3502 31444 3554
rect 30940 3500 31444 3502
rect 28476 3444 28532 3454
rect 27356 3442 28532 3444
rect 27356 3390 28478 3442
rect 28530 3390 28532 3442
rect 27356 3388 28532 3390
rect 27356 2212 27412 3388
rect 28476 3378 28532 3388
rect 30940 3442 30996 3500
rect 31388 3490 31444 3500
rect 45612 3554 45668 3612
rect 45612 3502 45614 3554
rect 45666 3502 45668 3554
rect 45612 3490 45668 3502
rect 46060 3556 46116 25004
rect 46172 23380 46228 25228
rect 46172 22372 46228 23324
rect 46172 22278 46228 22316
rect 46396 21924 46452 21934
rect 46396 21810 46452 21868
rect 46396 21758 46398 21810
rect 46450 21758 46452 21810
rect 46396 21746 46452 21758
rect 46508 5236 46564 25340
rect 46732 24388 46788 26236
rect 48188 26292 48244 26798
rect 48188 26226 48244 26236
rect 46620 24332 46788 24388
rect 46620 22484 46676 24332
rect 46732 24164 46788 24174
rect 46732 24052 46788 24108
rect 46732 24050 47012 24052
rect 46732 23998 46734 24050
rect 46786 23998 47012 24050
rect 46732 23996 47012 23998
rect 46732 23986 46788 23996
rect 46956 23938 47012 23996
rect 46956 23886 46958 23938
rect 47010 23886 47012 23938
rect 46956 23874 47012 23886
rect 48076 23828 48132 23838
rect 48076 23734 48132 23772
rect 46620 22428 46788 22484
rect 46732 21028 46788 22428
rect 47068 22372 47124 22382
rect 46844 22260 46900 22270
rect 46844 22166 46900 22204
rect 47068 22258 47124 22316
rect 47068 22206 47070 22258
rect 47122 22206 47124 22258
rect 47068 22194 47124 22206
rect 46956 22148 47012 22158
rect 46956 22054 47012 22092
rect 46620 20972 46788 21028
rect 46956 21586 47012 21598
rect 46956 21534 46958 21586
rect 47010 21534 47012 21586
rect 46620 16660 46676 20972
rect 46732 20804 46788 20814
rect 46956 20804 47012 21534
rect 48076 21474 48132 21486
rect 48076 21422 48078 21474
rect 48130 21422 48132 21474
rect 48076 21364 48132 21422
rect 48076 21298 48132 21308
rect 46788 20748 47012 20804
rect 46732 20710 46788 20748
rect 47404 20132 47460 20142
rect 47292 20130 47460 20132
rect 47292 20078 47406 20130
rect 47458 20078 47460 20130
rect 47292 20076 47460 20078
rect 47180 19908 47236 19918
rect 47068 19852 47180 19908
rect 47068 18900 47124 19852
rect 47180 19814 47236 19852
rect 47180 19236 47236 19246
rect 47292 19236 47348 20076
rect 47404 20066 47460 20076
rect 47628 20018 47684 20030
rect 47628 19966 47630 20018
rect 47682 19966 47684 20018
rect 47628 19908 47684 19966
rect 47628 19842 47684 19852
rect 47180 19234 47348 19236
rect 47180 19182 47182 19234
rect 47234 19182 47348 19234
rect 47180 19180 47348 19182
rect 47180 19170 47236 19180
rect 48076 19124 48132 19134
rect 48076 19030 48132 19068
rect 47068 18834 47124 18844
rect 47068 16884 47124 16894
rect 47068 16882 47460 16884
rect 47068 16830 47070 16882
rect 47122 16830 47460 16882
rect 47068 16828 47460 16830
rect 47068 16818 47124 16828
rect 46620 16604 47124 16660
rect 47068 16212 47124 16604
rect 47068 16118 47124 16156
rect 47404 15986 47460 16828
rect 47740 16882 47796 16894
rect 47740 16830 47742 16882
rect 47794 16830 47796 16882
rect 47740 16436 47796 16830
rect 47740 16370 47796 16380
rect 47628 16212 47684 16222
rect 47628 16098 47684 16156
rect 47628 16046 47630 16098
rect 47682 16046 47684 16098
rect 47628 16034 47684 16046
rect 47404 15934 47406 15986
rect 47458 15934 47460 15986
rect 47404 15922 47460 15934
rect 46732 14756 46788 14766
rect 46732 14644 46788 14700
rect 46732 14642 47012 14644
rect 46732 14590 46734 14642
rect 46786 14590 47012 14642
rect 46732 14588 47012 14590
rect 46732 14578 46788 14588
rect 46956 14530 47012 14588
rect 46956 14478 46958 14530
rect 47010 14478 47012 14530
rect 46956 14466 47012 14478
rect 48076 14418 48132 14430
rect 48076 14366 48078 14418
rect 48130 14366 48132 14418
rect 48076 13972 48132 14366
rect 48076 13906 48132 13916
rect 46620 13860 46676 13870
rect 46620 6692 46676 13804
rect 46732 12180 46788 12190
rect 46956 12180 47012 12190
rect 46788 12178 47012 12180
rect 46788 12126 46958 12178
rect 47010 12126 47012 12178
rect 46788 12124 47012 12126
rect 46732 12086 46788 12124
rect 46956 12114 47012 12124
rect 47740 11954 47796 11966
rect 47740 11902 47742 11954
rect 47794 11902 47796 11954
rect 47740 11508 47796 11902
rect 47740 11442 47796 11452
rect 46732 9940 46788 9950
rect 46788 9884 47012 9940
rect 46732 9846 46788 9884
rect 46956 9826 47012 9884
rect 46956 9774 46958 9826
rect 47010 9774 47012 9826
rect 46956 9762 47012 9774
rect 48076 9714 48132 9726
rect 48076 9662 48078 9714
rect 48130 9662 48132 9714
rect 48076 9044 48132 9662
rect 48076 8978 48132 8988
rect 46732 6692 46788 6702
rect 46956 6692 47012 6702
rect 46620 6690 47012 6692
rect 46620 6638 46734 6690
rect 46786 6638 46958 6690
rect 47010 6638 47012 6690
rect 46620 6636 47012 6638
rect 46732 6626 46788 6636
rect 46956 6626 47012 6636
rect 48076 6580 48132 6590
rect 48076 6486 48132 6524
rect 46620 5236 46676 5246
rect 46508 5234 47012 5236
rect 46508 5182 46622 5234
rect 46674 5182 47012 5234
rect 46508 5180 47012 5182
rect 46620 5170 46676 5180
rect 46956 5122 47012 5180
rect 46956 5070 46958 5122
rect 47010 5070 47012 5122
rect 46956 5058 47012 5070
rect 47740 5122 47796 5134
rect 47740 5070 47742 5122
rect 47794 5070 47796 5122
rect 46620 4452 46676 4462
rect 46676 4396 47012 4452
rect 46620 4358 46676 4396
rect 46956 4338 47012 4396
rect 46956 4286 46958 4338
rect 47010 4286 47012 4338
rect 46956 4274 47012 4286
rect 46060 3490 46116 3500
rect 30940 3390 30942 3442
rect 30994 3390 30996 3442
rect 22876 2156 23380 2212
rect 26908 2156 27412 2212
rect 22876 800 22932 2156
rect 26908 800 26964 2156
rect 30940 800 30996 3390
rect 39340 3444 39396 3482
rect 39788 3444 39844 3454
rect 39340 3442 39844 3444
rect 39340 3390 39342 3442
rect 39394 3390 39790 3442
rect 39842 3390 39844 3442
rect 39340 3388 39844 3390
rect 43148 3444 43204 3454
rect 43596 3444 43652 3454
rect 43148 3442 43652 3444
rect 43148 3390 43150 3442
rect 43202 3390 43598 3442
rect 43650 3390 43652 3442
rect 43148 3388 43652 3390
rect 31164 3332 31220 3342
rect 31164 3238 31220 3276
rect 39340 2212 39396 3388
rect 39788 3378 39844 3388
rect 39004 2156 39396 2212
rect 43036 3332 43204 3388
rect 43596 3378 43652 3388
rect 46396 3442 46452 3454
rect 46396 3390 46398 3442
rect 46450 3390 46452 3442
rect 46396 3388 46452 3390
rect 46396 3332 47124 3388
rect 39004 800 39060 2156
rect 43036 800 43092 3332
rect 47068 800 47124 3332
rect 47740 1652 47796 5070
rect 48076 4226 48132 4238
rect 48076 4174 48078 4226
rect 48130 4174 48132 4226
rect 48076 4116 48132 4174
rect 48076 4050 48132 4060
rect 47740 1586 47796 1596
rect 2688 0 2800 800
rect 6720 0 6832 800
rect 10752 0 10864 800
rect 14784 0 14896 800
rect 18816 0 18928 800
rect 22848 0 22960 800
rect 26880 0 26992 800
rect 30912 0 31024 800
rect 34944 0 35056 800
rect 38976 0 39088 800
rect 43008 0 43120 800
rect 47040 0 47152 800
<< via2 >>
rect 2604 77980 2660 78036
rect 1932 76412 1988 76468
rect 1708 75570 1764 75572
rect 1708 75518 1710 75570
rect 1710 75518 1762 75570
rect 1762 75518 1764 75570
rect 1708 75516 1764 75518
rect 2604 75740 2660 75796
rect 3164 75682 3220 75684
rect 3164 75630 3166 75682
rect 3166 75630 3218 75682
rect 3218 75630 3220 75682
rect 3164 75628 3220 75630
rect 1708 73052 1764 73108
rect 1260 72380 1316 72436
rect 1148 48076 1204 48132
rect 3724 76466 3780 76468
rect 3724 76414 3726 76466
rect 3726 76414 3778 76466
rect 3778 76414 3780 76466
rect 3724 76412 3780 76414
rect 13244 76636 13300 76692
rect 13916 76636 13972 76692
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 3612 75794 3668 75796
rect 3612 75742 3614 75794
rect 3614 75742 3666 75794
rect 3666 75742 3668 75794
rect 3612 75740 3668 75742
rect 5180 75628 5236 75684
rect 4172 74844 4228 74900
rect 3948 73948 4004 74004
rect 2156 71484 2212 71540
rect 1708 70588 1764 70644
rect 1820 68124 1876 68180
rect 1596 66220 1652 66276
rect 1484 62412 1540 62468
rect 1372 56924 1428 56980
rect 1820 65714 1876 65716
rect 1820 65662 1822 65714
rect 1822 65662 1874 65714
rect 1874 65662 1876 65714
rect 1820 65660 1876 65662
rect 2268 66274 2324 66276
rect 2268 66222 2270 66274
rect 2270 66222 2322 66274
rect 2322 66222 2324 66274
rect 2268 66220 2324 66222
rect 2156 65548 2212 65604
rect 1820 63250 1876 63252
rect 1820 63198 1822 63250
rect 1822 63198 1874 63250
rect 1874 63198 1876 63250
rect 1820 63196 1876 63198
rect 2268 62636 2324 62692
rect 1596 60396 1652 60452
rect 1708 60786 1764 60788
rect 1708 60734 1710 60786
rect 1710 60734 1762 60786
rect 1762 60734 1764 60786
rect 1708 60732 1764 60734
rect 1708 58322 1764 58324
rect 1708 58270 1710 58322
rect 1710 58270 1762 58322
rect 1762 58270 1764 58322
rect 1708 58268 1764 58270
rect 2044 57036 2100 57092
rect 1708 55804 1764 55860
rect 1932 54348 1988 54404
rect 1820 53730 1876 53732
rect 1820 53678 1822 53730
rect 1822 53678 1874 53730
rect 1874 53678 1876 53730
rect 1820 53676 1876 53678
rect 1708 52946 1764 52948
rect 1708 52894 1710 52946
rect 1710 52894 1762 52946
rect 1762 52894 1764 52946
rect 1708 52892 1764 52894
rect 2492 58322 2548 58324
rect 2492 58270 2494 58322
rect 2494 58270 2546 58322
rect 2546 58270 2548 58322
rect 2492 58268 2548 58270
rect 2940 61458 2996 61460
rect 2940 61406 2942 61458
rect 2942 61406 2994 61458
rect 2994 61406 2996 61458
rect 2940 61404 2996 61406
rect 2828 57036 2884 57092
rect 2492 55804 2548 55860
rect 2492 54402 2548 54404
rect 2492 54350 2494 54402
rect 2494 54350 2546 54402
rect 2546 54350 2548 54402
rect 2492 54348 2548 54350
rect 2268 52780 2324 52836
rect 1932 50204 1988 50260
rect 2044 50092 2100 50148
rect 1932 49698 1988 49700
rect 1932 49646 1934 49698
rect 1934 49646 1986 49698
rect 1986 49646 1988 49698
rect 1932 49644 1988 49646
rect 1484 46844 1540 46900
rect 1596 48748 1652 48804
rect 1708 48412 1764 48468
rect 1932 45330 1988 45332
rect 1932 45278 1934 45330
rect 1934 45278 1986 45330
rect 1986 45278 1988 45330
rect 1932 45276 1988 45278
rect 2716 51436 2772 51492
rect 2492 50594 2548 50596
rect 2492 50542 2494 50594
rect 2494 50542 2546 50594
rect 2546 50542 2548 50594
rect 2492 50540 2548 50542
rect 2380 50204 2436 50260
rect 2492 50092 2548 50148
rect 2380 49810 2436 49812
rect 2380 49758 2382 49810
rect 2382 49758 2434 49810
rect 2434 49758 2436 49810
rect 2380 49756 2436 49758
rect 2828 50482 2884 50484
rect 2828 50430 2830 50482
rect 2830 50430 2882 50482
rect 2882 50430 2884 50482
rect 2828 50428 2884 50430
rect 2492 48242 2548 48244
rect 2492 48190 2494 48242
rect 2494 48190 2546 48242
rect 2546 48190 2548 48242
rect 2492 48188 2548 48190
rect 2492 47458 2548 47460
rect 2492 47406 2494 47458
rect 2494 47406 2546 47458
rect 2546 47406 2548 47458
rect 2492 47404 2548 47406
rect 2940 49644 2996 49700
rect 2828 47404 2884 47460
rect 2380 45276 2436 45332
rect 2828 45276 2884 45332
rect 2268 45164 2324 45220
rect 2492 45106 2548 45108
rect 2492 45054 2494 45106
rect 2494 45054 2546 45106
rect 2546 45054 2548 45106
rect 2492 45052 2548 45054
rect 1820 39228 1876 39284
rect 1596 38668 1652 38724
rect 1708 38556 1764 38612
rect 2268 43596 2324 43652
rect 2380 43538 2436 43540
rect 2380 43486 2382 43538
rect 2382 43486 2434 43538
rect 2434 43486 2436 43538
rect 2380 43484 2436 43486
rect 2156 41074 2212 41076
rect 2156 41022 2158 41074
rect 2158 41022 2210 41074
rect 2210 41022 2212 41074
rect 2156 41020 2212 41022
rect 2604 44044 2660 44100
rect 2940 43260 2996 43316
rect 2716 41356 2772 41412
rect 2492 40962 2548 40964
rect 2492 40910 2494 40962
rect 2494 40910 2546 40962
rect 2546 40910 2548 40962
rect 2492 40908 2548 40910
rect 2604 39228 2660 39284
rect 2156 38722 2212 38724
rect 2156 38670 2158 38722
rect 2158 38670 2210 38722
rect 2210 38670 2212 38722
rect 2156 38668 2212 38670
rect 2044 37436 2100 37492
rect 1372 36652 1428 36708
rect 1596 36428 1652 36484
rect 1708 36092 1764 36148
rect 1708 33628 1764 33684
rect 2268 36594 2324 36596
rect 2268 36542 2270 36594
rect 2270 36542 2322 36594
rect 2322 36542 2324 36594
rect 2268 36540 2324 36542
rect 2268 35532 2324 35588
rect 2940 38108 2996 38164
rect 3164 50540 3220 50596
rect 3388 71372 3444 71428
rect 3388 60396 3444 60452
rect 4844 74898 4900 74900
rect 4844 74846 4846 74898
rect 4846 74846 4898 74898
rect 4898 74846 4900 74898
rect 4844 74844 4900 74846
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4732 74002 4788 74004
rect 4732 73950 4734 74002
rect 4734 73950 4786 74002
rect 4786 73950 4788 74002
rect 4732 73948 4788 73950
rect 5404 75010 5460 75012
rect 5404 74958 5406 75010
rect 5406 74958 5458 75010
rect 5458 74958 5460 75010
rect 5404 74956 5460 74958
rect 6636 75010 6692 75012
rect 6636 74958 6638 75010
rect 6638 74958 6690 75010
rect 6690 74958 6692 75010
rect 6636 74956 6692 74958
rect 5740 74844 5796 74900
rect 5740 74002 5796 74004
rect 5740 73950 5742 74002
rect 5742 73950 5794 74002
rect 5794 73950 5796 74002
rect 5740 73948 5796 73950
rect 4844 73218 4900 73220
rect 4844 73166 4846 73218
rect 4846 73166 4898 73218
rect 4898 73166 4900 73218
rect 4844 73164 4900 73166
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4956 71484 5012 71540
rect 4284 71372 4340 71428
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 4284 71036 4340 71092
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4172 65548 4228 65604
rect 4060 61404 4116 61460
rect 3276 50204 3332 50260
rect 3388 54348 3444 54404
rect 4396 65490 4452 65492
rect 4396 65438 4398 65490
rect 4398 65438 4450 65490
rect 4450 65438 4452 65490
rect 4396 65436 4452 65438
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4620 62636 4676 62692
rect 5068 65996 5124 66052
rect 5628 73164 5684 73220
rect 9100 74956 9156 75012
rect 9100 74732 9156 74788
rect 9660 74786 9716 74788
rect 9660 74734 9662 74786
rect 9662 74734 9714 74786
rect 9714 74734 9716 74786
rect 9660 74732 9716 74734
rect 9100 74114 9156 74116
rect 9100 74062 9102 74114
rect 9102 74062 9154 74114
rect 9154 74062 9156 74114
rect 9100 74060 9156 74062
rect 7532 73724 7588 73780
rect 8316 73388 8372 73444
rect 9548 73442 9604 73444
rect 9548 73390 9550 73442
rect 9550 73390 9602 73442
rect 9602 73390 9604 73442
rect 9548 73388 9604 73390
rect 5852 72380 5908 72436
rect 6524 72434 6580 72436
rect 6524 72382 6526 72434
rect 6526 72382 6578 72434
rect 6578 72382 6580 72434
rect 6524 72380 6580 72382
rect 6300 71090 6356 71092
rect 6300 71038 6302 71090
rect 6302 71038 6354 71090
rect 6354 71038 6356 71090
rect 6300 71036 6356 71038
rect 5628 66050 5684 66052
rect 5628 65998 5630 66050
rect 5630 65998 5682 66050
rect 5682 65998 5684 66050
rect 5628 65996 5684 65998
rect 5404 65772 5460 65828
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 5852 68626 5908 68628
rect 5852 68574 5854 68626
rect 5854 68574 5906 68626
rect 5906 68574 5908 68626
rect 5852 68572 5908 68574
rect 6188 70476 6244 70532
rect 6524 70364 6580 70420
rect 6636 69298 6692 69300
rect 6636 69246 6638 69298
rect 6638 69246 6690 69298
rect 6690 69246 6692 69298
rect 6636 69244 6692 69246
rect 8428 71148 8484 71204
rect 9212 71148 9268 71204
rect 8204 70700 8260 70756
rect 7084 70588 7140 70644
rect 7644 70418 7700 70420
rect 7644 70366 7646 70418
rect 7646 70366 7698 70418
rect 7698 70366 7700 70418
rect 7644 70364 7700 70366
rect 8428 70364 8484 70420
rect 8204 70252 8260 70308
rect 6972 69244 7028 69300
rect 7084 69186 7140 69188
rect 7084 69134 7086 69186
rect 7086 69134 7138 69186
rect 7138 69134 7140 69186
rect 7084 69132 7140 69134
rect 6412 68908 6468 68964
rect 6636 68572 6692 68628
rect 6524 67564 6580 67620
rect 7644 67954 7700 67956
rect 7644 67902 7646 67954
rect 7646 67902 7698 67954
rect 7698 67902 7700 67954
rect 7644 67900 7700 67902
rect 7532 67730 7588 67732
rect 7532 67678 7534 67730
rect 7534 67678 7586 67730
rect 7586 67678 7588 67730
rect 7532 67676 7588 67678
rect 7756 67618 7812 67620
rect 7756 67566 7758 67618
rect 7758 67566 7810 67618
rect 7810 67566 7812 67618
rect 7756 67564 7812 67566
rect 6636 67228 6692 67284
rect 7756 67228 7812 67284
rect 6748 66220 6804 66276
rect 6188 65212 6244 65268
rect 6524 64428 6580 64484
rect 6748 64652 6804 64708
rect 6636 63250 6692 63252
rect 6636 63198 6638 63250
rect 6638 63198 6690 63250
rect 6690 63198 6692 63250
rect 6636 63196 6692 63198
rect 6300 62914 6356 62916
rect 6300 62862 6302 62914
rect 6302 62862 6354 62914
rect 6354 62862 6356 62914
rect 6300 62860 6356 62862
rect 5740 62412 5796 62468
rect 6412 62300 6468 62356
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4956 58828 5012 58884
rect 5180 61516 5236 61572
rect 4684 58772 4740 58774
rect 5852 61516 5908 61572
rect 5516 61404 5572 61460
rect 5740 61292 5796 61348
rect 5516 60786 5572 60788
rect 5516 60734 5518 60786
rect 5518 60734 5570 60786
rect 5570 60734 5572 60786
rect 5516 60732 5572 60734
rect 5180 58380 5236 58436
rect 5852 61180 5908 61236
rect 6300 61570 6356 61572
rect 6300 61518 6302 61570
rect 6302 61518 6354 61570
rect 6354 61518 6356 61570
rect 6300 61516 6356 61518
rect 4620 58156 4676 58212
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4844 54572 4900 54628
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4172 53116 4228 53172
rect 3612 52050 3668 52052
rect 3612 51998 3614 52050
rect 3614 51998 3666 52050
rect 3666 51998 3668 52050
rect 3612 51996 3668 51998
rect 3836 51884 3892 51940
rect 3724 50706 3780 50708
rect 3724 50654 3726 50706
rect 3726 50654 3778 50706
rect 3778 50654 3780 50706
rect 3724 50652 3780 50654
rect 3836 50428 3892 50484
rect 3612 48354 3668 48356
rect 3612 48302 3614 48354
rect 3614 48302 3666 48354
rect 3666 48302 3668 48354
rect 3612 48300 3668 48302
rect 3388 47516 3444 47572
rect 3500 48188 3556 48244
rect 3612 47628 3668 47684
rect 3164 45218 3220 45220
rect 3164 45166 3166 45218
rect 3166 45166 3218 45218
rect 3218 45166 3220 45218
rect 3164 45164 3220 45166
rect 3388 45164 3444 45220
rect 3388 44156 3444 44212
rect 3612 44994 3668 44996
rect 3612 44942 3614 44994
rect 3614 44942 3666 44994
rect 3666 44942 3668 44994
rect 3612 44940 3668 44942
rect 3612 43932 3668 43988
rect 3164 41916 3220 41972
rect 3164 40908 3220 40964
rect 3164 39676 3220 39732
rect 2268 34130 2324 34132
rect 2268 34078 2270 34130
rect 2270 34078 2322 34130
rect 2322 34078 2324 34130
rect 2268 34076 2324 34078
rect 2044 33628 2100 33684
rect 2716 34018 2772 34020
rect 2716 33966 2718 34018
rect 2718 33966 2770 34018
rect 2770 33966 2772 34018
rect 2716 33964 2772 33966
rect 2156 33852 2212 33908
rect 1932 33068 1988 33124
rect 2044 32284 2100 32340
rect 1932 31666 1988 31668
rect 1932 31614 1934 31666
rect 1934 31614 1986 31666
rect 1986 31614 1988 31666
rect 1932 31612 1988 31614
rect 1932 31164 1988 31220
rect 1708 29932 1764 29988
rect 1932 30268 1988 30324
rect 1820 29260 1876 29316
rect 1820 28700 1876 28756
rect 1708 28642 1764 28644
rect 1708 28590 1710 28642
rect 1710 28590 1762 28642
rect 1762 28590 1764 28642
rect 1708 28588 1764 28590
rect 2380 33516 2436 33572
rect 2940 33906 2996 33908
rect 2940 33854 2942 33906
rect 2942 33854 2994 33906
rect 2994 33854 2996 33906
rect 2940 33852 2996 33854
rect 2492 32732 2548 32788
rect 2828 32732 2884 32788
rect 2716 32060 2772 32116
rect 2940 32562 2996 32564
rect 2940 32510 2942 32562
rect 2942 32510 2994 32562
rect 2994 32510 2996 32562
rect 2940 32508 2996 32510
rect 2492 31612 2548 31668
rect 2268 29986 2324 29988
rect 2268 29934 2270 29986
rect 2270 29934 2322 29986
rect 2322 29934 2324 29986
rect 2268 29932 2324 29934
rect 2940 30828 2996 30884
rect 2604 28588 2660 28644
rect 3836 47570 3892 47572
rect 3836 47518 3838 47570
rect 3838 47518 3890 47570
rect 3890 47518 3892 47570
rect 3836 47516 3892 47518
rect 3836 46674 3892 46676
rect 3836 46622 3838 46674
rect 3838 46622 3890 46674
rect 3890 46622 3892 46674
rect 3836 46620 3892 46622
rect 3836 45276 3892 45332
rect 4172 52162 4228 52164
rect 4172 52110 4174 52162
rect 4174 52110 4226 52162
rect 4226 52110 4228 52162
rect 4172 52108 4228 52110
rect 4172 51490 4228 51492
rect 4172 51438 4174 51490
rect 4174 51438 4226 51490
rect 4226 51438 4228 51490
rect 4172 51436 4228 51438
rect 4060 50428 4116 50484
rect 5068 53506 5124 53508
rect 5068 53454 5070 53506
rect 5070 53454 5122 53506
rect 5122 53454 5124 53506
rect 5068 53452 5124 53454
rect 5180 54460 5236 54516
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4732 52332 4788 52388
rect 4844 52220 4900 52276
rect 4956 52050 5012 52052
rect 4956 51998 4958 52050
rect 4958 51998 5010 52050
rect 5010 51998 5012 52050
rect 4956 51996 5012 51998
rect 4844 51324 4900 51380
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4508 50594 4564 50596
rect 4508 50542 4510 50594
rect 4510 50542 4562 50594
rect 4562 50542 4564 50594
rect 4508 50540 4564 50542
rect 4060 49756 4116 49812
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4396 48412 4452 48468
rect 4844 48466 4900 48468
rect 4844 48414 4846 48466
rect 4846 48414 4898 48466
rect 4898 48414 4900 48466
rect 4844 48412 4900 48414
rect 4284 48242 4340 48244
rect 4284 48190 4286 48242
rect 4286 48190 4338 48242
rect 4338 48190 4340 48242
rect 4284 48188 4340 48190
rect 4172 47404 4228 47460
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4732 47628 4788 47684
rect 4844 47458 4900 47460
rect 4844 47406 4846 47458
rect 4846 47406 4898 47458
rect 4898 47406 4900 47458
rect 4844 47404 4900 47406
rect 4396 47346 4452 47348
rect 4396 47294 4398 47346
rect 4398 47294 4450 47346
rect 4450 47294 4452 47346
rect 4396 47292 4452 47294
rect 4956 47346 5012 47348
rect 4956 47294 4958 47346
rect 4958 47294 5010 47346
rect 5010 47294 5012 47346
rect 4956 47292 5012 47294
rect 4172 46620 4228 46676
rect 4844 47068 4900 47124
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 3948 44380 4004 44436
rect 3724 44268 3780 44324
rect 4172 44268 4228 44324
rect 3948 44210 4004 44212
rect 3948 44158 3950 44210
rect 3950 44158 4002 44210
rect 4002 44158 4004 44210
rect 3948 44156 4004 44158
rect 4060 44098 4116 44100
rect 4060 44046 4062 44098
rect 4062 44046 4114 44098
rect 4114 44046 4116 44098
rect 4060 44044 4116 44046
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4732 44098 4788 44100
rect 4732 44046 4734 44098
rect 4734 44046 4786 44098
rect 4786 44046 4788 44098
rect 4732 44044 4788 44046
rect 3612 43596 3668 43652
rect 3388 39452 3444 39508
rect 3500 41020 3556 41076
rect 3388 38892 3444 38948
rect 3388 34018 3444 34020
rect 3388 33966 3390 34018
rect 3390 33966 3442 34018
rect 3442 33966 3444 34018
rect 3388 33964 3444 33966
rect 3388 33516 3444 33572
rect 3388 32732 3444 32788
rect 2268 27858 2324 27860
rect 2268 27806 2270 27858
rect 2270 27806 2322 27858
rect 2322 27806 2324 27858
rect 2268 27804 2324 27806
rect 2604 27020 2660 27076
rect 1708 26236 1764 26292
rect 3276 30268 3332 30324
rect 3724 42754 3780 42756
rect 3724 42702 3726 42754
rect 3726 42702 3778 42754
rect 3778 42702 3780 42754
rect 3724 42700 3780 42702
rect 3724 41074 3780 41076
rect 3724 41022 3726 41074
rect 3726 41022 3778 41074
rect 3778 41022 3780 41074
rect 3724 41020 3780 41022
rect 3948 39058 4004 39060
rect 3948 39006 3950 39058
rect 3950 39006 4002 39058
rect 4002 39006 4004 39058
rect 3948 39004 4004 39006
rect 3612 38444 3668 38500
rect 3948 37772 4004 37828
rect 3724 34972 3780 35028
rect 3836 36370 3892 36372
rect 3836 36318 3838 36370
rect 3838 36318 3890 36370
rect 3890 36318 3892 36370
rect 3836 36316 3892 36318
rect 3612 34300 3668 34356
rect 3836 33964 3892 34020
rect 3836 32508 3892 32564
rect 3836 31948 3892 32004
rect 3836 31612 3892 31668
rect 2940 27858 2996 27860
rect 2940 27806 2942 27858
rect 2942 27806 2994 27858
rect 2994 27806 2996 27858
rect 2940 27804 2996 27806
rect 3276 27074 3332 27076
rect 3276 27022 3278 27074
rect 3278 27022 3330 27074
rect 3330 27022 3332 27074
rect 3276 27020 3332 27022
rect 3612 27804 3668 27860
rect 2940 26962 2996 26964
rect 2940 26910 2942 26962
rect 2942 26910 2994 26962
rect 2994 26910 2996 26962
rect 2940 26908 2996 26910
rect 1596 23996 1652 24052
rect 2268 24050 2324 24052
rect 2268 23998 2270 24050
rect 2270 23998 2322 24050
rect 2322 23998 2324 24050
rect 2268 23996 2324 23998
rect 1708 23826 1764 23828
rect 1708 23774 1710 23826
rect 1710 23774 1762 23826
rect 1762 23774 1764 23826
rect 1708 23772 1764 23774
rect 1260 21644 1316 21700
rect 2268 21756 2324 21812
rect 1708 21308 1764 21364
rect 1148 20188 1204 20244
rect 3612 23548 3668 23604
rect 4060 35026 4116 35028
rect 4060 34974 4062 35026
rect 4062 34974 4114 35026
rect 4114 34974 4116 35026
rect 4060 34972 4116 34974
rect 5180 45164 5236 45220
rect 4956 44044 5012 44100
rect 4732 43596 4788 43652
rect 4620 43538 4676 43540
rect 4620 43486 4622 43538
rect 4622 43486 4674 43538
rect 4674 43486 4676 43538
rect 4620 43484 4676 43486
rect 4732 43372 4788 43428
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5068 43148 5124 43204
rect 4956 42700 5012 42756
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5740 58210 5796 58212
rect 5740 58158 5742 58210
rect 5742 58158 5794 58210
rect 5794 58158 5796 58210
rect 5740 58156 5796 58158
rect 6188 59052 6244 59108
rect 6636 60732 6692 60788
rect 6972 63196 7028 63252
rect 6860 61346 6916 61348
rect 6860 61294 6862 61346
rect 6862 61294 6914 61346
rect 6914 61294 6916 61346
rect 6860 61292 6916 61294
rect 6972 61180 7028 61236
rect 6412 59052 6468 59108
rect 5964 58492 6020 58548
rect 6300 58546 6356 58548
rect 6300 58494 6302 58546
rect 6302 58494 6354 58546
rect 6354 58494 6356 58546
rect 6300 58492 6356 58494
rect 5964 57708 6020 57764
rect 5740 56924 5796 56980
rect 6860 59106 6916 59108
rect 6860 59054 6862 59106
rect 6862 59054 6914 59106
rect 6914 59054 6916 59106
rect 6860 59052 6916 59054
rect 6524 58940 6580 58996
rect 6748 58492 6804 58548
rect 6636 58434 6692 58436
rect 6636 58382 6638 58434
rect 6638 58382 6690 58434
rect 6690 58382 6692 58434
rect 6636 58380 6692 58382
rect 6524 57708 6580 57764
rect 6076 57372 6132 57428
rect 5740 56140 5796 56196
rect 5516 53452 5572 53508
rect 5628 52162 5684 52164
rect 5628 52110 5630 52162
rect 5630 52110 5682 52162
rect 5682 52110 5684 52162
rect 5628 52108 5684 52110
rect 5628 51378 5684 51380
rect 5628 51326 5630 51378
rect 5630 51326 5682 51378
rect 5682 51326 5684 51378
rect 5628 51324 5684 51326
rect 5628 50652 5684 50708
rect 5852 54514 5908 54516
rect 5852 54462 5854 54514
rect 5854 54462 5906 54514
rect 5906 54462 5908 54514
rect 5852 54460 5908 54462
rect 6076 54684 6132 54740
rect 6188 54626 6244 54628
rect 6188 54574 6190 54626
rect 6190 54574 6242 54626
rect 6242 54574 6244 54626
rect 6188 54572 6244 54574
rect 6076 53900 6132 53956
rect 5852 52444 5908 52500
rect 5964 53564 6020 53620
rect 5964 52332 6020 52388
rect 7308 65772 7364 65828
rect 7196 65548 7252 65604
rect 7196 64652 7252 64708
rect 7196 64482 7252 64484
rect 7196 64430 7198 64482
rect 7198 64430 7250 64482
rect 7250 64430 7252 64482
rect 7196 64428 7252 64430
rect 7196 63084 7252 63140
rect 7084 60396 7140 60452
rect 7196 62860 7252 62916
rect 7644 65602 7700 65604
rect 7644 65550 7646 65602
rect 7646 65550 7698 65602
rect 7698 65550 7700 65602
rect 7644 65548 7700 65550
rect 7756 65324 7812 65380
rect 7644 65266 7700 65268
rect 7644 65214 7646 65266
rect 7646 65214 7698 65266
rect 7698 65214 7700 65266
rect 7644 65212 7700 65214
rect 7756 63196 7812 63252
rect 7644 63084 7700 63140
rect 7308 61740 7364 61796
rect 7196 61292 7252 61348
rect 7420 59388 7476 59444
rect 7196 57820 7252 57876
rect 7084 57484 7140 57540
rect 7084 56812 7140 56868
rect 6524 54460 6580 54516
rect 7420 58434 7476 58436
rect 7420 58382 7422 58434
rect 7422 58382 7474 58434
rect 7474 58382 7476 58434
rect 7420 58380 7476 58382
rect 7420 58044 7476 58100
rect 6636 53564 6692 53620
rect 7756 62354 7812 62356
rect 7756 62302 7758 62354
rect 7758 62302 7810 62354
rect 7810 62302 7812 62354
rect 7756 62300 7812 62302
rect 8428 69970 8484 69972
rect 8428 69918 8430 69970
rect 8430 69918 8482 69970
rect 8482 69918 8484 69970
rect 8428 69916 8484 69918
rect 8092 68572 8148 68628
rect 10668 74732 10724 74788
rect 10892 73948 10948 74004
rect 13580 76412 13636 76468
rect 15148 76466 15204 76468
rect 15148 76414 15150 76466
rect 15150 76414 15202 76466
rect 15202 76414 15204 76466
rect 15148 76412 15204 76414
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 14700 75628 14756 75684
rect 15932 75628 15988 75684
rect 12460 74002 12516 74004
rect 12460 73950 12462 74002
rect 12462 73950 12514 74002
rect 12514 73950 12516 74002
rect 12460 73948 12516 73950
rect 15596 74284 15652 74340
rect 14028 73948 14084 74004
rect 11788 73388 11844 73444
rect 11116 71260 11172 71316
rect 12796 72380 12852 72436
rect 9884 70588 9940 70644
rect 9996 70364 10052 70420
rect 8204 67676 8260 67732
rect 7980 67564 8036 67620
rect 8316 65490 8372 65492
rect 8316 65438 8318 65490
rect 8318 65438 8370 65490
rect 8370 65438 8372 65490
rect 8316 65436 8372 65438
rect 8540 68908 8596 68964
rect 8764 69244 8820 69300
rect 8764 68908 8820 68964
rect 10444 70418 10500 70420
rect 10444 70366 10446 70418
rect 10446 70366 10498 70418
rect 10498 70366 10500 70418
rect 10444 70364 10500 70366
rect 10220 70194 10276 70196
rect 10220 70142 10222 70194
rect 10222 70142 10274 70194
rect 10274 70142 10276 70194
rect 10220 70140 10276 70142
rect 9996 68908 10052 68964
rect 9548 68626 9604 68628
rect 9548 68574 9550 68626
rect 9550 68574 9602 68626
rect 9602 68574 9604 68626
rect 9548 68572 9604 68574
rect 9436 66274 9492 66276
rect 9436 66222 9438 66274
rect 9438 66222 9490 66274
rect 9490 66222 9492 66274
rect 9436 66220 9492 66222
rect 10668 67340 10724 67396
rect 10108 66220 10164 66276
rect 8652 65378 8708 65380
rect 8652 65326 8654 65378
rect 8654 65326 8706 65378
rect 8706 65326 8708 65378
rect 8652 65324 8708 65326
rect 9548 64706 9604 64708
rect 9548 64654 9550 64706
rect 9550 64654 9602 64706
rect 9602 64654 9604 64706
rect 9548 64652 9604 64654
rect 8764 64594 8820 64596
rect 8764 64542 8766 64594
rect 8766 64542 8818 64594
rect 8818 64542 8820 64594
rect 8764 64540 8820 64542
rect 7644 57874 7700 57876
rect 7644 57822 7646 57874
rect 7646 57822 7698 57874
rect 7698 57822 7700 57874
rect 7644 57820 7700 57822
rect 8204 62300 8260 62356
rect 7644 56866 7700 56868
rect 7644 56814 7646 56866
rect 7646 56814 7698 56866
rect 7698 56814 7700 56866
rect 7644 56812 7700 56814
rect 7868 61740 7924 61796
rect 8092 60396 8148 60452
rect 7980 59164 8036 59220
rect 7868 58940 7924 58996
rect 8428 61740 8484 61796
rect 8652 62300 8708 62356
rect 8316 58322 8372 58324
rect 8316 58270 8318 58322
rect 8318 58270 8370 58322
rect 8370 58270 8372 58322
rect 8316 58268 8372 58270
rect 7868 58044 7924 58100
rect 8428 57932 8484 57988
rect 8092 57820 8148 57876
rect 8652 59388 8708 59444
rect 8652 58828 8708 58884
rect 8988 64146 9044 64148
rect 8988 64094 8990 64146
rect 8990 64094 9042 64146
rect 9042 64094 9044 64146
rect 8988 64092 9044 64094
rect 10892 65378 10948 65380
rect 10892 65326 10894 65378
rect 10894 65326 10946 65378
rect 10946 65326 10948 65378
rect 10892 65324 10948 65326
rect 10892 64988 10948 65044
rect 10780 64764 10836 64820
rect 10108 64652 10164 64708
rect 10668 64652 10724 64708
rect 9884 64092 9940 64148
rect 10220 64594 10276 64596
rect 10220 64542 10222 64594
rect 10222 64542 10274 64594
rect 10274 64542 10276 64594
rect 10220 64540 10276 64542
rect 10332 64316 10388 64372
rect 10556 64204 10612 64260
rect 8988 62242 9044 62244
rect 8988 62190 8990 62242
rect 8990 62190 9042 62242
rect 9042 62190 9044 62242
rect 8988 62188 9044 62190
rect 10444 62524 10500 62580
rect 10780 64034 10836 64036
rect 10780 63982 10782 64034
rect 10782 63982 10834 64034
rect 10834 63982 10836 64034
rect 10780 63980 10836 63982
rect 11788 70812 11844 70868
rect 11452 70588 11508 70644
rect 11116 64204 11172 64260
rect 11228 64316 11284 64372
rect 12908 72268 12964 72324
rect 11788 70252 11844 70308
rect 12460 70364 12516 70420
rect 12012 69468 12068 69524
rect 11676 67340 11732 67396
rect 12796 69522 12852 69524
rect 12796 69470 12798 69522
rect 12798 69470 12850 69522
rect 12850 69470 12852 69522
rect 12796 69468 12852 69470
rect 13692 70364 13748 70420
rect 14140 70140 14196 70196
rect 12236 66162 12292 66164
rect 12236 66110 12238 66162
rect 12238 66110 12290 66162
rect 12290 66110 12292 66162
rect 12236 66108 12292 66110
rect 11564 64876 11620 64932
rect 11788 65490 11844 65492
rect 11788 65438 11790 65490
rect 11790 65438 11842 65490
rect 11842 65438 11844 65490
rect 11788 65436 11844 65438
rect 11564 64594 11620 64596
rect 11564 64542 11566 64594
rect 11566 64542 11618 64594
rect 11618 64542 11620 64594
rect 11564 64540 11620 64542
rect 12572 65490 12628 65492
rect 12572 65438 12574 65490
rect 12574 65438 12626 65490
rect 12626 65438 12628 65490
rect 12572 65436 12628 65438
rect 12348 65212 12404 65268
rect 12012 64876 12068 64932
rect 11452 64204 11508 64260
rect 11788 64034 11844 64036
rect 11788 63982 11790 64034
rect 11790 63982 11842 64034
rect 11842 63982 11844 64034
rect 11788 63980 11844 63982
rect 10780 63756 10836 63812
rect 10108 62188 10164 62244
rect 9660 60786 9716 60788
rect 9660 60734 9662 60786
rect 9662 60734 9714 60786
rect 9714 60734 9716 60786
rect 9660 60732 9716 60734
rect 10108 60396 10164 60452
rect 10668 60396 10724 60452
rect 9548 59218 9604 59220
rect 9548 59166 9550 59218
rect 9550 59166 9602 59218
rect 9602 59166 9604 59218
rect 9548 59164 9604 59166
rect 8764 58604 8820 58660
rect 9436 58604 9492 58660
rect 8764 57762 8820 57764
rect 8764 57710 8766 57762
rect 8766 57710 8818 57762
rect 8818 57710 8820 57762
rect 8764 57708 8820 57710
rect 8092 56812 8148 56868
rect 8764 57538 8820 57540
rect 8764 57486 8766 57538
rect 8766 57486 8818 57538
rect 8818 57486 8820 57538
rect 8764 57484 8820 57486
rect 8540 57426 8596 57428
rect 8540 57374 8542 57426
rect 8542 57374 8594 57426
rect 8594 57374 8596 57426
rect 8540 57372 8596 57374
rect 8988 57148 9044 57204
rect 7868 55804 7924 55860
rect 6300 52668 6356 52724
rect 6188 52332 6244 52388
rect 6748 52668 6804 52724
rect 6300 51996 6356 52052
rect 6748 52050 6804 52052
rect 6748 51998 6750 52050
rect 6750 51998 6802 52050
rect 6802 51998 6804 52050
rect 6748 51996 6804 51998
rect 6524 51324 6580 51380
rect 6188 50988 6244 51044
rect 5516 49420 5572 49476
rect 5404 47068 5460 47124
rect 5404 46786 5460 46788
rect 5404 46734 5406 46786
rect 5406 46734 5458 46786
rect 5458 46734 5460 46786
rect 5404 46732 5460 46734
rect 5852 49532 5908 49588
rect 5740 46786 5796 46788
rect 5740 46734 5742 46786
rect 5742 46734 5794 46786
rect 5794 46734 5796 46786
rect 5740 46732 5796 46734
rect 5852 46284 5908 46340
rect 5740 45890 5796 45892
rect 5740 45838 5742 45890
rect 5742 45838 5794 45890
rect 5794 45838 5796 45890
rect 5740 45836 5796 45838
rect 5516 44044 5572 44100
rect 5404 42812 5460 42868
rect 5180 42476 5236 42532
rect 5404 42476 5460 42532
rect 5740 43036 5796 43092
rect 5852 43484 5908 43540
rect 5628 42754 5684 42756
rect 5628 42702 5630 42754
rect 5630 42702 5682 42754
rect 5682 42702 5684 42754
rect 5628 42700 5684 42702
rect 5068 41020 5124 41076
rect 4732 40626 4788 40628
rect 4732 40574 4734 40626
rect 4734 40574 4786 40626
rect 4786 40574 4788 40626
rect 4732 40572 4788 40574
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4284 39452 4340 39508
rect 4620 39004 4676 39060
rect 4844 38892 4900 38948
rect 4284 38556 4340 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4396 37266 4452 37268
rect 4396 37214 4398 37266
rect 4398 37214 4450 37266
rect 4450 37214 4452 37266
rect 4396 37212 4452 37214
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4396 36652 4452 36708
rect 5516 41580 5572 41636
rect 5516 40626 5572 40628
rect 5516 40574 5518 40626
rect 5518 40574 5570 40626
rect 5570 40574 5572 40626
rect 5516 40572 5572 40574
rect 5740 42530 5796 42532
rect 5740 42478 5742 42530
rect 5742 42478 5794 42530
rect 5794 42478 5796 42530
rect 5740 42476 5796 42478
rect 6860 50652 6916 50708
rect 6076 48466 6132 48468
rect 6076 48414 6078 48466
rect 6078 48414 6130 48466
rect 6130 48414 6132 48466
rect 6076 48412 6132 48414
rect 6636 49420 6692 49476
rect 6636 48412 6692 48468
rect 6748 46844 6804 46900
rect 6860 45276 6916 45332
rect 6300 44434 6356 44436
rect 6300 44382 6302 44434
rect 6302 44382 6354 44434
rect 6354 44382 6356 44434
rect 6300 44380 6356 44382
rect 6524 44044 6580 44100
rect 6636 43820 6692 43876
rect 6188 43036 6244 43092
rect 6636 43484 6692 43540
rect 6636 42700 6692 42756
rect 7532 53170 7588 53172
rect 7532 53118 7534 53170
rect 7534 53118 7586 53170
rect 7586 53118 7588 53170
rect 7532 53116 7588 53118
rect 7644 51324 7700 51380
rect 7644 50482 7700 50484
rect 7644 50430 7646 50482
rect 7646 50430 7698 50482
rect 7698 50430 7700 50482
rect 7644 50428 7700 50430
rect 7756 50988 7812 51044
rect 7196 48188 7252 48244
rect 7084 45276 7140 45332
rect 8204 55804 8260 55860
rect 8092 54514 8148 54516
rect 8092 54462 8094 54514
rect 8094 54462 8146 54514
rect 8146 54462 8148 54514
rect 8092 54460 8148 54462
rect 8092 52444 8148 52500
rect 8540 54738 8596 54740
rect 8540 54686 8542 54738
rect 8542 54686 8594 54738
rect 8594 54686 8596 54738
rect 8540 54684 8596 54686
rect 8428 54348 8484 54404
rect 8428 52668 8484 52724
rect 8316 51996 8372 52052
rect 8988 56866 9044 56868
rect 8988 56814 8990 56866
rect 8990 56814 9042 56866
rect 9042 56814 9044 56866
rect 8988 56812 9044 56814
rect 9548 58044 9604 58100
rect 9996 59106 10052 59108
rect 9996 59054 9998 59106
rect 9998 59054 10050 59106
rect 10050 59054 10052 59106
rect 9996 59052 10052 59054
rect 10668 58940 10724 58996
rect 9996 58210 10052 58212
rect 9996 58158 9998 58210
rect 9998 58158 10050 58210
rect 10050 58158 10052 58210
rect 9996 58156 10052 58158
rect 10668 58716 10724 58772
rect 10556 58210 10612 58212
rect 10556 58158 10558 58210
rect 10558 58158 10610 58210
rect 10610 58158 10612 58210
rect 10556 58156 10612 58158
rect 9884 57762 9940 57764
rect 9884 57710 9886 57762
rect 9886 57710 9938 57762
rect 9938 57710 9940 57762
rect 9884 57708 9940 57710
rect 9884 56866 9940 56868
rect 9884 56814 9886 56866
rect 9886 56814 9938 56866
rect 9938 56814 9940 56866
rect 9884 56812 9940 56814
rect 10108 57932 10164 57988
rect 10668 57820 10724 57876
rect 10108 57484 10164 57540
rect 11116 62578 11172 62580
rect 11116 62526 11118 62578
rect 11118 62526 11170 62578
rect 11170 62526 11172 62578
rect 11116 62524 11172 62526
rect 13020 65772 13076 65828
rect 12796 65212 12852 65268
rect 12572 64594 12628 64596
rect 12572 64542 12574 64594
rect 12574 64542 12626 64594
rect 12626 64542 12628 64594
rect 12572 64540 12628 64542
rect 12236 64092 12292 64148
rect 11900 63644 11956 63700
rect 11452 62524 11508 62580
rect 11228 61570 11284 61572
rect 11228 61518 11230 61570
rect 11230 61518 11282 61570
rect 11282 61518 11284 61570
rect 11228 61516 11284 61518
rect 11228 60396 11284 60452
rect 11004 58044 11060 58100
rect 10780 57596 10836 57652
rect 10444 57484 10500 57540
rect 10332 56812 10388 56868
rect 9660 55804 9716 55860
rect 9660 55580 9716 55636
rect 8876 53170 8932 53172
rect 8876 53118 8878 53170
rect 8878 53118 8930 53170
rect 8930 53118 8932 53170
rect 8876 53116 8932 53118
rect 8876 52556 8932 52612
rect 9548 52780 9604 52836
rect 8764 52444 8820 52500
rect 8652 51884 8708 51940
rect 8540 51548 8596 51604
rect 8316 50540 8372 50596
rect 8428 50428 8484 50484
rect 8204 48972 8260 49028
rect 7644 47234 7700 47236
rect 7644 47182 7646 47234
rect 7646 47182 7698 47234
rect 7698 47182 7700 47234
rect 7644 47180 7700 47182
rect 7532 46898 7588 46900
rect 7532 46846 7534 46898
rect 7534 46846 7586 46898
rect 7586 46846 7588 46898
rect 7532 46844 7588 46846
rect 7420 44940 7476 44996
rect 7084 44098 7140 44100
rect 7084 44046 7086 44098
rect 7086 44046 7138 44098
rect 7138 44046 7140 44098
rect 7084 44044 7140 44046
rect 7644 44380 7700 44436
rect 7084 43372 7140 43428
rect 6972 43036 7028 43092
rect 7084 42978 7140 42980
rect 7084 42926 7086 42978
rect 7086 42926 7138 42978
rect 7138 42926 7140 42978
rect 7084 42924 7140 42926
rect 6972 42642 7028 42644
rect 6972 42590 6974 42642
rect 6974 42590 7026 42642
rect 7026 42590 7028 42642
rect 6972 42588 7028 42590
rect 6748 42364 6804 42420
rect 6188 41580 6244 41636
rect 7084 41580 7140 41636
rect 6076 41020 6132 41076
rect 5404 38946 5460 38948
rect 5404 38894 5406 38946
rect 5406 38894 5458 38946
rect 5458 38894 5460 38946
rect 5404 38892 5460 38894
rect 5068 36370 5124 36372
rect 5068 36318 5070 36370
rect 5070 36318 5122 36370
rect 5122 36318 5124 36370
rect 5068 36316 5124 36318
rect 5180 36258 5236 36260
rect 5180 36206 5182 36258
rect 5182 36206 5234 36258
rect 5234 36206 5236 36258
rect 5180 36204 5236 36206
rect 4956 35586 5012 35588
rect 4956 35534 4958 35586
rect 4958 35534 5010 35586
rect 5010 35534 5012 35586
rect 4956 35532 5012 35534
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4956 35308 5012 35364
rect 5628 35308 5684 35364
rect 4284 34914 4340 34916
rect 4284 34862 4286 34914
rect 4286 34862 4338 34914
rect 4338 34862 4340 34914
rect 4284 34860 4340 34862
rect 5068 35026 5124 35028
rect 5068 34974 5070 35026
rect 5070 34974 5122 35026
rect 5122 34974 5124 35026
rect 5068 34972 5124 34974
rect 6076 36258 6132 36260
rect 6076 36206 6078 36258
rect 6078 36206 6130 36258
rect 6130 36206 6132 36258
rect 6076 36204 6132 36206
rect 4396 34748 4452 34804
rect 5964 34914 6020 34916
rect 5964 34862 5966 34914
rect 5966 34862 6018 34914
rect 6018 34862 6020 34914
rect 5964 34860 6020 34862
rect 4620 34354 4676 34356
rect 4620 34302 4622 34354
rect 4622 34302 4674 34354
rect 4674 34302 4676 34354
rect 4620 34300 4676 34302
rect 5068 34300 5124 34356
rect 4284 34188 4340 34244
rect 5180 34242 5236 34244
rect 5180 34190 5182 34242
rect 5182 34190 5234 34242
rect 5234 34190 5236 34242
rect 5180 34188 5236 34190
rect 4732 33964 4788 34020
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4284 33404 4340 33460
rect 4284 32786 4340 32788
rect 4284 32734 4286 32786
rect 4286 32734 4338 32786
rect 4338 32734 4340 32786
rect 4284 32732 4340 32734
rect 4844 33180 4900 33236
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4620 31388 4676 31444
rect 4956 31388 5012 31444
rect 4844 30940 4900 30996
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4956 30882 5012 30884
rect 4956 30830 4958 30882
rect 4958 30830 5010 30882
rect 5010 30830 5012 30882
rect 4956 30828 5012 30830
rect 4060 26962 4116 26964
rect 4060 26910 4062 26962
rect 4062 26910 4114 26962
rect 4114 26910 4116 26962
rect 4060 26908 4116 26910
rect 5180 30210 5236 30212
rect 5180 30158 5182 30210
rect 5182 30158 5234 30210
rect 5234 30158 5236 30210
rect 5180 30156 5236 30158
rect 5740 34690 5796 34692
rect 5740 34638 5742 34690
rect 5742 34638 5794 34690
rect 5794 34638 5796 34690
rect 5740 34636 5796 34638
rect 5740 33234 5796 33236
rect 5740 33182 5742 33234
rect 5742 33182 5794 33234
rect 5794 33182 5796 33234
rect 5740 33180 5796 33182
rect 5740 31388 5796 31444
rect 5516 30604 5572 30660
rect 4396 29596 4452 29652
rect 5404 29650 5460 29652
rect 5404 29598 5406 29650
rect 5406 29598 5458 29650
rect 5458 29598 5460 29650
rect 5404 29596 5460 29598
rect 5740 29820 5796 29876
rect 5740 29538 5796 29540
rect 5740 29486 5742 29538
rect 5742 29486 5794 29538
rect 5794 29486 5796 29538
rect 5740 29484 5796 29486
rect 4844 29314 4900 29316
rect 4844 29262 4846 29314
rect 4846 29262 4898 29314
rect 4898 29262 4900 29314
rect 4844 29260 4900 29262
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4620 28754 4676 28756
rect 4620 28702 4622 28754
rect 4622 28702 4674 28754
rect 4674 28702 4676 28754
rect 4620 28700 4676 28702
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5740 29036 5796 29092
rect 5068 28642 5124 28644
rect 5068 28590 5070 28642
rect 5070 28590 5122 28642
rect 5122 28590 5124 28642
rect 5068 28588 5124 28590
rect 4956 26908 5012 26964
rect 6188 34524 6244 34580
rect 6188 34300 6244 34356
rect 6076 32508 6132 32564
rect 5964 32338 6020 32340
rect 5964 32286 5966 32338
rect 5966 32286 6018 32338
rect 6018 32286 6020 32338
rect 5964 32284 6020 32286
rect 6076 31500 6132 31556
rect 5964 30156 6020 30212
rect 6748 41020 6804 41076
rect 7308 42754 7364 42756
rect 7308 42702 7310 42754
rect 7310 42702 7362 42754
rect 7362 42702 7364 42754
rect 7308 42700 7364 42702
rect 7308 42364 7364 42420
rect 7196 40796 7252 40852
rect 6860 39842 6916 39844
rect 6860 39790 6862 39842
rect 6862 39790 6914 39842
rect 6914 39790 6916 39842
rect 6860 39788 6916 39790
rect 8204 48242 8260 48244
rect 8204 48190 8206 48242
rect 8206 48190 8258 48242
rect 8258 48190 8260 48242
rect 8204 48188 8260 48190
rect 8204 47404 8260 47460
rect 8652 51660 8708 51716
rect 8540 48412 8596 48468
rect 7980 45836 8036 45892
rect 7868 45106 7924 45108
rect 7868 45054 7870 45106
rect 7870 45054 7922 45106
rect 7922 45054 7924 45106
rect 7868 45052 7924 45054
rect 7644 41916 7700 41972
rect 7532 40012 7588 40068
rect 7420 39618 7476 39620
rect 7420 39566 7422 39618
rect 7422 39566 7474 39618
rect 7474 39566 7476 39618
rect 7420 39564 7476 39566
rect 6524 37100 6580 37156
rect 7084 39340 7140 39396
rect 6860 36652 6916 36708
rect 6860 36316 6916 36372
rect 6860 35196 6916 35252
rect 6748 34748 6804 34804
rect 6412 34188 6468 34244
rect 6300 33404 6356 33460
rect 6524 33852 6580 33908
rect 6972 34860 7028 34916
rect 6972 33516 7028 33572
rect 6300 32620 6356 32676
rect 6524 32450 6580 32452
rect 6524 32398 6526 32450
rect 6526 32398 6578 32450
rect 6578 32398 6580 32450
rect 6524 32396 6580 32398
rect 6748 31948 6804 32004
rect 6188 31388 6244 31444
rect 6524 31388 6580 31444
rect 6412 30994 6468 30996
rect 6412 30942 6414 30994
rect 6414 30942 6466 30994
rect 6466 30942 6468 30994
rect 6412 30940 6468 30942
rect 6076 29820 6132 29876
rect 6636 29820 6692 29876
rect 6076 29036 6132 29092
rect 5852 28700 5908 28756
rect 5852 26962 5908 26964
rect 5852 26910 5854 26962
rect 5854 26910 5906 26962
rect 5906 26910 5908 26962
rect 5852 26908 5908 26910
rect 5068 26236 5124 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4620 25506 4676 25508
rect 4620 25454 4622 25506
rect 4622 25454 4674 25506
rect 4674 25454 4676 25506
rect 4620 25452 4676 25454
rect 4284 25116 4340 25172
rect 5628 26290 5684 26292
rect 5628 26238 5630 26290
rect 5630 26238 5682 26290
rect 5682 26238 5684 26290
rect 5628 26236 5684 26238
rect 5292 25452 5348 25508
rect 4844 25004 4900 25060
rect 5180 25116 5236 25172
rect 4732 24834 4788 24836
rect 4732 24782 4734 24834
rect 4734 24782 4786 24834
rect 4786 24782 4788 24834
rect 4732 24780 4788 24782
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5068 21586 5124 21588
rect 5068 21534 5070 21586
rect 5070 21534 5122 21586
rect 5122 21534 5124 21586
rect 5068 21532 5124 21534
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4060 20748 4116 20804
rect 3948 19964 4004 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5852 25564 5908 25620
rect 5628 25506 5684 25508
rect 5628 25454 5630 25506
rect 5630 25454 5682 25506
rect 5682 25454 5684 25506
rect 5628 25452 5684 25454
rect 6860 31836 6916 31892
rect 6748 27244 6804 27300
rect 6748 25564 6804 25620
rect 5852 25228 5908 25284
rect 6076 25004 6132 25060
rect 6412 24780 6468 24836
rect 6860 25004 6916 25060
rect 5852 23324 5908 23380
rect 6412 23548 6468 23604
rect 6188 23042 6244 23044
rect 6188 22990 6190 23042
rect 6190 22990 6242 23042
rect 6242 22990 6244 23042
rect 6188 22988 6244 22990
rect 5628 21532 5684 21588
rect 5964 20802 6020 20804
rect 5964 20750 5966 20802
rect 5966 20750 6018 20802
rect 6018 20750 6020 20802
rect 5964 20748 6020 20750
rect 6860 23378 6916 23380
rect 6860 23326 6862 23378
rect 6862 23326 6914 23378
rect 6914 23326 6916 23378
rect 6860 23324 6916 23326
rect 7756 39788 7812 39844
rect 7756 39452 7812 39508
rect 7196 38946 7252 38948
rect 7196 38894 7198 38946
rect 7198 38894 7250 38946
rect 7250 38894 7252 38946
rect 7196 38892 7252 38894
rect 7308 38834 7364 38836
rect 7308 38782 7310 38834
rect 7310 38782 7362 38834
rect 7362 38782 7364 38834
rect 7308 38780 7364 38782
rect 7644 38444 7700 38500
rect 7644 37660 7700 37716
rect 7644 37212 7700 37268
rect 7532 37100 7588 37156
rect 7420 35196 7476 35252
rect 8316 46898 8372 46900
rect 8316 46846 8318 46898
rect 8318 46846 8370 46898
rect 8370 46846 8372 46898
rect 8316 46844 8372 46846
rect 8316 45164 8372 45220
rect 8540 45276 8596 45332
rect 8764 51378 8820 51380
rect 8764 51326 8766 51378
rect 8766 51326 8818 51378
rect 8818 51326 8820 51378
rect 8764 51324 8820 51326
rect 8876 50428 8932 50484
rect 8764 50204 8820 50260
rect 8764 46956 8820 47012
rect 8988 49026 9044 49028
rect 8988 48974 8990 49026
rect 8990 48974 9042 49026
rect 9042 48974 9044 49026
rect 8988 48972 9044 48974
rect 9772 53564 9828 53620
rect 10220 54348 10276 54404
rect 9884 52946 9940 52948
rect 9884 52894 9886 52946
rect 9886 52894 9938 52946
rect 9938 52894 9940 52946
rect 9884 52892 9940 52894
rect 10780 55186 10836 55188
rect 10780 55134 10782 55186
rect 10782 55134 10834 55186
rect 10834 55134 10836 55186
rect 10780 55132 10836 55134
rect 10556 53618 10612 53620
rect 10556 53566 10558 53618
rect 10558 53566 10610 53618
rect 10610 53566 10612 53618
rect 10556 53564 10612 53566
rect 10332 52946 10388 52948
rect 10332 52894 10334 52946
rect 10334 52894 10386 52946
rect 10386 52894 10388 52946
rect 10332 52892 10388 52894
rect 10780 53004 10836 53060
rect 10556 52668 10612 52724
rect 9660 51660 9716 51716
rect 9772 51602 9828 51604
rect 9772 51550 9774 51602
rect 9774 51550 9826 51602
rect 9826 51550 9828 51602
rect 9772 51548 9828 51550
rect 10332 51266 10388 51268
rect 10332 51214 10334 51266
rect 10334 51214 10386 51266
rect 10386 51214 10388 51266
rect 10332 51212 10388 51214
rect 10556 51212 10612 51268
rect 10668 52946 10724 52948
rect 10668 52894 10670 52946
rect 10670 52894 10722 52946
rect 10722 52894 10724 52946
rect 10668 52892 10724 52894
rect 9772 50594 9828 50596
rect 9772 50542 9774 50594
rect 9774 50542 9826 50594
rect 9826 50542 9828 50594
rect 9772 50540 9828 50542
rect 10220 50482 10276 50484
rect 10220 50430 10222 50482
rect 10222 50430 10274 50482
rect 10274 50430 10276 50482
rect 10220 50428 10276 50430
rect 8988 48466 9044 48468
rect 8988 48414 8990 48466
rect 8990 48414 9042 48466
rect 9042 48414 9044 48466
rect 8988 48412 9044 48414
rect 8988 48188 9044 48244
rect 9548 48466 9604 48468
rect 9548 48414 9550 48466
rect 9550 48414 9602 48466
rect 9602 48414 9604 48466
rect 9548 48412 9604 48414
rect 9884 48412 9940 48468
rect 8988 46732 9044 46788
rect 8876 45276 8932 45332
rect 8316 44604 8372 44660
rect 8428 44716 8484 44772
rect 8652 44940 8708 44996
rect 8876 45052 8932 45108
rect 8540 43426 8596 43428
rect 8540 43374 8542 43426
rect 8542 43374 8594 43426
rect 8594 43374 8596 43426
rect 8540 43372 8596 43374
rect 8652 44604 8708 44660
rect 9100 44940 9156 44996
rect 9212 47180 9268 47236
rect 8988 43596 9044 43652
rect 8876 42924 8932 42980
rect 9100 43484 9156 43540
rect 8428 41356 8484 41412
rect 8540 41916 8596 41972
rect 8092 39564 8148 39620
rect 7980 39506 8036 39508
rect 7980 39454 7982 39506
rect 7982 39454 8034 39506
rect 8034 39454 8036 39506
rect 7980 39452 8036 39454
rect 8204 39452 8260 39508
rect 8092 39340 8148 39396
rect 8092 38946 8148 38948
rect 8092 38894 8094 38946
rect 8094 38894 8146 38946
rect 8146 38894 8148 38946
rect 8092 38892 8148 38894
rect 7868 38668 7924 38724
rect 7980 38780 8036 38836
rect 7644 34972 7700 35028
rect 7532 34636 7588 34692
rect 7420 32844 7476 32900
rect 7084 31724 7140 31780
rect 7196 32396 7252 32452
rect 8428 40962 8484 40964
rect 8428 40910 8430 40962
rect 8430 40910 8482 40962
rect 8482 40910 8484 40962
rect 8428 40908 8484 40910
rect 8988 41858 9044 41860
rect 8988 41806 8990 41858
rect 8990 41806 9042 41858
rect 9042 41806 9044 41858
rect 8988 41804 9044 41806
rect 8540 40572 8596 40628
rect 8316 40236 8372 40292
rect 9324 45724 9380 45780
rect 9324 43596 9380 43652
rect 8988 39452 9044 39508
rect 8540 39340 8596 39396
rect 8316 38834 8372 38836
rect 8316 38782 8318 38834
rect 8318 38782 8370 38834
rect 8370 38782 8372 38834
rect 8316 38780 8372 38782
rect 8988 38780 9044 38836
rect 7980 36540 8036 36596
rect 8092 38332 8148 38388
rect 8204 38274 8260 38276
rect 8204 38222 8206 38274
rect 8206 38222 8258 38274
rect 8258 38222 8260 38274
rect 8204 38220 8260 38222
rect 8876 38108 8932 38164
rect 8204 37212 8260 37268
rect 8316 37100 8372 37156
rect 8764 36594 8820 36596
rect 8764 36542 8766 36594
rect 8766 36542 8818 36594
rect 8818 36542 8820 36594
rect 8764 36540 8820 36542
rect 7756 34802 7812 34804
rect 7756 34750 7758 34802
rect 7758 34750 7810 34802
rect 7810 34750 7812 34802
rect 7756 34748 7812 34750
rect 7756 32732 7812 32788
rect 7644 32396 7700 32452
rect 7196 31052 7252 31108
rect 7532 31836 7588 31892
rect 7420 31500 7476 31556
rect 7308 30940 7364 30996
rect 7532 29650 7588 29652
rect 7532 29598 7534 29650
rect 7534 29598 7586 29650
rect 7586 29598 7588 29650
rect 7532 29596 7588 29598
rect 7420 27244 7476 27300
rect 7756 31052 7812 31108
rect 7980 34300 8036 34356
rect 8092 33292 8148 33348
rect 8204 33180 8260 33236
rect 7980 32508 8036 32564
rect 8092 32732 8148 32788
rect 7868 30828 7924 30884
rect 7756 30268 7812 30324
rect 8092 31724 8148 31780
rect 8540 34300 8596 34356
rect 8428 33906 8484 33908
rect 8428 33854 8430 33906
rect 8430 33854 8482 33906
rect 8482 33854 8484 33906
rect 8428 33852 8484 33854
rect 8652 33404 8708 33460
rect 8876 35252 8932 35308
rect 8652 32844 8708 32900
rect 8092 31164 8148 31220
rect 8428 32620 8484 32676
rect 8316 30994 8372 30996
rect 8316 30942 8318 30994
rect 8318 30942 8370 30994
rect 8370 30942 8372 30994
rect 8316 30940 8372 30942
rect 8428 30268 8484 30324
rect 8540 32284 8596 32340
rect 8652 31500 8708 31556
rect 8652 30828 8708 30884
rect 8876 31500 8932 31556
rect 8876 30044 8932 30100
rect 9548 45778 9604 45780
rect 9548 45726 9550 45778
rect 9550 45726 9602 45778
rect 9602 45726 9604 45778
rect 9548 45724 9604 45726
rect 10332 50316 10388 50372
rect 9884 46898 9940 46900
rect 9884 46846 9886 46898
rect 9886 46846 9938 46898
rect 9938 46846 9940 46898
rect 9884 46844 9940 46846
rect 9996 45836 10052 45892
rect 10220 45778 10276 45780
rect 10220 45726 10222 45778
rect 10222 45726 10274 45778
rect 10274 45726 10276 45778
rect 10220 45724 10276 45726
rect 9772 45052 9828 45108
rect 9660 44994 9716 44996
rect 9660 44942 9662 44994
rect 9662 44942 9714 44994
rect 9714 44942 9716 44994
rect 9660 44940 9716 44942
rect 9436 43260 9492 43316
rect 9548 43538 9604 43540
rect 9548 43486 9550 43538
rect 9550 43486 9602 43538
rect 9602 43486 9604 43538
rect 9548 43484 9604 43486
rect 10108 43708 10164 43764
rect 11116 56642 11172 56644
rect 11116 56590 11118 56642
rect 11118 56590 11170 56642
rect 11170 56590 11172 56642
rect 11116 56588 11172 56590
rect 11788 61516 11844 61572
rect 11564 61180 11620 61236
rect 12012 61292 12068 61348
rect 12124 60508 12180 60564
rect 11564 58940 11620 58996
rect 11004 55580 11060 55636
rect 11004 53564 11060 53620
rect 11228 53058 11284 53060
rect 11228 53006 11230 53058
rect 11230 53006 11282 53058
rect 11282 53006 11284 53058
rect 11228 53004 11284 53006
rect 10780 52444 10836 52500
rect 10668 50316 10724 50372
rect 10444 50204 10500 50260
rect 11004 49922 11060 49924
rect 11004 49870 11006 49922
rect 11006 49870 11058 49922
rect 11058 49870 11060 49922
rect 11004 49868 11060 49870
rect 11116 49810 11172 49812
rect 11116 49758 11118 49810
rect 11118 49758 11170 49810
rect 11170 49758 11172 49810
rect 11116 49756 11172 49758
rect 10556 49698 10612 49700
rect 10556 49646 10558 49698
rect 10558 49646 10610 49698
rect 10610 49646 10612 49698
rect 10556 49644 10612 49646
rect 11116 49532 11172 49588
rect 11564 58268 11620 58324
rect 12572 62076 12628 62132
rect 13020 64316 13076 64372
rect 14476 67564 14532 67620
rect 15372 70588 15428 70644
rect 20076 76300 20132 76356
rect 19068 75794 19124 75796
rect 19068 75742 19070 75794
rect 19070 75742 19122 75794
rect 19122 75742 19124 75794
rect 19068 75740 19124 75742
rect 19068 75180 19124 75236
rect 16380 73948 16436 74004
rect 16828 74002 16884 74004
rect 16828 73950 16830 74002
rect 16830 73950 16882 74002
rect 16882 73950 16884 74002
rect 16828 73948 16884 73950
rect 18172 74786 18228 74788
rect 18172 74734 18174 74786
rect 18174 74734 18226 74786
rect 18226 74734 18228 74786
rect 18172 74732 18228 74734
rect 18172 74172 18228 74228
rect 17388 73948 17444 74004
rect 16604 73218 16660 73220
rect 16604 73166 16606 73218
rect 16606 73166 16658 73218
rect 16658 73166 16660 73218
rect 16604 73164 16660 73166
rect 17164 73164 17220 73220
rect 17612 73164 17668 73220
rect 17948 73276 18004 73332
rect 18620 73330 18676 73332
rect 18620 73278 18622 73330
rect 18622 73278 18674 73330
rect 18674 73278 18676 73330
rect 18620 73276 18676 73278
rect 19068 73948 19124 74004
rect 18844 72828 18900 72884
rect 18956 73276 19012 73332
rect 18172 72658 18228 72660
rect 18172 72606 18174 72658
rect 18174 72606 18226 72658
rect 18226 72606 18228 72658
rect 18172 72604 18228 72606
rect 18956 72658 19012 72660
rect 18956 72606 18958 72658
rect 18958 72606 19010 72658
rect 19010 72606 19012 72658
rect 18956 72604 19012 72606
rect 16604 71372 16660 71428
rect 16716 71260 16772 71316
rect 16268 70140 16324 70196
rect 14812 67058 14868 67060
rect 14812 67006 14814 67058
rect 14814 67006 14866 67058
rect 14866 67006 14868 67058
rect 14812 67004 14868 67006
rect 13580 65490 13636 65492
rect 13580 65438 13582 65490
rect 13582 65438 13634 65490
rect 13634 65438 13636 65490
rect 13580 65436 13636 65438
rect 13468 65324 13524 65380
rect 13916 65996 13972 66052
rect 14252 65772 14308 65828
rect 14140 65602 14196 65604
rect 14140 65550 14142 65602
rect 14142 65550 14194 65602
rect 14194 65550 14196 65602
rect 14140 65548 14196 65550
rect 14252 65436 14308 65492
rect 13244 63980 13300 64036
rect 13132 63196 13188 63252
rect 12684 61570 12740 61572
rect 12684 61518 12686 61570
rect 12686 61518 12738 61570
rect 12738 61518 12740 61570
rect 12684 61516 12740 61518
rect 12796 61068 12852 61124
rect 12908 62188 12964 62244
rect 12236 58380 12292 58436
rect 12684 59948 12740 60004
rect 11676 57708 11732 57764
rect 12348 58156 12404 58212
rect 12124 56700 12180 56756
rect 11564 56642 11620 56644
rect 11564 56590 11566 56642
rect 11566 56590 11618 56642
rect 11618 56590 11620 56642
rect 11564 56588 11620 56590
rect 11564 56194 11620 56196
rect 11564 56142 11566 56194
rect 11566 56142 11618 56194
rect 11618 56142 11620 56194
rect 11564 56140 11620 56142
rect 12124 56194 12180 56196
rect 12124 56142 12126 56194
rect 12126 56142 12178 56194
rect 12178 56142 12180 56194
rect 12124 56140 12180 56142
rect 12124 55468 12180 55524
rect 11900 55132 11956 55188
rect 12572 57596 12628 57652
rect 12348 56754 12404 56756
rect 12348 56702 12350 56754
rect 12350 56702 12402 56754
rect 12402 56702 12404 56754
rect 12348 56700 12404 56702
rect 13020 61458 13076 61460
rect 13020 61406 13022 61458
rect 13022 61406 13074 61458
rect 13074 61406 13076 61458
rect 13020 61404 13076 61406
rect 12684 56588 12740 56644
rect 11452 54012 11508 54068
rect 11900 54012 11956 54068
rect 11564 53564 11620 53620
rect 11788 51884 11844 51940
rect 11340 50204 11396 50260
rect 11564 50092 11620 50148
rect 11228 48748 11284 48804
rect 11452 49980 11508 50036
rect 10780 47964 10836 48020
rect 10556 47458 10612 47460
rect 10556 47406 10558 47458
rect 10558 47406 10610 47458
rect 10610 47406 10612 47458
rect 10556 47404 10612 47406
rect 10668 46844 10724 46900
rect 10556 46284 10612 46340
rect 10444 44380 10500 44436
rect 10892 47180 10948 47236
rect 11228 46786 11284 46788
rect 11228 46734 11230 46786
rect 11230 46734 11282 46786
rect 11282 46734 11284 46786
rect 11228 46732 11284 46734
rect 11116 46284 11172 46340
rect 12348 51938 12404 51940
rect 12348 51886 12350 51938
rect 12350 51886 12402 51938
rect 12402 51886 12404 51938
rect 12348 51884 12404 51886
rect 12236 50316 12292 50372
rect 12348 49922 12404 49924
rect 12348 49870 12350 49922
rect 12350 49870 12402 49922
rect 12402 49870 12404 49922
rect 12348 49868 12404 49870
rect 12124 49756 12180 49812
rect 12236 49586 12292 49588
rect 12236 49534 12238 49586
rect 12238 49534 12290 49586
rect 12290 49534 12292 49586
rect 12236 49532 12292 49534
rect 11564 46844 11620 46900
rect 11676 46508 11732 46564
rect 11228 45778 11284 45780
rect 11228 45726 11230 45778
rect 11230 45726 11282 45778
rect 11282 45726 11284 45778
rect 11228 45724 11284 45726
rect 11004 45500 11060 45556
rect 10892 44380 10948 44436
rect 9548 43148 9604 43204
rect 9660 43372 9716 43428
rect 9996 42364 10052 42420
rect 10220 42476 10276 42532
rect 9996 41804 10052 41860
rect 9772 40908 9828 40964
rect 9660 40626 9716 40628
rect 9660 40574 9662 40626
rect 9662 40574 9714 40626
rect 9714 40574 9716 40626
rect 9660 40572 9716 40574
rect 9436 38108 9492 38164
rect 9436 37324 9492 37380
rect 9548 37266 9604 37268
rect 9548 37214 9550 37266
rect 9550 37214 9602 37266
rect 9602 37214 9604 37266
rect 9548 37212 9604 37214
rect 10108 40290 10164 40292
rect 10108 40238 10110 40290
rect 10110 40238 10162 40290
rect 10162 40238 10164 40290
rect 10108 40236 10164 40238
rect 11004 43596 11060 43652
rect 10556 43538 10612 43540
rect 10556 43486 10558 43538
rect 10558 43486 10610 43538
rect 10610 43486 10612 43538
rect 10556 43484 10612 43486
rect 10556 42476 10612 42532
rect 10556 40012 10612 40068
rect 9548 35980 9604 36036
rect 9100 34354 9156 34356
rect 9100 34302 9102 34354
rect 9102 34302 9154 34354
rect 9154 34302 9156 34354
rect 9100 34300 9156 34302
rect 9100 31836 9156 31892
rect 8988 29148 9044 29204
rect 8204 27132 8260 27188
rect 7420 25228 7476 25284
rect 9772 34524 9828 34580
rect 9324 34300 9380 34356
rect 9548 33346 9604 33348
rect 9548 33294 9550 33346
rect 9550 33294 9602 33346
rect 9602 33294 9604 33346
rect 9548 33292 9604 33294
rect 9324 33234 9380 33236
rect 9324 33182 9326 33234
rect 9326 33182 9378 33234
rect 9378 33182 9380 33234
rect 9324 33180 9380 33182
rect 9548 33122 9604 33124
rect 9548 33070 9550 33122
rect 9550 33070 9602 33122
rect 9602 33070 9604 33122
rect 9548 33068 9604 33070
rect 9548 32674 9604 32676
rect 9548 32622 9550 32674
rect 9550 32622 9602 32674
rect 9602 32622 9604 32674
rect 9548 32620 9604 32622
rect 9660 32508 9716 32564
rect 9996 33180 10052 33236
rect 9996 31948 10052 32004
rect 12572 52162 12628 52164
rect 12572 52110 12574 52162
rect 12574 52110 12626 52162
rect 12626 52110 12628 52162
rect 12572 52108 12628 52110
rect 12908 54908 12964 54964
rect 13468 63922 13524 63924
rect 13468 63870 13470 63922
rect 13470 63870 13522 63922
rect 13522 63870 13524 63922
rect 13468 63868 13524 63870
rect 15260 67618 15316 67620
rect 15260 67566 15262 67618
rect 15262 67566 15314 67618
rect 15314 67566 15316 67618
rect 15260 67564 15316 67566
rect 15036 66274 15092 66276
rect 15036 66222 15038 66274
rect 15038 66222 15090 66274
rect 15090 66222 15092 66274
rect 15036 66220 15092 66222
rect 15932 66946 15988 66948
rect 15932 66894 15934 66946
rect 15934 66894 15986 66946
rect 15986 66894 15988 66946
rect 15932 66892 15988 66894
rect 14924 65772 14980 65828
rect 14700 65490 14756 65492
rect 14700 65438 14702 65490
rect 14702 65438 14754 65490
rect 14754 65438 14756 65490
rect 14700 65436 14756 65438
rect 13916 64540 13972 64596
rect 14588 64594 14644 64596
rect 14588 64542 14590 64594
rect 14590 64542 14642 64594
rect 14642 64542 14644 64594
rect 14588 64540 14644 64542
rect 14252 63980 14308 64036
rect 13916 63868 13972 63924
rect 14028 62524 14084 62580
rect 13692 61404 13748 61460
rect 13580 61346 13636 61348
rect 13580 61294 13582 61346
rect 13582 61294 13634 61346
rect 13634 61294 13636 61346
rect 13580 61292 13636 61294
rect 13804 61292 13860 61348
rect 13468 61180 13524 61236
rect 13356 59612 13412 59668
rect 13356 56754 13412 56756
rect 13356 56702 13358 56754
rect 13358 56702 13410 56754
rect 13410 56702 13412 56754
rect 13356 56700 13412 56702
rect 13804 58156 13860 58212
rect 13804 57708 13860 57764
rect 13468 56194 13524 56196
rect 13468 56142 13470 56194
rect 13470 56142 13522 56194
rect 13522 56142 13524 56194
rect 13468 56140 13524 56142
rect 13356 55916 13412 55972
rect 13580 55522 13636 55524
rect 13580 55470 13582 55522
rect 13582 55470 13634 55522
rect 13634 55470 13636 55522
rect 13580 55468 13636 55470
rect 14812 65266 14868 65268
rect 14812 65214 14814 65266
rect 14814 65214 14866 65266
rect 14866 65214 14868 65266
rect 14812 65212 14868 65214
rect 15036 65660 15092 65716
rect 15596 66050 15652 66052
rect 15596 65998 15598 66050
rect 15598 65998 15650 66050
rect 15650 65998 15652 66050
rect 15596 65996 15652 65998
rect 15260 65602 15316 65604
rect 15260 65550 15262 65602
rect 15262 65550 15314 65602
rect 15314 65550 15316 65602
rect 15260 65548 15316 65550
rect 15596 65436 15652 65492
rect 15596 65100 15652 65156
rect 15148 64652 15204 64708
rect 15484 64482 15540 64484
rect 15484 64430 15486 64482
rect 15486 64430 15538 64482
rect 15538 64430 15540 64482
rect 15484 64428 15540 64430
rect 14924 63532 14980 63588
rect 14700 62578 14756 62580
rect 14700 62526 14702 62578
rect 14702 62526 14754 62578
rect 14754 62526 14756 62578
rect 14700 62524 14756 62526
rect 14924 62354 14980 62356
rect 14924 62302 14926 62354
rect 14926 62302 14978 62354
rect 14978 62302 14980 62354
rect 14924 62300 14980 62302
rect 14364 61516 14420 61572
rect 14028 60844 14084 60900
rect 14140 61068 14196 61124
rect 13916 56194 13972 56196
rect 13916 56142 13918 56194
rect 13918 56142 13970 56194
rect 13970 56142 13972 56194
rect 13916 56140 13972 56142
rect 13804 56082 13860 56084
rect 13804 56030 13806 56082
rect 13806 56030 13858 56082
rect 13858 56030 13860 56082
rect 13804 56028 13860 56030
rect 13916 55916 13972 55972
rect 13580 54908 13636 54964
rect 12908 52780 12964 52836
rect 12684 50988 12740 51044
rect 13580 54626 13636 54628
rect 13580 54574 13582 54626
rect 13582 54574 13634 54626
rect 13634 54574 13636 54626
rect 13580 54572 13636 54574
rect 12684 50316 12740 50372
rect 13132 53788 13188 53844
rect 12572 48354 12628 48356
rect 12572 48302 12574 48354
rect 12574 48302 12626 48354
rect 12626 48302 12628 48354
rect 12572 48300 12628 48302
rect 12572 46060 12628 46116
rect 11900 45778 11956 45780
rect 11900 45726 11902 45778
rect 11902 45726 11954 45778
rect 11954 45726 11956 45778
rect 11900 45724 11956 45726
rect 11676 43538 11732 43540
rect 11676 43486 11678 43538
rect 11678 43486 11730 43538
rect 11730 43486 11732 43538
rect 11676 43484 11732 43486
rect 11228 42812 11284 42868
rect 10892 42476 10948 42532
rect 12012 43596 12068 43652
rect 12236 45612 12292 45668
rect 12348 45500 12404 45556
rect 13020 48412 13076 48468
rect 13020 47740 13076 47796
rect 11228 39676 11284 39732
rect 11116 39394 11172 39396
rect 11116 39342 11118 39394
rect 11118 39342 11170 39394
rect 11170 39342 11172 39394
rect 11116 39340 11172 39342
rect 10332 33516 10388 33572
rect 10332 33234 10388 33236
rect 10332 33182 10334 33234
rect 10334 33182 10386 33234
rect 10386 33182 10388 33234
rect 10332 33180 10388 33182
rect 10108 32732 10164 32788
rect 9548 31666 9604 31668
rect 9548 31614 9550 31666
rect 9550 31614 9602 31666
rect 9602 31614 9604 31666
rect 9548 31612 9604 31614
rect 9996 31554 10052 31556
rect 9996 31502 9998 31554
rect 9998 31502 10050 31554
rect 10050 31502 10052 31554
rect 9996 31500 10052 31502
rect 9660 31164 9716 31220
rect 9548 30940 9604 30996
rect 10220 33122 10276 33124
rect 10220 33070 10222 33122
rect 10222 33070 10274 33122
rect 10274 33070 10276 33122
rect 10220 33068 10276 33070
rect 10668 33122 10724 33124
rect 10668 33070 10670 33122
rect 10670 33070 10722 33122
rect 10722 33070 10724 33122
rect 10668 33068 10724 33070
rect 11004 32674 11060 32676
rect 11004 32622 11006 32674
rect 11006 32622 11058 32674
rect 11058 32622 11060 32674
rect 11004 32620 11060 32622
rect 10220 32284 10276 32340
rect 10668 32508 10724 32564
rect 10892 31948 10948 32004
rect 9884 30994 9940 30996
rect 9884 30942 9886 30994
rect 9886 30942 9938 30994
rect 9938 30942 9940 30994
rect 9884 30940 9940 30942
rect 9436 28700 9492 28756
rect 8876 27186 8932 27188
rect 8876 27134 8878 27186
rect 8878 27134 8930 27186
rect 8930 27134 8932 27186
rect 8876 27132 8932 27134
rect 10108 31052 10164 31108
rect 10556 29596 10612 29652
rect 10780 30828 10836 30884
rect 9772 29148 9828 29204
rect 10780 28588 10836 28644
rect 9884 28476 9940 28532
rect 7756 25618 7812 25620
rect 7756 25566 7758 25618
rect 7758 25566 7810 25618
rect 7810 25566 7812 25618
rect 7756 25564 7812 25566
rect 8316 25228 8372 25284
rect 7644 22988 7700 23044
rect 7644 22428 7700 22484
rect 8540 22482 8596 22484
rect 8540 22430 8542 22482
rect 8542 22430 8594 22482
rect 8594 22430 8596 22482
rect 8540 22428 8596 22430
rect 8428 22370 8484 22372
rect 8428 22318 8430 22370
rect 8430 22318 8482 22370
rect 8482 22318 8484 22370
rect 8428 22316 8484 22318
rect 6972 21756 7028 21812
rect 8316 21586 8372 21588
rect 8316 21534 8318 21586
rect 8318 21534 8370 21586
rect 8370 21534 8372 21586
rect 8316 21532 8372 21534
rect 6412 18060 6468 18116
rect 5516 17388 5572 17444
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 7308 3442 7364 3444
rect 7308 3390 7310 3442
rect 7310 3390 7362 3442
rect 7362 3390 7364 3442
rect 7308 3388 7364 3390
rect 8988 26290 9044 26292
rect 8988 26238 8990 26290
rect 8990 26238 9042 26290
rect 9042 26238 9044 26290
rect 8988 26236 9044 26238
rect 10668 28530 10724 28532
rect 10668 28478 10670 28530
rect 10670 28478 10722 28530
rect 10722 28478 10724 28530
rect 10668 28476 10724 28478
rect 10108 27804 10164 27860
rect 10780 28140 10836 28196
rect 9996 26572 10052 26628
rect 9772 26124 9828 26180
rect 10332 26572 10388 26628
rect 8988 25340 9044 25396
rect 9100 25228 9156 25284
rect 10556 26178 10612 26180
rect 10556 26126 10558 26178
rect 10558 26126 10610 26178
rect 10610 26126 10612 26178
rect 10556 26124 10612 26126
rect 10108 23884 10164 23940
rect 9996 22428 10052 22484
rect 9772 22370 9828 22372
rect 9772 22318 9774 22370
rect 9774 22318 9826 22370
rect 9826 22318 9828 22370
rect 9772 22316 9828 22318
rect 11228 32338 11284 32340
rect 11228 32286 11230 32338
rect 11230 32286 11282 32338
rect 11282 32286 11284 32338
rect 11228 32284 11284 32286
rect 11116 31948 11172 32004
rect 11116 31666 11172 31668
rect 11116 31614 11118 31666
rect 11118 31614 11170 31666
rect 11170 31614 11172 31666
rect 11116 31612 11172 31614
rect 11900 42140 11956 42196
rect 11788 42028 11844 42084
rect 11900 39730 11956 39732
rect 11900 39678 11902 39730
rect 11902 39678 11954 39730
rect 11954 39678 11956 39730
rect 11900 39676 11956 39678
rect 11564 37324 11620 37380
rect 11564 36540 11620 36596
rect 12124 39116 12180 39172
rect 12012 36428 12068 36484
rect 11788 35980 11844 36036
rect 11900 33292 11956 33348
rect 11676 33068 11732 33124
rect 11452 32620 11508 32676
rect 11340 30098 11396 30100
rect 11340 30046 11342 30098
rect 11342 30046 11394 30098
rect 11394 30046 11396 30098
rect 11340 30044 11396 30046
rect 11452 29932 11508 29988
rect 11004 28252 11060 28308
rect 12908 44322 12964 44324
rect 12908 44270 12910 44322
rect 12910 44270 12962 44322
rect 12962 44270 12964 44322
rect 12908 44268 12964 44270
rect 12348 44044 12404 44100
rect 12348 42028 12404 42084
rect 12348 39116 12404 39172
rect 12796 43538 12852 43540
rect 12796 43486 12798 43538
rect 12798 43486 12850 43538
rect 12850 43486 12852 43538
rect 12796 43484 12852 43486
rect 13244 53676 13300 53732
rect 14924 62076 14980 62132
rect 14812 60620 14868 60676
rect 14700 57650 14756 57652
rect 14700 57598 14702 57650
rect 14702 57598 14754 57650
rect 14754 57598 14756 57650
rect 14700 57596 14756 57598
rect 14588 57036 14644 57092
rect 14924 56364 14980 56420
rect 14476 54796 14532 54852
rect 14252 54572 14308 54628
rect 14140 54124 14196 54180
rect 14028 53564 14084 53620
rect 13580 53116 13636 53172
rect 13356 52162 13412 52164
rect 13356 52110 13358 52162
rect 13358 52110 13410 52162
rect 13410 52110 13412 52162
rect 13356 52108 13412 52110
rect 13580 52108 13636 52164
rect 15596 63644 15652 63700
rect 15260 62636 15316 62692
rect 15596 62300 15652 62356
rect 15372 62188 15428 62244
rect 15484 61570 15540 61572
rect 15484 61518 15486 61570
rect 15486 61518 15538 61570
rect 15538 61518 15540 61570
rect 15484 61516 15540 61518
rect 15372 61068 15428 61124
rect 15260 60732 15316 60788
rect 15260 57932 15316 57988
rect 15260 57596 15316 57652
rect 15036 54572 15092 54628
rect 15148 57484 15204 57540
rect 14924 54124 14980 54180
rect 14812 53730 14868 53732
rect 14812 53678 14814 53730
rect 14814 53678 14866 53730
rect 14866 53678 14868 53730
rect 14812 53676 14868 53678
rect 13916 52108 13972 52164
rect 13916 50988 13972 51044
rect 13468 49868 13524 49924
rect 13804 49810 13860 49812
rect 13804 49758 13806 49810
rect 13806 49758 13858 49810
rect 13858 49758 13860 49810
rect 13804 49756 13860 49758
rect 13804 48914 13860 48916
rect 13804 48862 13806 48914
rect 13806 48862 13858 48914
rect 13858 48862 13860 48914
rect 13804 48860 13860 48862
rect 13580 48300 13636 48356
rect 13804 48636 13860 48692
rect 13356 47740 13412 47796
rect 13580 48076 13636 48132
rect 13356 47068 13412 47124
rect 13468 46898 13524 46900
rect 13468 46846 13470 46898
rect 13470 46846 13522 46898
rect 13522 46846 13524 46898
rect 13468 46844 13524 46846
rect 13356 45276 13412 45332
rect 14700 53564 14756 53620
rect 14140 52946 14196 52948
rect 14140 52894 14142 52946
rect 14142 52894 14194 52946
rect 14194 52894 14196 52946
rect 14140 52892 14196 52894
rect 14476 52946 14532 52948
rect 14476 52894 14478 52946
rect 14478 52894 14530 52946
rect 14530 52894 14532 52946
rect 14476 52892 14532 52894
rect 14140 48860 14196 48916
rect 14252 48802 14308 48804
rect 14252 48750 14254 48802
rect 14254 48750 14306 48802
rect 14306 48750 14308 48802
rect 14252 48748 14308 48750
rect 13692 46844 13748 46900
rect 14140 45890 14196 45892
rect 14140 45838 14142 45890
rect 14142 45838 14194 45890
rect 14194 45838 14196 45890
rect 14140 45836 14196 45838
rect 13692 45724 13748 45780
rect 14476 45778 14532 45780
rect 14476 45726 14478 45778
rect 14478 45726 14530 45778
rect 14530 45726 14532 45778
rect 14476 45724 14532 45726
rect 14140 44828 14196 44884
rect 13580 44268 13636 44324
rect 13916 44380 13972 44436
rect 13356 44044 13412 44100
rect 13804 44156 13860 44212
rect 13356 43708 13412 43764
rect 12796 42866 12852 42868
rect 12796 42814 12798 42866
rect 12798 42814 12850 42866
rect 12850 42814 12852 42866
rect 12796 42812 12852 42814
rect 12908 42028 12964 42084
rect 13468 43484 13524 43540
rect 14028 43538 14084 43540
rect 14028 43486 14030 43538
rect 14030 43486 14082 43538
rect 14082 43486 14084 43538
rect 14028 43484 14084 43486
rect 14588 45330 14644 45332
rect 14588 45278 14590 45330
rect 14590 45278 14642 45330
rect 14642 45278 14644 45330
rect 14588 45276 14644 45278
rect 14588 44604 14644 44660
rect 14588 44156 14644 44212
rect 14812 45890 14868 45892
rect 14812 45838 14814 45890
rect 14814 45838 14866 45890
rect 14866 45838 14868 45890
rect 14812 45836 14868 45838
rect 14476 43932 14532 43988
rect 13468 39618 13524 39620
rect 13468 39566 13470 39618
rect 13470 39566 13522 39618
rect 13522 39566 13524 39618
rect 13468 39564 13524 39566
rect 13468 38892 13524 38948
rect 12572 36594 12628 36596
rect 12572 36542 12574 36594
rect 12574 36542 12626 36594
rect 12626 36542 12628 36594
rect 12572 36540 12628 36542
rect 12236 34076 12292 34132
rect 12460 34636 12516 34692
rect 12236 33346 12292 33348
rect 12236 33294 12238 33346
rect 12238 33294 12290 33346
rect 12290 33294 12292 33346
rect 12236 33292 12292 33294
rect 12124 33068 12180 33124
rect 12684 34188 12740 34244
rect 12572 33404 12628 33460
rect 12684 33292 12740 33348
rect 12348 32562 12404 32564
rect 12348 32510 12350 32562
rect 12350 32510 12402 32562
rect 12402 32510 12404 32562
rect 12348 32508 12404 32510
rect 12348 31948 12404 32004
rect 11788 30882 11844 30884
rect 11788 30830 11790 30882
rect 11790 30830 11842 30882
rect 11842 30830 11844 30882
rect 11788 30828 11844 30830
rect 11228 29538 11284 29540
rect 11228 29486 11230 29538
rect 11230 29486 11282 29538
rect 11282 29486 11284 29538
rect 11228 29484 11284 29486
rect 11228 28700 11284 28756
rect 11116 28476 11172 28532
rect 11004 28028 11060 28084
rect 11116 27132 11172 27188
rect 11004 26962 11060 26964
rect 11004 26910 11006 26962
rect 11006 26910 11058 26962
rect 11058 26910 11060 26962
rect 11004 26908 11060 26910
rect 10332 23212 10388 23268
rect 10780 23884 10836 23940
rect 10892 25228 10948 25284
rect 10780 23660 10836 23716
rect 11116 24946 11172 24948
rect 11116 24894 11118 24946
rect 11118 24894 11170 24946
rect 11170 24894 11172 24946
rect 11116 24892 11172 24894
rect 11116 24444 11172 24500
rect 11452 29148 11508 29204
rect 12124 30940 12180 30996
rect 11900 29426 11956 29428
rect 11900 29374 11902 29426
rect 11902 29374 11954 29426
rect 11954 29374 11956 29426
rect 11900 29372 11956 29374
rect 13132 33292 13188 33348
rect 13804 38556 13860 38612
rect 12796 31612 12852 31668
rect 13356 31948 13412 32004
rect 11564 28588 11620 28644
rect 11564 28140 11620 28196
rect 11788 28028 11844 28084
rect 11788 27580 11844 27636
rect 12236 28140 12292 28196
rect 12348 28082 12404 28084
rect 12348 28030 12350 28082
rect 12350 28030 12402 28082
rect 12402 28030 12404 28082
rect 12348 28028 12404 28030
rect 12796 28140 12852 28196
rect 12012 27858 12068 27860
rect 12012 27806 12014 27858
rect 12014 27806 12066 27858
rect 12066 27806 12068 27858
rect 12012 27804 12068 27806
rect 12012 27132 12068 27188
rect 12124 26852 12180 26908
rect 12348 27804 12404 27860
rect 12460 27746 12516 27748
rect 12460 27694 12462 27746
rect 12462 27694 12514 27746
rect 12514 27694 12516 27746
rect 12460 27692 12516 27694
rect 12348 27132 12404 27188
rect 12796 27580 12852 27636
rect 13020 27132 13076 27188
rect 12684 26908 12740 26964
rect 12572 26850 12628 26852
rect 12572 26798 12574 26850
rect 12574 26798 12626 26850
rect 12626 26798 12628 26850
rect 12572 26796 12628 26798
rect 11788 25340 11844 25396
rect 11452 24444 11508 24500
rect 11788 24892 11844 24948
rect 10220 23100 10276 23156
rect 10780 22988 10836 23044
rect 9884 21756 9940 21812
rect 9212 18396 9268 18452
rect 10892 21810 10948 21812
rect 10892 21758 10894 21810
rect 10894 21758 10946 21810
rect 10946 21758 10948 21810
rect 10892 21756 10948 21758
rect 9884 19852 9940 19908
rect 9996 19794 10052 19796
rect 9996 19742 9998 19794
rect 9998 19742 10050 19794
rect 10050 19742 10052 19794
rect 9996 19740 10052 19742
rect 9884 18508 9940 18564
rect 9772 18396 9828 18452
rect 11116 22428 11172 22484
rect 11340 23714 11396 23716
rect 11340 23662 11342 23714
rect 11342 23662 11394 23714
rect 11394 23662 11396 23714
rect 11340 23660 11396 23662
rect 11004 20076 11060 20132
rect 11340 23212 11396 23268
rect 11116 19906 11172 19908
rect 11116 19854 11118 19906
rect 11118 19854 11170 19906
rect 11170 19854 11172 19906
rect 11116 19852 11172 19854
rect 11228 20524 11284 20580
rect 10556 19740 10612 19796
rect 10444 19180 10500 19236
rect 10444 18620 10500 18676
rect 10332 18450 10388 18452
rect 10332 18398 10334 18450
rect 10334 18398 10386 18450
rect 10386 18398 10388 18450
rect 10332 18396 10388 18398
rect 11676 23100 11732 23156
rect 12460 25282 12516 25284
rect 12460 25230 12462 25282
rect 12462 25230 12514 25282
rect 12514 25230 12516 25282
rect 12460 25228 12516 25230
rect 11788 22482 11844 22484
rect 11788 22430 11790 22482
rect 11790 22430 11842 22482
rect 11842 22430 11844 22482
rect 11788 22428 11844 22430
rect 11900 22370 11956 22372
rect 11900 22318 11902 22370
rect 11902 22318 11954 22370
rect 11954 22318 11956 22370
rect 11900 22316 11956 22318
rect 12236 23996 12292 24052
rect 12124 23938 12180 23940
rect 12124 23886 12126 23938
rect 12126 23886 12178 23938
rect 12178 23886 12180 23938
rect 12124 23884 12180 23886
rect 13020 26908 13076 26964
rect 12796 23884 12852 23940
rect 13244 27692 13300 27748
rect 12796 23154 12852 23156
rect 12796 23102 12798 23154
rect 12798 23102 12850 23154
rect 12850 23102 12852 23154
rect 12796 23100 12852 23102
rect 13132 23212 13188 23268
rect 12684 22988 12740 23044
rect 11452 21810 11508 21812
rect 11452 21758 11454 21810
rect 11454 21758 11506 21810
rect 11506 21758 11508 21810
rect 11452 21756 11508 21758
rect 14252 37100 14308 37156
rect 14700 39004 14756 39060
rect 15596 61068 15652 61124
rect 15596 60786 15652 60788
rect 15596 60734 15598 60786
rect 15598 60734 15650 60786
rect 15650 60734 15652 60786
rect 15596 60732 15652 60734
rect 15484 57650 15540 57652
rect 15484 57598 15486 57650
rect 15486 57598 15538 57650
rect 15538 57598 15540 57650
rect 15484 57596 15540 57598
rect 15820 65324 15876 65380
rect 16492 65436 16548 65492
rect 16380 65378 16436 65380
rect 16380 65326 16382 65378
rect 16382 65326 16434 65378
rect 16434 65326 16436 65378
rect 16380 65324 16436 65326
rect 16044 64652 16100 64708
rect 16268 64540 16324 64596
rect 16044 63980 16100 64036
rect 16380 62914 16436 62916
rect 16380 62862 16382 62914
rect 16382 62862 16434 62914
rect 16434 62862 16436 62914
rect 16380 62860 16436 62862
rect 15932 62524 15988 62580
rect 17052 71260 17108 71316
rect 16716 64764 16772 64820
rect 16828 70082 16884 70084
rect 16828 70030 16830 70082
rect 16830 70030 16882 70082
rect 16882 70030 16884 70082
rect 16828 70028 16884 70030
rect 17164 70588 17220 70644
rect 17948 72268 18004 72324
rect 17724 71372 17780 71428
rect 17836 70588 17892 70644
rect 18508 70700 18564 70756
rect 17612 70028 17668 70084
rect 17388 67618 17444 67620
rect 17388 67566 17390 67618
rect 17390 67566 17442 67618
rect 17442 67566 17444 67618
rect 17388 67564 17444 67566
rect 17276 66892 17332 66948
rect 17500 66892 17556 66948
rect 17388 66220 17444 66276
rect 18284 70364 18340 70420
rect 18396 70588 18452 70644
rect 18732 70364 18788 70420
rect 20076 75740 20132 75796
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19180 74172 19236 74228
rect 19404 74732 19460 74788
rect 22092 76354 22148 76356
rect 22092 76302 22094 76354
rect 22094 76302 22146 76354
rect 22146 76302 22148 76354
rect 22092 76300 22148 76302
rect 20524 75404 20580 75460
rect 20636 75628 20692 75684
rect 24332 76524 24388 76580
rect 22428 75628 22484 75684
rect 23548 74898 23604 74900
rect 23548 74846 23550 74898
rect 23550 74846 23602 74898
rect 23602 74846 23604 74898
rect 23548 74844 23604 74846
rect 22764 74786 22820 74788
rect 22764 74734 22766 74786
rect 22766 74734 22818 74786
rect 22818 74734 22820 74786
rect 22764 74732 22820 74734
rect 22764 74396 22820 74452
rect 20524 74172 20580 74228
rect 23996 74898 24052 74900
rect 23996 74846 23998 74898
rect 23998 74846 24050 74898
rect 24050 74846 24052 74898
rect 23996 74844 24052 74846
rect 29372 77196 29428 77252
rect 30380 77196 30436 77252
rect 27580 76636 27636 76692
rect 29260 76636 29316 76692
rect 27244 76466 27300 76468
rect 27244 76414 27246 76466
rect 27246 76414 27298 76466
rect 27298 76414 27300 76466
rect 27244 76412 27300 76414
rect 24780 75852 24836 75908
rect 24668 74898 24724 74900
rect 24668 74846 24670 74898
rect 24670 74846 24722 74898
rect 24722 74846 24724 74898
rect 24668 74844 24724 74846
rect 24332 74396 24388 74452
rect 22316 74226 22372 74228
rect 22316 74174 22318 74226
rect 22318 74174 22370 74226
rect 22370 74174 22372 74226
rect 22316 74172 22372 74174
rect 19740 74002 19796 74004
rect 19740 73950 19742 74002
rect 19742 73950 19794 74002
rect 19794 73950 19796 74002
rect 19740 73948 19796 73950
rect 20748 74002 20804 74004
rect 20748 73950 20750 74002
rect 20750 73950 20802 74002
rect 20802 73950 20804 74002
rect 20748 73948 20804 73950
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 20636 73612 20692 73668
rect 19180 72604 19236 72660
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19404 70588 19460 70644
rect 17948 67116 18004 67172
rect 18172 67228 18228 67284
rect 17612 65660 17668 65716
rect 17276 64594 17332 64596
rect 17276 64542 17278 64594
rect 17278 64542 17330 64594
rect 17330 64542 17332 64594
rect 17276 64540 17332 64542
rect 17052 64428 17108 64484
rect 16940 63980 16996 64036
rect 16828 63196 16884 63252
rect 17276 63138 17332 63140
rect 17276 63086 17278 63138
rect 17278 63086 17330 63138
rect 17330 63086 17332 63138
rect 17276 63084 17332 63086
rect 16828 62914 16884 62916
rect 16828 62862 16830 62914
rect 16830 62862 16882 62914
rect 16882 62862 16884 62914
rect 16828 62860 16884 62862
rect 16604 62524 16660 62580
rect 15932 61068 15988 61124
rect 16044 62300 16100 62356
rect 15820 59948 15876 60004
rect 15932 60898 15988 60900
rect 15932 60846 15934 60898
rect 15934 60846 15986 60898
rect 15986 60846 15988 60898
rect 15932 60844 15988 60846
rect 16716 62300 16772 62356
rect 16492 61516 16548 61572
rect 15708 57596 15764 57652
rect 15820 57484 15876 57540
rect 15260 57148 15316 57204
rect 15708 57090 15764 57092
rect 15708 57038 15710 57090
rect 15710 57038 15762 57090
rect 15762 57038 15764 57090
rect 15708 57036 15764 57038
rect 16492 60732 16548 60788
rect 17612 65100 17668 65156
rect 17612 64482 17668 64484
rect 17612 64430 17614 64482
rect 17614 64430 17666 64482
rect 17666 64430 17668 64482
rect 17612 64428 17668 64430
rect 17836 63362 17892 63364
rect 17836 63310 17838 63362
rect 17838 63310 17890 63362
rect 17890 63310 17892 63362
rect 17836 63308 17892 63310
rect 17500 62860 17556 62916
rect 17836 62748 17892 62804
rect 17164 61180 17220 61236
rect 16940 60508 16996 60564
rect 16492 59276 16548 59332
rect 16380 58546 16436 58548
rect 16380 58494 16382 58546
rect 16382 58494 16434 58546
rect 16434 58494 16436 58546
rect 16380 58492 16436 58494
rect 16716 58492 16772 58548
rect 16940 57932 16996 57988
rect 15932 57036 15988 57092
rect 15708 56754 15764 56756
rect 15708 56702 15710 56754
rect 15710 56702 15762 56754
rect 15762 56702 15764 56754
rect 15708 56700 15764 56702
rect 16828 57650 16884 57652
rect 16828 57598 16830 57650
rect 16830 57598 16882 57650
rect 16882 57598 16884 57650
rect 16828 57596 16884 57598
rect 16828 57372 16884 57428
rect 16492 56700 16548 56756
rect 16716 57148 16772 57204
rect 15932 55186 15988 55188
rect 15932 55134 15934 55186
rect 15934 55134 15986 55186
rect 15986 55134 15988 55186
rect 15932 55132 15988 55134
rect 15484 54572 15540 54628
rect 15820 53564 15876 53620
rect 15260 52946 15316 52948
rect 15260 52894 15262 52946
rect 15262 52894 15314 52946
rect 15314 52894 15316 52946
rect 15260 52892 15316 52894
rect 15260 52668 15316 52724
rect 15372 51996 15428 52052
rect 15372 50706 15428 50708
rect 15372 50654 15374 50706
rect 15374 50654 15426 50706
rect 15426 50654 15428 50706
rect 15372 50652 15428 50654
rect 15260 49644 15316 49700
rect 15036 49532 15092 49588
rect 15260 48748 15316 48804
rect 15708 52946 15764 52948
rect 15708 52894 15710 52946
rect 15710 52894 15762 52946
rect 15762 52894 15764 52946
rect 15708 52892 15764 52894
rect 16940 56364 16996 56420
rect 17164 56140 17220 56196
rect 16940 55298 16996 55300
rect 16940 55246 16942 55298
rect 16942 55246 16994 55298
rect 16994 55246 16996 55298
rect 16940 55244 16996 55246
rect 17052 55132 17108 55188
rect 17164 55580 17220 55636
rect 18620 67170 18676 67172
rect 18620 67118 18622 67170
rect 18622 67118 18674 67170
rect 18674 67118 18676 67170
rect 18620 67116 18676 67118
rect 18172 65212 18228 65268
rect 18172 63644 18228 63700
rect 18396 64594 18452 64596
rect 18396 64542 18398 64594
rect 18398 64542 18450 64594
rect 18450 64542 18452 64594
rect 18396 64540 18452 64542
rect 18284 63532 18340 63588
rect 18396 63980 18452 64036
rect 18172 63308 18228 63364
rect 18172 62748 18228 62804
rect 19292 70252 19348 70308
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 20188 70306 20244 70308
rect 20188 70254 20190 70306
rect 20190 70254 20242 70306
rect 20242 70254 20244 70306
rect 20188 70252 20244 70254
rect 19068 67228 19124 67284
rect 18844 65266 18900 65268
rect 18844 65214 18846 65266
rect 18846 65214 18898 65266
rect 18898 65214 18900 65266
rect 18844 65212 18900 65214
rect 17948 62354 18004 62356
rect 17948 62302 17950 62354
rect 17950 62302 18002 62354
rect 18002 62302 18004 62354
rect 17948 62300 18004 62302
rect 17612 61180 17668 61236
rect 17612 60620 17668 60676
rect 17836 60620 17892 60676
rect 17276 54572 17332 54628
rect 17388 59724 17444 59780
rect 17500 59612 17556 59668
rect 19516 64428 19572 64484
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 20748 72828 20804 72884
rect 20524 70866 20580 70868
rect 20524 70814 20526 70866
rect 20526 70814 20578 70866
rect 20578 70814 20580 70866
rect 20524 70812 20580 70814
rect 20636 69580 20692 69636
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 20188 65100 20244 65156
rect 19740 64594 19796 64596
rect 19740 64542 19742 64594
rect 19742 64542 19794 64594
rect 19794 64542 19796 64594
rect 19740 64540 19796 64542
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 19180 63362 19236 63364
rect 19180 63310 19182 63362
rect 19182 63310 19234 63362
rect 19234 63310 19236 63362
rect 19180 63308 19236 63310
rect 19964 63362 20020 63364
rect 19964 63310 19966 63362
rect 19966 63310 20018 63362
rect 20018 63310 20020 63362
rect 19964 63308 20020 63310
rect 20300 63250 20356 63252
rect 20300 63198 20302 63250
rect 20302 63198 20354 63250
rect 20354 63198 20356 63250
rect 20300 63196 20356 63198
rect 18508 62188 18564 62244
rect 18844 63138 18900 63140
rect 18844 63086 18846 63138
rect 18846 63086 18898 63138
rect 18898 63086 18900 63138
rect 18844 63084 18900 63086
rect 18060 61010 18116 61012
rect 18060 60958 18062 61010
rect 18062 60958 18114 61010
rect 18114 60958 18116 61010
rect 18060 60956 18116 60958
rect 18284 60508 18340 60564
rect 18060 59724 18116 59780
rect 18060 59330 18116 59332
rect 18060 59278 18062 59330
rect 18062 59278 18114 59330
rect 18114 59278 18116 59330
rect 18060 59276 18116 59278
rect 17724 59106 17780 59108
rect 17724 59054 17726 59106
rect 17726 59054 17778 59106
rect 17778 59054 17780 59106
rect 17724 59052 17780 59054
rect 17500 57762 17556 57764
rect 17500 57710 17502 57762
rect 17502 57710 17554 57762
rect 17554 57710 17556 57762
rect 17500 57708 17556 57710
rect 17612 57650 17668 57652
rect 17612 57598 17614 57650
rect 17614 57598 17666 57650
rect 17666 57598 17668 57650
rect 17612 57596 17668 57598
rect 17500 56194 17556 56196
rect 17500 56142 17502 56194
rect 17502 56142 17554 56194
rect 17554 56142 17556 56194
rect 17500 56140 17556 56142
rect 18172 59164 18228 59220
rect 17836 57596 17892 57652
rect 18060 58434 18116 58436
rect 18060 58382 18062 58434
rect 18062 58382 18114 58434
rect 18114 58382 18116 58434
rect 18060 58380 18116 58382
rect 18508 61852 18564 61908
rect 18620 61180 18676 61236
rect 19404 62860 19460 62916
rect 19740 62914 19796 62916
rect 19740 62862 19742 62914
rect 19742 62862 19794 62914
rect 19794 62862 19796 62914
rect 19740 62860 19796 62862
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 18508 60786 18564 60788
rect 18508 60734 18510 60786
rect 18510 60734 18562 60786
rect 18562 60734 18564 60786
rect 18508 60732 18564 60734
rect 18396 58716 18452 58772
rect 18844 62242 18900 62244
rect 18844 62190 18846 62242
rect 18846 62190 18898 62242
rect 18898 62190 18900 62242
rect 18844 62188 18900 62190
rect 19404 61852 19460 61908
rect 20300 62188 20356 62244
rect 20860 65436 20916 65492
rect 20748 65324 20804 65380
rect 20972 64540 21028 64596
rect 20636 64428 20692 64484
rect 21644 72434 21700 72436
rect 21644 72382 21646 72434
rect 21646 72382 21698 72434
rect 21698 72382 21700 72434
rect 21644 72380 21700 72382
rect 23212 74172 23268 74228
rect 23884 74226 23940 74228
rect 23884 74174 23886 74226
rect 23886 74174 23938 74226
rect 23938 74174 23940 74226
rect 23884 74172 23940 74174
rect 22204 72380 22260 72436
rect 21980 71372 22036 71428
rect 22428 71708 22484 71764
rect 21420 70754 21476 70756
rect 21420 70702 21422 70754
rect 21422 70702 21474 70754
rect 21474 70702 21476 70754
rect 21420 70700 21476 70702
rect 22764 71708 22820 71764
rect 22652 71260 22708 71316
rect 25228 74172 25284 74228
rect 26012 74898 26068 74900
rect 26012 74846 26014 74898
rect 26014 74846 26066 74898
rect 26066 74846 26068 74898
rect 26012 74844 26068 74846
rect 26348 74284 26404 74340
rect 24780 73276 24836 73332
rect 24892 73052 24948 73108
rect 24556 72604 24612 72660
rect 23884 72268 23940 72324
rect 21420 70364 21476 70420
rect 21308 69580 21364 69636
rect 23100 71090 23156 71092
rect 23100 71038 23102 71090
rect 23102 71038 23154 71090
rect 23154 71038 23156 71090
rect 23100 71036 23156 71038
rect 23436 69916 23492 69972
rect 23660 67452 23716 67508
rect 21308 67116 21364 67172
rect 23324 67170 23380 67172
rect 23324 67118 23326 67170
rect 23326 67118 23378 67170
rect 23378 67118 23380 67170
rect 23324 67116 23380 67118
rect 21308 65100 21364 65156
rect 21756 66108 21812 66164
rect 22428 66162 22484 66164
rect 22428 66110 22430 66162
rect 22430 66110 22482 66162
rect 22482 66110 22484 66162
rect 22428 66108 22484 66110
rect 22092 65490 22148 65492
rect 22092 65438 22094 65490
rect 22094 65438 22146 65490
rect 22146 65438 22148 65490
rect 22092 65436 22148 65438
rect 22988 65324 23044 65380
rect 22092 64706 22148 64708
rect 22092 64654 22094 64706
rect 22094 64654 22146 64706
rect 22146 64654 22148 64706
rect 22092 64652 22148 64654
rect 21868 64594 21924 64596
rect 21868 64542 21870 64594
rect 21870 64542 21922 64594
rect 21922 64542 21924 64594
rect 21868 64540 21924 64542
rect 23660 64428 23716 64484
rect 21644 63196 21700 63252
rect 21532 62860 21588 62916
rect 18956 61570 19012 61572
rect 18956 61518 18958 61570
rect 18958 61518 19010 61570
rect 19010 61518 19012 61570
rect 18956 61516 19012 61518
rect 18844 61292 18900 61348
rect 19516 61458 19572 61460
rect 19516 61406 19518 61458
rect 19518 61406 19570 61458
rect 19570 61406 19572 61458
rect 19516 61404 19572 61406
rect 19292 61346 19348 61348
rect 19292 61294 19294 61346
rect 19294 61294 19346 61346
rect 19346 61294 19348 61346
rect 19292 61292 19348 61294
rect 19180 61180 19236 61236
rect 19516 61180 19572 61236
rect 19836 61178 19892 61180
rect 18732 60508 18788 60564
rect 19068 61068 19124 61124
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 18956 58716 19012 58772
rect 17612 54626 17668 54628
rect 17612 54574 17614 54626
rect 17614 54574 17666 54626
rect 17666 54574 17668 54626
rect 17612 54572 17668 54574
rect 17948 55580 18004 55636
rect 18172 56140 18228 56196
rect 17948 54738 18004 54740
rect 17948 54686 17950 54738
rect 17950 54686 18002 54738
rect 18002 54686 18004 54738
rect 17948 54684 18004 54686
rect 18620 58380 18676 58436
rect 18508 56924 18564 56980
rect 18396 55804 18452 55860
rect 18396 55244 18452 55300
rect 16268 53618 16324 53620
rect 16268 53566 16270 53618
rect 16270 53566 16322 53618
rect 16322 53566 16324 53618
rect 16268 53564 16324 53566
rect 16380 53452 16436 53508
rect 15596 49810 15652 49812
rect 15596 49758 15598 49810
rect 15598 49758 15650 49810
rect 15650 49758 15652 49810
rect 15596 49756 15652 49758
rect 16604 52946 16660 52948
rect 16604 52894 16606 52946
rect 16606 52894 16658 52946
rect 16658 52894 16660 52946
rect 16604 52892 16660 52894
rect 16604 52556 16660 52612
rect 15932 50092 15988 50148
rect 16156 52220 16212 52276
rect 15484 46844 15540 46900
rect 15596 49308 15652 49364
rect 15036 45836 15092 45892
rect 15708 49026 15764 49028
rect 15708 48974 15710 49026
rect 15710 48974 15762 49026
rect 15762 48974 15764 49026
rect 15708 48972 15764 48974
rect 16380 50092 16436 50148
rect 16156 49644 16212 49700
rect 15820 48748 15876 48804
rect 16044 49084 16100 49140
rect 15148 45276 15204 45332
rect 15260 45388 15316 45444
rect 15708 46956 15764 47012
rect 15932 46844 15988 46900
rect 15708 46172 15764 46228
rect 15036 43932 15092 43988
rect 15372 43708 15428 43764
rect 15596 45666 15652 45668
rect 15596 45614 15598 45666
rect 15598 45614 15650 45666
rect 15650 45614 15652 45666
rect 15596 45612 15652 45614
rect 15820 46396 15876 46452
rect 15932 45948 15988 46004
rect 16268 49586 16324 49588
rect 16268 49534 16270 49586
rect 16270 49534 16322 49586
rect 16322 49534 16324 49586
rect 16268 49532 16324 49534
rect 16268 48860 16324 48916
rect 16156 48748 16212 48804
rect 15708 45388 15764 45444
rect 15708 45106 15764 45108
rect 15708 45054 15710 45106
rect 15710 45054 15762 45106
rect 15762 45054 15764 45106
rect 15708 45052 15764 45054
rect 16604 45724 16660 45780
rect 17052 50652 17108 50708
rect 17724 53452 17780 53508
rect 18732 57372 18788 57428
rect 18956 57426 19012 57428
rect 18956 57374 18958 57426
rect 18958 57374 19010 57426
rect 19010 57374 19012 57426
rect 18956 57372 19012 57374
rect 19180 60674 19236 60676
rect 19180 60622 19182 60674
rect 19182 60622 19234 60674
rect 19234 60622 19236 60674
rect 19180 60620 19236 60622
rect 19964 60620 20020 60676
rect 19292 60060 19348 60116
rect 19852 60002 19908 60004
rect 19852 59950 19854 60002
rect 19854 59950 19906 60002
rect 19906 59950 19908 60002
rect 19852 59948 19908 59950
rect 20300 59948 20356 60004
rect 20524 61292 20580 61348
rect 20524 60956 20580 61012
rect 20412 60620 20468 60676
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19628 59218 19684 59220
rect 19628 59166 19630 59218
rect 19630 59166 19682 59218
rect 19682 59166 19684 59218
rect 19628 59164 19684 59166
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19964 57650 20020 57652
rect 19964 57598 19966 57650
rect 19966 57598 20018 57650
rect 20018 57598 20020 57650
rect 19964 57596 20020 57598
rect 20524 59890 20580 59892
rect 20524 59838 20526 59890
rect 20526 59838 20578 59890
rect 20578 59838 20580 59890
rect 20524 59836 20580 59838
rect 20636 59052 20692 59108
rect 20524 58156 20580 58212
rect 19404 57372 19460 57428
rect 18956 56364 19012 56420
rect 18732 55858 18788 55860
rect 18732 55806 18734 55858
rect 18734 55806 18786 55858
rect 18786 55806 18788 55858
rect 18732 55804 18788 55806
rect 19068 55858 19124 55860
rect 19068 55806 19070 55858
rect 19070 55806 19122 55858
rect 19122 55806 19124 55858
rect 19068 55804 19124 55806
rect 19180 55580 19236 55636
rect 19852 57036 19908 57092
rect 20188 57148 20244 57204
rect 18620 53506 18676 53508
rect 18620 53454 18622 53506
rect 18622 53454 18674 53506
rect 18674 53454 18676 53506
rect 18620 53452 18676 53454
rect 18508 52946 18564 52948
rect 18508 52894 18510 52946
rect 18510 52894 18562 52946
rect 18562 52894 18564 52946
rect 18508 52892 18564 52894
rect 17836 51660 17892 51716
rect 18396 52444 18452 52500
rect 17612 49980 17668 50036
rect 17948 50034 18004 50036
rect 17948 49982 17950 50034
rect 17950 49982 18002 50034
rect 18002 49982 18004 50034
rect 17948 49980 18004 49982
rect 19180 53900 19236 53956
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20076 55020 20132 55076
rect 20188 55804 20244 55860
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 20636 56194 20692 56196
rect 20636 56142 20638 56194
rect 20638 56142 20690 56194
rect 20690 56142 20692 56194
rect 20636 56140 20692 56142
rect 20412 55356 20468 55412
rect 20300 55132 20356 55188
rect 20188 54236 20244 54292
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19852 52892 19908 52948
rect 19180 52780 19236 52836
rect 19068 52108 19124 52164
rect 18844 52050 18900 52052
rect 18844 51998 18846 52050
rect 18846 51998 18898 52050
rect 18898 51998 18900 52050
rect 18844 51996 18900 51998
rect 18956 51772 19012 51828
rect 18732 51660 18788 51716
rect 18620 50876 18676 50932
rect 18508 50540 18564 50596
rect 18956 50988 19012 51044
rect 17724 49308 17780 49364
rect 17724 47516 17780 47572
rect 17500 46898 17556 46900
rect 17500 46846 17502 46898
rect 17502 46846 17554 46898
rect 17554 46846 17556 46898
rect 17500 46844 17556 46846
rect 16716 45276 16772 45332
rect 16380 44322 16436 44324
rect 16380 44270 16382 44322
rect 16382 44270 16434 44322
rect 16434 44270 16436 44322
rect 16380 44268 16436 44270
rect 15260 43484 15316 43540
rect 15596 42812 15652 42868
rect 15036 42252 15092 42308
rect 15484 42252 15540 42308
rect 15596 41804 15652 41860
rect 15932 42364 15988 42420
rect 16044 42028 16100 42084
rect 15484 40962 15540 40964
rect 15484 40910 15486 40962
rect 15486 40910 15538 40962
rect 15538 40910 15540 40962
rect 15484 40908 15540 40910
rect 14924 38556 14980 38612
rect 15484 38946 15540 38948
rect 15484 38894 15486 38946
rect 15486 38894 15538 38946
rect 15538 38894 15540 38946
rect 15484 38892 15540 38894
rect 15820 38780 15876 38836
rect 16604 44492 16660 44548
rect 16604 43708 16660 43764
rect 16716 45052 16772 45108
rect 16828 44156 16884 44212
rect 17500 46450 17556 46452
rect 17500 46398 17502 46450
rect 17502 46398 17554 46450
rect 17554 46398 17556 46450
rect 17500 46396 17556 46398
rect 17164 46002 17220 46004
rect 17164 45950 17166 46002
rect 17166 45950 17218 46002
rect 17218 45950 17220 46002
rect 17164 45948 17220 45950
rect 17948 48354 18004 48356
rect 17948 48302 17950 48354
rect 17950 48302 18002 48354
rect 18002 48302 18004 48354
rect 17948 48300 18004 48302
rect 18060 48018 18116 48020
rect 18060 47966 18062 48018
rect 18062 47966 18114 48018
rect 18114 47966 18116 48018
rect 18060 47964 18116 47966
rect 18396 49196 18452 49252
rect 17836 45276 17892 45332
rect 17500 45106 17556 45108
rect 17500 45054 17502 45106
rect 17502 45054 17554 45106
rect 17554 45054 17556 45106
rect 17500 45052 17556 45054
rect 17052 44268 17108 44324
rect 17836 44322 17892 44324
rect 17836 44270 17838 44322
rect 17838 44270 17890 44322
rect 17890 44270 17892 44322
rect 17836 44268 17892 44270
rect 17500 44156 17556 44212
rect 18844 50034 18900 50036
rect 18844 49982 18846 50034
rect 18846 49982 18898 50034
rect 18898 49982 18900 50034
rect 18844 49980 18900 49982
rect 18620 49308 18676 49364
rect 18620 49026 18676 49028
rect 18620 48974 18622 49026
rect 18622 48974 18674 49026
rect 18674 48974 18676 49026
rect 18620 48972 18676 48974
rect 18620 48130 18676 48132
rect 18620 48078 18622 48130
rect 18622 48078 18674 48130
rect 18674 48078 18676 48130
rect 18620 48076 18676 48078
rect 19852 52162 19908 52164
rect 19852 52110 19854 52162
rect 19854 52110 19906 52162
rect 19906 52110 19908 52162
rect 19852 52108 19908 52110
rect 19404 51938 19460 51940
rect 19404 51886 19406 51938
rect 19406 51886 19458 51938
rect 19458 51886 19460 51938
rect 19404 51884 19460 51886
rect 19516 51772 19572 51828
rect 19068 50594 19124 50596
rect 19068 50542 19070 50594
rect 19070 50542 19122 50594
rect 19122 50542 19124 50594
rect 19068 50540 19124 50542
rect 19404 50540 19460 50596
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20076 50876 20132 50932
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19068 49532 19124 49588
rect 18396 45276 18452 45332
rect 18060 44828 18116 44884
rect 19068 46844 19124 46900
rect 18956 45612 19012 45668
rect 18732 44268 18788 44324
rect 19740 49810 19796 49812
rect 19740 49758 19742 49810
rect 19742 49758 19794 49810
rect 19794 49758 19796 49810
rect 19740 49756 19796 49758
rect 19628 49308 19684 49364
rect 19404 48972 19460 49028
rect 20524 53676 20580 53732
rect 20748 53340 20804 53396
rect 20524 53116 20580 53172
rect 20300 52556 20356 52612
rect 20748 52892 20804 52948
rect 20972 61628 21028 61684
rect 21644 61404 21700 61460
rect 22876 62188 22932 62244
rect 22652 61292 22708 61348
rect 22540 60844 22596 60900
rect 21756 60786 21812 60788
rect 21756 60734 21758 60786
rect 21758 60734 21810 60786
rect 21810 60734 21812 60786
rect 21756 60732 21812 60734
rect 21308 60674 21364 60676
rect 21308 60622 21310 60674
rect 21310 60622 21362 60674
rect 21362 60622 21364 60674
rect 21308 60620 21364 60622
rect 22092 60060 22148 60116
rect 21644 60002 21700 60004
rect 21644 59950 21646 60002
rect 21646 59950 21698 60002
rect 21698 59950 21700 60002
rect 21644 59948 21700 59950
rect 22316 59890 22372 59892
rect 22316 59838 22318 59890
rect 22318 59838 22370 59890
rect 22370 59838 22372 59890
rect 22316 59836 22372 59838
rect 22764 60060 22820 60116
rect 22764 59890 22820 59892
rect 22764 59838 22766 59890
rect 22766 59838 22818 59890
rect 22818 59838 22820 59890
rect 22764 59836 22820 59838
rect 21868 59442 21924 59444
rect 21868 59390 21870 59442
rect 21870 59390 21922 59442
rect 21922 59390 21924 59442
rect 21868 59388 21924 59390
rect 21420 57148 21476 57204
rect 21756 57090 21812 57092
rect 21756 57038 21758 57090
rect 21758 57038 21810 57090
rect 21810 57038 21812 57090
rect 21756 57036 21812 57038
rect 22652 57820 22708 57876
rect 22204 57650 22260 57652
rect 22204 57598 22206 57650
rect 22206 57598 22258 57650
rect 22258 57598 22260 57650
rect 22204 57596 22260 57598
rect 22428 57090 22484 57092
rect 22428 57038 22430 57090
rect 22430 57038 22482 57090
rect 22482 57038 22484 57090
rect 22428 57036 22484 57038
rect 22428 55916 22484 55972
rect 21532 55410 21588 55412
rect 21532 55358 21534 55410
rect 21534 55358 21586 55410
rect 21586 55358 21588 55410
rect 21532 55356 21588 55358
rect 22316 55298 22372 55300
rect 22316 55246 22318 55298
rect 22318 55246 22370 55298
rect 22370 55246 22372 55298
rect 22316 55244 22372 55246
rect 21420 55132 21476 55188
rect 21980 55020 22036 55076
rect 21196 54572 21252 54628
rect 20972 54236 21028 54292
rect 24332 71762 24388 71764
rect 24332 71710 24334 71762
rect 24334 71710 24386 71762
rect 24386 71710 24388 71762
rect 24332 71708 24388 71710
rect 24220 69186 24276 69188
rect 24220 69134 24222 69186
rect 24222 69134 24274 69186
rect 24274 69134 24276 69186
rect 24220 69132 24276 69134
rect 24668 69186 24724 69188
rect 24668 69134 24670 69186
rect 24670 69134 24722 69186
rect 24722 69134 24724 69186
rect 24668 69132 24724 69134
rect 24444 67452 24500 67508
rect 23996 67116 24052 67172
rect 23884 62188 23940 62244
rect 24556 64540 24612 64596
rect 23324 60620 23380 60676
rect 23324 59836 23380 59892
rect 23100 58828 23156 58884
rect 23100 58322 23156 58324
rect 23100 58270 23102 58322
rect 23102 58270 23154 58322
rect 23154 58270 23156 58322
rect 23100 58268 23156 58270
rect 22988 55244 23044 55300
rect 23100 56924 23156 56980
rect 23548 58940 23604 58996
rect 24444 61516 24500 61572
rect 24108 60732 24164 60788
rect 24668 62242 24724 62244
rect 24668 62190 24670 62242
rect 24670 62190 24722 62242
rect 24722 62190 24724 62242
rect 24668 62188 24724 62190
rect 25004 70140 25060 70196
rect 25452 73442 25508 73444
rect 25452 73390 25454 73442
rect 25454 73390 25506 73442
rect 25506 73390 25508 73442
rect 25452 73388 25508 73390
rect 25340 72268 25396 72324
rect 25452 70082 25508 70084
rect 25452 70030 25454 70082
rect 25454 70030 25506 70082
rect 25506 70030 25508 70082
rect 25452 70028 25508 70030
rect 26236 73218 26292 73220
rect 26236 73166 26238 73218
rect 26238 73166 26290 73218
rect 26290 73166 26292 73218
rect 26236 73164 26292 73166
rect 25676 72658 25732 72660
rect 25676 72606 25678 72658
rect 25678 72606 25730 72658
rect 25730 72606 25732 72658
rect 25676 72604 25732 72606
rect 26236 72268 26292 72324
rect 27244 74732 27300 74788
rect 28588 74732 28644 74788
rect 26684 73500 26740 73556
rect 26684 73052 26740 73108
rect 27692 73554 27748 73556
rect 27692 73502 27694 73554
rect 27694 73502 27746 73554
rect 27746 73502 27748 73554
rect 27692 73500 27748 73502
rect 28028 72044 28084 72100
rect 28140 71820 28196 71876
rect 25900 70924 25956 70980
rect 25900 69580 25956 69636
rect 26908 70978 26964 70980
rect 26908 70926 26910 70978
rect 26910 70926 26962 70978
rect 26962 70926 26964 70978
rect 26908 70924 26964 70926
rect 27356 70252 27412 70308
rect 27804 70252 27860 70308
rect 27132 69804 27188 69860
rect 25676 69132 25732 69188
rect 25452 66946 25508 66948
rect 25452 66894 25454 66946
rect 25454 66894 25506 66946
rect 25506 66894 25508 66946
rect 25452 66892 25508 66894
rect 25340 64818 25396 64820
rect 25340 64766 25342 64818
rect 25342 64766 25394 64818
rect 25394 64766 25396 64818
rect 25340 64764 25396 64766
rect 25340 63532 25396 63588
rect 25452 63308 25508 63364
rect 25340 63026 25396 63028
rect 25340 62974 25342 63026
rect 25342 62974 25394 63026
rect 25394 62974 25396 63026
rect 25340 62972 25396 62974
rect 28028 69804 28084 69860
rect 26572 67004 26628 67060
rect 26684 66892 26740 66948
rect 26236 64092 26292 64148
rect 25788 63810 25844 63812
rect 25788 63758 25790 63810
rect 25790 63758 25842 63810
rect 25842 63758 25844 63810
rect 25788 63756 25844 63758
rect 26348 62972 26404 63028
rect 25340 61628 25396 61684
rect 25676 62860 25732 62916
rect 24892 61516 24948 61572
rect 24444 60620 24500 60676
rect 23996 58828 24052 58884
rect 24220 58940 24276 58996
rect 23884 58210 23940 58212
rect 23884 58158 23886 58210
rect 23886 58158 23938 58210
rect 23938 58158 23940 58210
rect 23884 58156 23940 58158
rect 23884 57820 23940 57876
rect 23212 56364 23268 56420
rect 22876 55132 22932 55188
rect 22764 55074 22820 55076
rect 22764 55022 22766 55074
rect 22766 55022 22818 55074
rect 22818 55022 22820 55074
rect 22764 55020 22820 55022
rect 22428 54738 22484 54740
rect 22428 54686 22430 54738
rect 22430 54686 22482 54738
rect 22482 54686 22484 54738
rect 22428 54684 22484 54686
rect 22316 53788 22372 53844
rect 21532 53730 21588 53732
rect 21532 53678 21534 53730
rect 21534 53678 21586 53730
rect 21586 53678 21588 53730
rect 21532 53676 21588 53678
rect 20524 51490 20580 51492
rect 20524 51438 20526 51490
rect 20526 51438 20578 51490
rect 20578 51438 20580 51490
rect 20524 51436 20580 51438
rect 20636 50316 20692 50372
rect 20412 49980 20468 50036
rect 20300 49308 20356 49364
rect 20188 48972 20244 49028
rect 19516 48914 19572 48916
rect 19516 48862 19518 48914
rect 19518 48862 19570 48914
rect 19570 48862 19572 48914
rect 19516 48860 19572 48862
rect 20188 48802 20244 48804
rect 20188 48750 20190 48802
rect 20190 48750 20242 48802
rect 20242 48750 20244 48802
rect 20188 48748 20244 48750
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19404 45276 19460 45332
rect 19516 47964 19572 48020
rect 20300 47964 20356 48020
rect 19740 47570 19796 47572
rect 19740 47518 19742 47570
rect 19742 47518 19794 47570
rect 19794 47518 19796 47570
rect 19740 47516 19796 47518
rect 20972 50316 21028 50372
rect 20636 49532 20692 49588
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20300 47234 20356 47236
rect 20300 47182 20302 47234
rect 20302 47182 20354 47234
rect 20354 47182 20356 47234
rect 20300 47180 20356 47182
rect 20748 49026 20804 49028
rect 20748 48974 20750 49026
rect 20750 48974 20802 49026
rect 20802 48974 20804 49026
rect 20748 48972 20804 48974
rect 20748 47180 20804 47236
rect 19628 45666 19684 45668
rect 19628 45614 19630 45666
rect 19630 45614 19682 45666
rect 19682 45614 19684 45666
rect 19628 45612 19684 45614
rect 20188 45666 20244 45668
rect 20188 45614 20190 45666
rect 20190 45614 20242 45666
rect 20242 45614 20244 45666
rect 20188 45612 20244 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19628 44994 19684 44996
rect 19628 44942 19630 44994
rect 19630 44942 19682 44994
rect 19682 44942 19684 44994
rect 19628 44940 19684 44942
rect 18956 43820 19012 43876
rect 19852 44882 19908 44884
rect 19852 44830 19854 44882
rect 19854 44830 19906 44882
rect 19906 44830 19908 44882
rect 19852 44828 19908 44830
rect 20748 46674 20804 46676
rect 20748 46622 20750 46674
rect 20750 46622 20802 46674
rect 20802 46622 20804 46674
rect 20748 46620 20804 46622
rect 20412 45948 20468 46004
rect 20636 46396 20692 46452
rect 20412 44940 20468 44996
rect 20524 45164 20580 45220
rect 20748 45778 20804 45780
rect 20748 45726 20750 45778
rect 20750 45726 20802 45778
rect 20802 45726 20804 45778
rect 20748 45724 20804 45726
rect 20188 44882 20244 44884
rect 20188 44830 20190 44882
rect 20190 44830 20242 44882
rect 20242 44830 20244 44882
rect 20188 44828 20244 44830
rect 20188 44604 20244 44660
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20412 44434 20468 44436
rect 20412 44382 20414 44434
rect 20414 44382 20466 44434
rect 20466 44382 20468 44434
rect 20412 44380 20468 44382
rect 20188 43820 20244 43876
rect 20300 44268 20356 44324
rect 16380 42866 16436 42868
rect 16380 42814 16382 42866
rect 16382 42814 16434 42866
rect 16434 42814 16436 42866
rect 16380 42812 16436 42814
rect 16828 43484 16884 43540
rect 16380 42252 16436 42308
rect 16492 42364 16548 42420
rect 16268 41692 16324 41748
rect 16380 41804 16436 41860
rect 16380 41186 16436 41188
rect 16380 41134 16382 41186
rect 16382 41134 16434 41186
rect 16434 41134 16436 41186
rect 16380 41132 16436 41134
rect 16156 40124 16212 40180
rect 16492 41020 16548 41076
rect 16268 39788 16324 39844
rect 16492 40236 16548 40292
rect 16268 38668 16324 38724
rect 16604 40124 16660 40180
rect 16492 39058 16548 39060
rect 16492 39006 16494 39058
rect 16494 39006 16546 39058
rect 16546 39006 16548 39058
rect 16492 39004 16548 39006
rect 14588 36988 14644 37044
rect 16268 37324 16324 37380
rect 14364 34300 14420 34356
rect 15036 37100 15092 37156
rect 13916 34242 13972 34244
rect 13916 34190 13918 34242
rect 13918 34190 13970 34242
rect 13970 34190 13972 34242
rect 13916 34188 13972 34190
rect 14364 34076 14420 34132
rect 14140 33628 14196 33684
rect 14028 33516 14084 33572
rect 13580 33234 13636 33236
rect 13580 33182 13582 33234
rect 13582 33182 13634 33234
rect 13634 33182 13636 33234
rect 13580 33180 13636 33182
rect 14476 33404 14532 33460
rect 13468 31724 13524 31780
rect 14028 30994 14084 30996
rect 14028 30942 14030 30994
rect 14030 30942 14082 30994
rect 14082 30942 14084 30994
rect 14028 30940 14084 30942
rect 14028 30380 14084 30436
rect 14140 30322 14196 30324
rect 14140 30270 14142 30322
rect 14142 30270 14194 30322
rect 14194 30270 14196 30322
rect 14140 30268 14196 30270
rect 14364 30156 14420 30212
rect 14700 33516 14756 33572
rect 14924 33740 14980 33796
rect 14588 32060 14644 32116
rect 14812 33234 14868 33236
rect 14812 33182 14814 33234
rect 14814 33182 14866 33234
rect 14866 33182 14868 33234
rect 14812 33180 14868 33182
rect 14700 31948 14756 32004
rect 14700 31612 14756 31668
rect 14924 31778 14980 31780
rect 14924 31726 14926 31778
rect 14926 31726 14978 31778
rect 14978 31726 14980 31778
rect 14924 31724 14980 31726
rect 14812 31388 14868 31444
rect 15372 37154 15428 37156
rect 15372 37102 15374 37154
rect 15374 37102 15426 37154
rect 15426 37102 15428 37154
rect 15372 37100 15428 37102
rect 16044 34914 16100 34916
rect 16044 34862 16046 34914
rect 16046 34862 16098 34914
rect 16098 34862 16100 34914
rect 16044 34860 16100 34862
rect 15932 34748 15988 34804
rect 15484 33404 15540 33460
rect 15820 33964 15876 34020
rect 16492 34242 16548 34244
rect 16492 34190 16494 34242
rect 16494 34190 16546 34242
rect 16546 34190 16548 34242
rect 16492 34188 16548 34190
rect 16268 34130 16324 34132
rect 16268 34078 16270 34130
rect 16270 34078 16322 34130
rect 16322 34078 16324 34130
rect 16268 34076 16324 34078
rect 16380 34018 16436 34020
rect 16380 33966 16382 34018
rect 16382 33966 16434 34018
rect 16434 33966 16436 34018
rect 16380 33964 16436 33966
rect 16044 33180 16100 33236
rect 15708 31890 15764 31892
rect 15708 31838 15710 31890
rect 15710 31838 15762 31890
rect 15762 31838 15764 31890
rect 15708 31836 15764 31838
rect 16156 31836 16212 31892
rect 15372 31724 15428 31780
rect 15036 31276 15092 31332
rect 15260 31276 15316 31332
rect 15148 30322 15204 30324
rect 15148 30270 15150 30322
rect 15150 30270 15202 30322
rect 15202 30270 15204 30322
rect 15148 30268 15204 30270
rect 14812 30210 14868 30212
rect 14812 30158 14814 30210
rect 14814 30158 14866 30210
rect 14866 30158 14868 30210
rect 14812 30156 14868 30158
rect 14588 29986 14644 29988
rect 14588 29934 14590 29986
rect 14590 29934 14642 29986
rect 14642 29934 14644 29986
rect 14588 29932 14644 29934
rect 14700 29538 14756 29540
rect 14700 29486 14702 29538
rect 14702 29486 14754 29538
rect 14754 29486 14756 29538
rect 14700 29484 14756 29486
rect 15372 30882 15428 30884
rect 15372 30830 15374 30882
rect 15374 30830 15426 30882
rect 15426 30830 15428 30882
rect 15372 30828 15428 30830
rect 16044 31052 16100 31108
rect 16380 30940 16436 30996
rect 16268 30828 16324 30884
rect 18620 43260 18676 43316
rect 18844 42476 18900 42532
rect 19180 43314 19236 43316
rect 19180 43262 19182 43314
rect 19182 43262 19234 43314
rect 19234 43262 19236 43314
rect 19180 43260 19236 43262
rect 17276 41186 17332 41188
rect 17276 41134 17278 41186
rect 17278 41134 17330 41186
rect 17330 41134 17332 41186
rect 17276 41132 17332 41134
rect 17052 40796 17108 40852
rect 18060 40796 18116 40852
rect 17500 40572 17556 40628
rect 17500 40236 17556 40292
rect 17276 40124 17332 40180
rect 16940 39788 16996 39844
rect 16716 36876 16772 36932
rect 16716 34972 16772 35028
rect 16828 33628 16884 33684
rect 17052 35308 17108 35364
rect 18956 41916 19012 41972
rect 19852 43260 19908 43316
rect 20076 42642 20132 42644
rect 20076 42590 20078 42642
rect 20078 42590 20130 42642
rect 20130 42590 20132 42642
rect 20076 42588 20132 42590
rect 19740 42530 19796 42532
rect 19740 42478 19742 42530
rect 19742 42478 19794 42530
rect 19794 42478 19796 42530
rect 19740 42476 19796 42478
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19628 41970 19684 41972
rect 19628 41918 19630 41970
rect 19630 41918 19682 41970
rect 19682 41918 19684 41970
rect 19628 41916 19684 41918
rect 18620 38556 18676 38612
rect 17836 36764 17892 36820
rect 18060 37490 18116 37492
rect 18060 37438 18062 37490
rect 18062 37438 18114 37490
rect 18114 37438 18116 37490
rect 18060 37436 18116 37438
rect 17500 35868 17556 35924
rect 18508 37490 18564 37492
rect 18508 37438 18510 37490
rect 18510 37438 18562 37490
rect 18562 37438 18564 37490
rect 18508 37436 18564 37438
rect 18956 41132 19012 41188
rect 18284 36204 18340 36260
rect 17948 35810 18004 35812
rect 17948 35758 17950 35810
rect 17950 35758 18002 35810
rect 18002 35758 18004 35810
rect 17948 35756 18004 35758
rect 17724 35644 17780 35700
rect 17388 34690 17444 34692
rect 17388 34638 17390 34690
rect 17390 34638 17442 34690
rect 17442 34638 17444 34690
rect 17388 34636 17444 34638
rect 17836 35586 17892 35588
rect 17836 35534 17838 35586
rect 17838 35534 17890 35586
rect 17890 35534 17892 35586
rect 17836 35532 17892 35534
rect 18396 35420 18452 35476
rect 17836 34972 17892 35028
rect 17948 34860 18004 34916
rect 17724 34354 17780 34356
rect 17724 34302 17726 34354
rect 17726 34302 17778 34354
rect 17778 34302 17780 34354
rect 17724 34300 17780 34302
rect 17388 33740 17444 33796
rect 17052 32284 17108 32340
rect 16716 30882 16772 30884
rect 16716 30830 16718 30882
rect 16718 30830 16770 30882
rect 16770 30830 16772 30882
rect 16716 30828 16772 30830
rect 16380 30322 16436 30324
rect 16380 30270 16382 30322
rect 16382 30270 16434 30322
rect 16434 30270 16436 30322
rect 16380 30268 16436 30270
rect 15596 30210 15652 30212
rect 15596 30158 15598 30210
rect 15598 30158 15650 30210
rect 15650 30158 15652 30210
rect 15596 30156 15652 30158
rect 14028 28140 14084 28196
rect 14700 28530 14756 28532
rect 14700 28478 14702 28530
rect 14702 28478 14754 28530
rect 14754 28478 14756 28530
rect 14700 28476 14756 28478
rect 13580 27916 13636 27972
rect 14476 27970 14532 27972
rect 14476 27918 14478 27970
rect 14478 27918 14530 27970
rect 14530 27918 14532 27970
rect 14476 27916 14532 27918
rect 13804 27692 13860 27748
rect 13580 27074 13636 27076
rect 13580 27022 13582 27074
rect 13582 27022 13634 27074
rect 13634 27022 13636 27074
rect 13580 27020 13636 27022
rect 14924 28418 14980 28420
rect 14924 28366 14926 28418
rect 14926 28366 14978 28418
rect 14978 28366 14980 28418
rect 14924 28364 14980 28366
rect 15260 28364 15316 28420
rect 13916 27020 13972 27076
rect 13580 26796 13636 26852
rect 14476 26962 14532 26964
rect 14476 26910 14478 26962
rect 14478 26910 14530 26962
rect 14530 26910 14532 26962
rect 14476 26908 14532 26910
rect 14700 27132 14756 27188
rect 15260 27804 15316 27860
rect 14252 25730 14308 25732
rect 14252 25678 14254 25730
rect 14254 25678 14306 25730
rect 14306 25678 14308 25730
rect 14252 25676 14308 25678
rect 14364 25452 14420 25508
rect 15148 25676 15204 25732
rect 14252 25282 14308 25284
rect 14252 25230 14254 25282
rect 14254 25230 14306 25282
rect 14306 25230 14308 25282
rect 14252 25228 14308 25230
rect 14700 25228 14756 25284
rect 13356 22316 13412 22372
rect 14028 24332 14084 24388
rect 13804 23548 13860 23604
rect 12124 20524 12180 20580
rect 12684 20860 12740 20916
rect 11004 18562 11060 18564
rect 11004 18510 11006 18562
rect 11006 18510 11058 18562
rect 11058 18510 11060 18562
rect 11004 18508 11060 18510
rect 11116 18396 11172 18452
rect 11564 19180 11620 19236
rect 11340 19122 11396 19124
rect 11340 19070 11342 19122
rect 11342 19070 11394 19122
rect 11394 19070 11396 19122
rect 11340 19068 11396 19070
rect 11452 19010 11508 19012
rect 11452 18958 11454 19010
rect 11454 18958 11506 19010
rect 11506 18958 11508 19010
rect 11452 18956 11508 18958
rect 11004 18284 11060 18340
rect 9548 17500 9604 17556
rect 11116 17500 11172 17556
rect 11340 18226 11396 18228
rect 11340 18174 11342 18226
rect 11342 18174 11394 18226
rect 11394 18174 11396 18226
rect 11340 18172 11396 18174
rect 8988 16044 9044 16100
rect 10444 16098 10500 16100
rect 10444 16046 10446 16098
rect 10446 16046 10498 16098
rect 10498 16046 10500 16098
rect 10444 16044 10500 16046
rect 11004 15874 11060 15876
rect 11004 15822 11006 15874
rect 11006 15822 11058 15874
rect 11058 15822 11060 15874
rect 11004 15820 11060 15822
rect 11340 15596 11396 15652
rect 11676 16828 11732 16884
rect 12012 19234 12068 19236
rect 12012 19182 12014 19234
rect 12014 19182 12066 19234
rect 12066 19182 12068 19234
rect 12012 19180 12068 19182
rect 11900 18508 11956 18564
rect 12796 20130 12852 20132
rect 12796 20078 12798 20130
rect 12798 20078 12850 20130
rect 12850 20078 12852 20130
rect 12796 20076 12852 20078
rect 12124 18956 12180 19012
rect 12236 18562 12292 18564
rect 12236 18510 12238 18562
rect 12238 18510 12290 18562
rect 12290 18510 12292 18562
rect 12236 18508 12292 18510
rect 12236 18284 12292 18340
rect 11452 15426 11508 15428
rect 11452 15374 11454 15426
rect 11454 15374 11506 15426
rect 11506 15374 11508 15426
rect 11452 15372 11508 15374
rect 11564 15484 11620 15540
rect 11900 15484 11956 15540
rect 12572 19010 12628 19012
rect 12572 18958 12574 19010
rect 12574 18958 12626 19010
rect 12626 18958 12628 19010
rect 12572 18956 12628 18958
rect 12460 18172 12516 18228
rect 13916 23266 13972 23268
rect 13916 23214 13918 23266
rect 13918 23214 13970 23266
rect 13970 23214 13972 23266
rect 13916 23212 13972 23214
rect 13916 21868 13972 21924
rect 14028 19964 14084 20020
rect 13468 19122 13524 19124
rect 13468 19070 13470 19122
rect 13470 19070 13522 19122
rect 13522 19070 13524 19122
rect 13468 19068 13524 19070
rect 13692 19010 13748 19012
rect 13692 18958 13694 19010
rect 13694 18958 13746 19010
rect 13746 18958 13748 19010
rect 13692 18956 13748 18958
rect 12908 18620 12964 18676
rect 12796 18508 12852 18564
rect 13244 18450 13300 18452
rect 13244 18398 13246 18450
rect 13246 18398 13298 18450
rect 13298 18398 13300 18450
rect 13244 18396 13300 18398
rect 12348 16828 12404 16884
rect 12348 15874 12404 15876
rect 12348 15822 12350 15874
rect 12350 15822 12402 15874
rect 12402 15822 12404 15874
rect 12348 15820 12404 15822
rect 12348 15596 12404 15652
rect 11900 14252 11956 14308
rect 12572 15538 12628 15540
rect 12572 15486 12574 15538
rect 12574 15486 12626 15538
rect 12626 15486 12628 15538
rect 12572 15484 12628 15486
rect 12572 14530 12628 14532
rect 12572 14478 12574 14530
rect 12574 14478 12626 14530
rect 12626 14478 12628 14530
rect 12572 14476 12628 14478
rect 12348 13580 12404 13636
rect 11228 11676 11284 11732
rect 11340 11282 11396 11284
rect 11340 11230 11342 11282
rect 11342 11230 11394 11282
rect 11394 11230 11396 11282
rect 11340 11228 11396 11230
rect 12236 12962 12292 12964
rect 12236 12910 12238 12962
rect 12238 12910 12290 12962
rect 12290 12910 12292 12962
rect 12236 12908 12292 12910
rect 12796 12908 12852 12964
rect 13132 15596 13188 15652
rect 13020 15426 13076 15428
rect 13020 15374 13022 15426
rect 13022 15374 13074 15426
rect 13074 15374 13076 15426
rect 13020 15372 13076 15374
rect 13020 14252 13076 14308
rect 12908 13916 12964 13972
rect 13692 17666 13748 17668
rect 13692 17614 13694 17666
rect 13694 17614 13746 17666
rect 13746 17614 13748 17666
rect 13692 17612 13748 17614
rect 14588 23548 14644 23604
rect 14364 22876 14420 22932
rect 14364 18396 14420 18452
rect 14140 17724 14196 17780
rect 14588 22988 14644 23044
rect 14588 22428 14644 22484
rect 14924 22988 14980 23044
rect 15036 25116 15092 25172
rect 14812 22876 14868 22932
rect 15036 22652 15092 22708
rect 14700 22540 14756 22596
rect 14924 21810 14980 21812
rect 14924 21758 14926 21810
rect 14926 21758 14978 21810
rect 14978 21758 14980 21810
rect 14924 21756 14980 21758
rect 15036 21532 15092 21588
rect 14812 21196 14868 21252
rect 15148 21084 15204 21140
rect 15148 19404 15204 19460
rect 15036 19346 15092 19348
rect 15036 19294 15038 19346
rect 15038 19294 15090 19346
rect 15090 19294 15092 19346
rect 15036 19292 15092 19294
rect 14588 18562 14644 18564
rect 14588 18510 14590 18562
rect 14590 18510 14642 18562
rect 14642 18510 14644 18562
rect 14588 18508 14644 18510
rect 14924 18450 14980 18452
rect 14924 18398 14926 18450
rect 14926 18398 14978 18450
rect 14978 18398 14980 18450
rect 14924 18396 14980 18398
rect 14588 17778 14644 17780
rect 14588 17726 14590 17778
rect 14590 17726 14642 17778
rect 14642 17726 14644 17778
rect 14588 17724 14644 17726
rect 14476 17612 14532 17668
rect 14140 16882 14196 16884
rect 14140 16830 14142 16882
rect 14142 16830 14194 16882
rect 14194 16830 14196 16882
rect 14140 16828 14196 16830
rect 14252 16716 14308 16772
rect 13356 13804 13412 13860
rect 14140 16604 14196 16660
rect 12236 11788 12292 11844
rect 12684 12348 12740 12404
rect 12348 11676 12404 11732
rect 13020 11676 13076 11732
rect 12460 11228 12516 11284
rect 12796 11170 12852 11172
rect 12796 11118 12798 11170
rect 12798 11118 12850 11170
rect 12850 11118 12852 11170
rect 12796 11116 12852 11118
rect 13580 14418 13636 14420
rect 13580 14366 13582 14418
rect 13582 14366 13634 14418
rect 13634 14366 13636 14418
rect 13580 14364 13636 14366
rect 13468 13580 13524 13636
rect 13804 14028 13860 14084
rect 13692 12962 13748 12964
rect 13692 12910 13694 12962
rect 13694 12910 13746 12962
rect 13746 12910 13748 12962
rect 13692 12908 13748 12910
rect 13580 12850 13636 12852
rect 13580 12798 13582 12850
rect 13582 12798 13634 12850
rect 13634 12798 13636 12850
rect 13580 12796 13636 12798
rect 13356 12348 13412 12404
rect 13244 9996 13300 10052
rect 13692 12012 13748 12068
rect 12012 9772 12068 9828
rect 14476 16882 14532 16884
rect 14476 16830 14478 16882
rect 14478 16830 14530 16882
rect 14530 16830 14532 16882
rect 14476 16828 14532 16830
rect 14588 16716 14644 16772
rect 14700 17500 14756 17556
rect 15484 23548 15540 23604
rect 15596 28700 15652 28756
rect 16716 30210 16772 30212
rect 16716 30158 16718 30210
rect 16718 30158 16770 30210
rect 16770 30158 16772 30210
rect 16716 30156 16772 30158
rect 16604 29820 16660 29876
rect 16380 28700 16436 28756
rect 16604 29596 16660 29652
rect 17052 28754 17108 28756
rect 17052 28702 17054 28754
rect 17054 28702 17106 28754
rect 17106 28702 17108 28754
rect 17052 28700 17108 28702
rect 15820 27858 15876 27860
rect 15820 27806 15822 27858
rect 15822 27806 15874 27858
rect 15874 27806 15876 27858
rect 15820 27804 15876 27806
rect 15932 27074 15988 27076
rect 15932 27022 15934 27074
rect 15934 27022 15986 27074
rect 15986 27022 15988 27074
rect 15932 27020 15988 27022
rect 16156 26850 16212 26852
rect 16156 26798 16158 26850
rect 16158 26798 16210 26850
rect 16210 26798 16212 26850
rect 16156 26796 16212 26798
rect 15708 25676 15764 25732
rect 15820 26066 15876 26068
rect 15820 26014 15822 26066
rect 15822 26014 15874 26066
rect 15874 26014 15876 26066
rect 15820 26012 15876 26014
rect 16492 26460 16548 26516
rect 16604 27020 16660 27076
rect 16380 26124 16436 26180
rect 16492 26066 16548 26068
rect 16492 26014 16494 26066
rect 16494 26014 16546 26066
rect 16546 26014 16548 26066
rect 16492 26012 16548 26014
rect 16716 26460 16772 26516
rect 17052 27580 17108 27636
rect 16940 27020 16996 27076
rect 16716 23548 16772 23604
rect 15596 23266 15652 23268
rect 15596 23214 15598 23266
rect 15598 23214 15650 23266
rect 15650 23214 15652 23266
rect 15596 23212 15652 23214
rect 16156 23266 16212 23268
rect 16156 23214 16158 23266
rect 16158 23214 16210 23266
rect 16210 23214 16212 23266
rect 16156 23212 16212 23214
rect 15708 22594 15764 22596
rect 15708 22542 15710 22594
rect 15710 22542 15762 22594
rect 15762 22542 15764 22594
rect 15708 22540 15764 22542
rect 15484 22482 15540 22484
rect 15484 22430 15486 22482
rect 15486 22430 15538 22482
rect 15538 22430 15540 22482
rect 15484 22428 15540 22430
rect 15484 21308 15540 21364
rect 15820 21532 15876 21588
rect 15708 21084 15764 21140
rect 15596 20690 15652 20692
rect 15596 20638 15598 20690
rect 15598 20638 15650 20690
rect 15650 20638 15652 20690
rect 15596 20636 15652 20638
rect 15036 17724 15092 17780
rect 15260 17388 15316 17444
rect 14700 16604 14756 16660
rect 14364 16156 14420 16212
rect 15484 19404 15540 19460
rect 16828 22146 16884 22148
rect 16828 22094 16830 22146
rect 16830 22094 16882 22146
rect 16882 22094 16884 22146
rect 16828 22092 16884 22094
rect 16940 20802 16996 20804
rect 16940 20750 16942 20802
rect 16942 20750 16994 20802
rect 16994 20750 16996 20802
rect 16940 20748 16996 20750
rect 16716 20412 16772 20468
rect 15820 17388 15876 17444
rect 15932 17500 15988 17556
rect 15484 16882 15540 16884
rect 15484 16830 15486 16882
rect 15486 16830 15538 16882
rect 15538 16830 15540 16882
rect 15484 16828 15540 16830
rect 15260 16210 15316 16212
rect 15260 16158 15262 16210
rect 15262 16158 15314 16210
rect 15314 16158 15316 16210
rect 15260 16156 15316 16158
rect 14700 14642 14756 14644
rect 14700 14590 14702 14642
rect 14702 14590 14754 14642
rect 14754 14590 14756 14642
rect 14700 14588 14756 14590
rect 14588 14364 14644 14420
rect 14476 13804 14532 13860
rect 14476 13468 14532 13524
rect 14364 13356 14420 13412
rect 14028 12796 14084 12852
rect 14252 12066 14308 12068
rect 14252 12014 14254 12066
rect 14254 12014 14306 12066
rect 14306 12014 14308 12066
rect 14252 12012 14308 12014
rect 13916 11788 13972 11844
rect 13916 9100 13972 9156
rect 15148 13858 15204 13860
rect 15148 13806 15150 13858
rect 15150 13806 15202 13858
rect 15202 13806 15204 13858
rect 15148 13804 15204 13806
rect 14924 13020 14980 13076
rect 16268 18226 16324 18228
rect 16268 18174 16270 18226
rect 16270 18174 16322 18226
rect 16322 18174 16324 18226
rect 16268 18172 16324 18174
rect 16604 18172 16660 18228
rect 17500 31106 17556 31108
rect 17500 31054 17502 31106
rect 17502 31054 17554 31106
rect 17554 31054 17556 31106
rect 17500 31052 17556 31054
rect 17388 30994 17444 30996
rect 17388 30942 17390 30994
rect 17390 30942 17442 30994
rect 17442 30942 17444 30994
rect 17388 30940 17444 30942
rect 17388 30098 17444 30100
rect 17388 30046 17390 30098
rect 17390 30046 17442 30098
rect 17442 30046 17444 30098
rect 17388 30044 17444 30046
rect 17612 29986 17668 29988
rect 17612 29934 17614 29986
rect 17614 29934 17666 29986
rect 17666 29934 17668 29986
rect 17612 29932 17668 29934
rect 17276 29484 17332 29540
rect 17724 27804 17780 27860
rect 18508 34636 18564 34692
rect 18620 34860 18676 34916
rect 18172 33516 18228 33572
rect 18620 34300 18676 34356
rect 18844 38444 18900 38500
rect 18844 35868 18900 35924
rect 20972 47740 21028 47796
rect 22988 53564 23044 53620
rect 21980 52946 22036 52948
rect 21980 52894 21982 52946
rect 21982 52894 22034 52946
rect 22034 52894 22036 52946
rect 21980 52892 22036 52894
rect 21868 52780 21924 52836
rect 21420 51996 21476 52052
rect 21196 51884 21252 51940
rect 21196 50652 21252 50708
rect 21420 50540 21476 50596
rect 21420 49868 21476 49924
rect 21196 49308 21252 49364
rect 21308 48748 21364 48804
rect 21196 46620 21252 46676
rect 22652 52892 22708 52948
rect 22876 52668 22932 52724
rect 22540 52444 22596 52500
rect 22316 52162 22372 52164
rect 22316 52110 22318 52162
rect 22318 52110 22370 52162
rect 22370 52110 22372 52162
rect 22316 52108 22372 52110
rect 22316 51772 22372 51828
rect 23212 53058 23268 53060
rect 23212 53006 23214 53058
rect 23214 53006 23266 53058
rect 23266 53006 23268 53058
rect 23212 53004 23268 53006
rect 23548 52668 23604 52724
rect 22988 52444 23044 52500
rect 23212 52556 23268 52612
rect 22764 51884 22820 51940
rect 22540 51602 22596 51604
rect 22540 51550 22542 51602
rect 22542 51550 22594 51602
rect 22594 51550 22596 51602
rect 22540 51548 22596 51550
rect 22204 50594 22260 50596
rect 22204 50542 22206 50594
rect 22206 50542 22258 50594
rect 22258 50542 22260 50594
rect 22204 50540 22260 50542
rect 21644 49980 21700 50036
rect 21868 49922 21924 49924
rect 21868 49870 21870 49922
rect 21870 49870 21922 49922
rect 21922 49870 21924 49922
rect 21868 49868 21924 49870
rect 21756 49532 21812 49588
rect 21420 46396 21476 46452
rect 21308 45724 21364 45780
rect 21532 45948 21588 46004
rect 22204 49026 22260 49028
rect 22204 48974 22206 49026
rect 22206 48974 22258 49026
rect 22258 48974 22260 49026
rect 22204 48972 22260 48974
rect 22204 47180 22260 47236
rect 21868 45778 21924 45780
rect 21868 45726 21870 45778
rect 21870 45726 21922 45778
rect 21922 45726 21924 45778
rect 21868 45724 21924 45726
rect 21196 44828 21252 44884
rect 21420 44940 21476 44996
rect 21420 44716 21476 44772
rect 21868 45052 21924 45108
rect 21532 44604 21588 44660
rect 21756 44828 21812 44884
rect 21532 44380 21588 44436
rect 21420 44044 21476 44100
rect 20972 43484 21028 43540
rect 20300 42642 20356 42644
rect 20300 42590 20302 42642
rect 20302 42590 20354 42642
rect 20354 42590 20356 42642
rect 20300 42588 20356 42590
rect 20748 43372 20804 43428
rect 20300 41970 20356 41972
rect 20300 41918 20302 41970
rect 20302 41918 20354 41970
rect 20354 41918 20356 41970
rect 20300 41916 20356 41918
rect 20076 41858 20132 41860
rect 20076 41806 20078 41858
rect 20078 41806 20130 41858
rect 20130 41806 20132 41858
rect 20076 41804 20132 41806
rect 19180 41132 19236 41188
rect 19628 41186 19684 41188
rect 19628 41134 19630 41186
rect 19630 41134 19682 41186
rect 19682 41134 19684 41186
rect 19628 41132 19684 41134
rect 19068 37324 19124 37380
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20636 41020 20692 41076
rect 20188 40348 20244 40404
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19516 38444 19572 38500
rect 19516 37378 19572 37380
rect 19516 37326 19518 37378
rect 19518 37326 19570 37378
rect 19570 37326 19572 37378
rect 19516 37324 19572 37326
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19852 37266 19908 37268
rect 19852 37214 19854 37266
rect 19854 37214 19906 37266
rect 19906 37214 19908 37266
rect 19852 37212 19908 37214
rect 19292 36428 19348 36484
rect 19180 36204 19236 36260
rect 19292 35756 19348 35812
rect 19404 36316 19460 36372
rect 19068 35586 19124 35588
rect 19068 35534 19070 35586
rect 19070 35534 19122 35586
rect 19122 35534 19124 35586
rect 19068 35532 19124 35534
rect 19964 36988 20020 37044
rect 19740 36428 19796 36484
rect 19852 36370 19908 36372
rect 19852 36318 19854 36370
rect 19854 36318 19906 36370
rect 19906 36318 19908 36370
rect 19852 36316 19908 36318
rect 20300 38444 20356 38500
rect 20300 37212 20356 37268
rect 19404 35420 19460 35476
rect 19180 35308 19236 35364
rect 18956 34914 19012 34916
rect 18956 34862 18958 34914
rect 18958 34862 19010 34914
rect 19010 34862 19012 34914
rect 18956 34860 19012 34862
rect 18732 33628 18788 33684
rect 19292 34018 19348 34020
rect 19292 33966 19294 34018
rect 19294 33966 19346 34018
rect 19346 33966 19348 34018
rect 19292 33964 19348 33966
rect 19068 33516 19124 33572
rect 18508 33292 18564 33348
rect 18732 33292 18788 33348
rect 17948 33068 18004 33124
rect 18396 33122 18452 33124
rect 18396 33070 18398 33122
rect 18398 33070 18450 33122
rect 18450 33070 18452 33122
rect 18396 33068 18452 33070
rect 19404 33122 19460 33124
rect 19404 33070 19406 33122
rect 19406 33070 19458 33122
rect 19458 33070 19460 33122
rect 19404 33068 19460 33070
rect 18396 30940 18452 30996
rect 18284 30828 18340 30884
rect 18956 32338 19012 32340
rect 18956 32286 18958 32338
rect 18958 32286 19010 32338
rect 19010 32286 19012 32338
rect 18956 32284 19012 32286
rect 18060 30044 18116 30100
rect 18172 29820 18228 29876
rect 18060 27634 18116 27636
rect 18060 27582 18062 27634
rect 18062 27582 18114 27634
rect 18114 27582 18116 27634
rect 18060 27580 18116 27582
rect 17612 27074 17668 27076
rect 17612 27022 17614 27074
rect 17614 27022 17666 27074
rect 17666 27022 17668 27074
rect 17612 27020 17668 27022
rect 17724 26908 17780 26964
rect 17836 27020 17892 27076
rect 17612 26684 17668 26740
rect 17276 24668 17332 24724
rect 17388 23436 17444 23492
rect 17164 21308 17220 21364
rect 17276 21756 17332 21812
rect 17052 20300 17108 20356
rect 17612 22540 17668 22596
rect 18620 30044 18676 30100
rect 18508 29708 18564 29764
rect 18396 29484 18452 29540
rect 19292 29932 19348 29988
rect 18956 29820 19012 29876
rect 18844 29538 18900 29540
rect 18844 29486 18846 29538
rect 18846 29486 18898 29538
rect 18898 29486 18900 29538
rect 18844 29484 18900 29486
rect 18508 28754 18564 28756
rect 18508 28702 18510 28754
rect 18510 28702 18562 28754
rect 18562 28702 18564 28754
rect 18508 28700 18564 28702
rect 19180 28642 19236 28644
rect 19180 28590 19182 28642
rect 19182 28590 19234 28642
rect 19234 28590 19236 28642
rect 19180 28588 19236 28590
rect 19404 29484 19460 29540
rect 19404 27858 19460 27860
rect 19404 27806 19406 27858
rect 19406 27806 19458 27858
rect 19458 27806 19460 27858
rect 19404 27804 19460 27806
rect 19404 27244 19460 27300
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19740 35810 19796 35812
rect 19740 35758 19742 35810
rect 19742 35758 19794 35810
rect 19794 35758 19796 35810
rect 19740 35756 19796 35758
rect 20188 34748 20244 34804
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19964 34076 20020 34132
rect 19628 33570 19684 33572
rect 19628 33518 19630 33570
rect 19630 33518 19682 33570
rect 19682 33518 19684 33570
rect 19628 33516 19684 33518
rect 19628 33180 19684 33236
rect 19852 33122 19908 33124
rect 19852 33070 19854 33122
rect 19854 33070 19906 33122
rect 19906 33070 19908 33122
rect 19852 33068 19908 33070
rect 20412 35756 20468 35812
rect 20412 35308 20468 35364
rect 20972 42588 21028 42644
rect 20972 40402 21028 40404
rect 20972 40350 20974 40402
rect 20974 40350 21026 40402
rect 21026 40350 21028 40402
rect 20972 40348 21028 40350
rect 20972 39676 21028 39732
rect 20636 39004 20692 39060
rect 20748 38274 20804 38276
rect 20748 38222 20750 38274
rect 20750 38222 20802 38274
rect 20802 38222 20804 38274
rect 20748 38220 20804 38222
rect 20860 36988 20916 37044
rect 20972 35922 21028 35924
rect 20972 35870 20974 35922
rect 20974 35870 21026 35922
rect 21026 35870 21028 35922
rect 20972 35868 21028 35870
rect 21532 41970 21588 41972
rect 21532 41918 21534 41970
rect 21534 41918 21586 41970
rect 21586 41918 21588 41970
rect 21532 41916 21588 41918
rect 21420 41804 21476 41860
rect 21756 44098 21812 44100
rect 21756 44046 21758 44098
rect 21758 44046 21810 44098
rect 21810 44046 21812 44098
rect 21756 44044 21812 44046
rect 22876 51772 22932 51828
rect 22764 51324 22820 51380
rect 22204 45164 22260 45220
rect 22204 44994 22260 44996
rect 22204 44942 22206 44994
rect 22206 44942 22258 44994
rect 22258 44942 22260 44994
rect 22204 44940 22260 44942
rect 22092 44380 22148 44436
rect 22652 47516 22708 47572
rect 22652 46562 22708 46564
rect 22652 46510 22654 46562
rect 22654 46510 22706 46562
rect 22706 46510 22708 46562
rect 22652 46508 22708 46510
rect 23436 52332 23492 52388
rect 23436 51212 23492 51268
rect 24444 58322 24500 58324
rect 24444 58270 24446 58322
rect 24446 58270 24498 58322
rect 24498 58270 24500 58322
rect 24444 58268 24500 58270
rect 24444 57874 24500 57876
rect 24444 57822 24446 57874
rect 24446 57822 24498 57874
rect 24498 57822 24500 57874
rect 24444 57820 24500 57822
rect 24108 56924 24164 56980
rect 24220 57036 24276 57092
rect 23884 51602 23940 51604
rect 23884 51550 23886 51602
rect 23886 51550 23938 51602
rect 23938 51550 23940 51602
rect 23884 51548 23940 51550
rect 23996 53676 24052 53732
rect 23436 49810 23492 49812
rect 23436 49758 23438 49810
rect 23438 49758 23490 49810
rect 23490 49758 23492 49810
rect 23436 49756 23492 49758
rect 23324 49420 23380 49476
rect 22764 46172 22820 46228
rect 22652 45948 22708 46004
rect 22988 47180 23044 47236
rect 22876 47068 22932 47124
rect 22988 46786 23044 46788
rect 22988 46734 22990 46786
rect 22990 46734 23042 46786
rect 23042 46734 23044 46786
rect 22988 46732 23044 46734
rect 23100 46620 23156 46676
rect 24108 52556 24164 52612
rect 24444 56306 24500 56308
rect 24444 56254 24446 56306
rect 24446 56254 24498 56306
rect 24498 56254 24500 56306
rect 24444 56252 24500 56254
rect 25228 60898 25284 60900
rect 25228 60846 25230 60898
rect 25230 60846 25282 60898
rect 25282 60846 25284 60898
rect 25228 60844 25284 60846
rect 24892 60732 24948 60788
rect 24892 60002 24948 60004
rect 24892 59950 24894 60002
rect 24894 59950 24946 60002
rect 24946 59950 24948 60002
rect 24892 59948 24948 59950
rect 25564 60786 25620 60788
rect 25564 60734 25566 60786
rect 25566 60734 25618 60786
rect 25618 60734 25620 60786
rect 25564 60732 25620 60734
rect 27356 67004 27412 67060
rect 27692 66892 27748 66948
rect 27356 66780 27412 66836
rect 27916 66892 27972 66948
rect 27804 64764 27860 64820
rect 26684 63756 26740 63812
rect 26572 63644 26628 63700
rect 26572 63138 26628 63140
rect 26572 63086 26574 63138
rect 26574 63086 26626 63138
rect 26626 63086 26628 63138
rect 26572 63084 26628 63086
rect 26460 61964 26516 62020
rect 27692 63644 27748 63700
rect 27020 63362 27076 63364
rect 27020 63310 27022 63362
rect 27022 63310 27074 63362
rect 27074 63310 27076 63362
rect 27020 63308 27076 63310
rect 27356 63138 27412 63140
rect 27356 63086 27358 63138
rect 27358 63086 27410 63138
rect 27410 63086 27412 63138
rect 27356 63084 27412 63086
rect 26684 62076 26740 62132
rect 27244 62130 27300 62132
rect 27244 62078 27246 62130
rect 27246 62078 27298 62130
rect 27298 62078 27300 62130
rect 27244 62076 27300 62078
rect 26796 61964 26852 62020
rect 26460 60002 26516 60004
rect 26460 59950 26462 60002
rect 26462 59950 26514 60002
rect 26514 59950 26516 60002
rect 26460 59948 26516 59950
rect 25564 59500 25620 59556
rect 25004 58210 25060 58212
rect 25004 58158 25006 58210
rect 25006 58158 25058 58210
rect 25058 58158 25060 58210
rect 25004 58156 25060 58158
rect 25228 58044 25284 58100
rect 25564 58492 25620 58548
rect 25900 58492 25956 58548
rect 26124 59052 26180 59108
rect 25676 58380 25732 58436
rect 25788 58268 25844 58324
rect 26348 58604 26404 58660
rect 26348 58156 26404 58212
rect 25564 58044 25620 58100
rect 24892 55356 24948 55412
rect 24668 55244 24724 55300
rect 24444 54124 24500 54180
rect 24780 54012 24836 54068
rect 24556 53058 24612 53060
rect 24556 53006 24558 53058
rect 24558 53006 24610 53058
rect 24610 53006 24612 53058
rect 24556 53004 24612 53006
rect 23996 49644 24052 49700
rect 24444 52668 24500 52724
rect 23660 49420 23716 49476
rect 23660 48242 23716 48244
rect 23660 48190 23662 48242
rect 23662 48190 23714 48242
rect 23714 48190 23716 48242
rect 23660 48188 23716 48190
rect 23548 48076 23604 48132
rect 23884 47516 23940 47572
rect 23436 47404 23492 47460
rect 23324 47234 23380 47236
rect 23324 47182 23326 47234
rect 23326 47182 23378 47234
rect 23378 47182 23380 47234
rect 23324 47180 23380 47182
rect 23996 47180 24052 47236
rect 22876 45724 22932 45780
rect 22428 44604 22484 44660
rect 22652 45052 22708 45108
rect 22428 44210 22484 44212
rect 22428 44158 22430 44210
rect 22430 44158 22482 44210
rect 22482 44158 22484 44210
rect 22428 44156 22484 44158
rect 22204 44044 22260 44100
rect 21980 43932 22036 43988
rect 22092 42924 22148 42980
rect 21980 41916 22036 41972
rect 21868 41692 21924 41748
rect 21756 41132 21812 41188
rect 21644 41020 21700 41076
rect 21532 40514 21588 40516
rect 21532 40462 21534 40514
rect 21534 40462 21586 40514
rect 21586 40462 21588 40514
rect 21532 40460 21588 40462
rect 21420 40348 21476 40404
rect 21532 39900 21588 39956
rect 21308 39058 21364 39060
rect 21308 39006 21310 39058
rect 21310 39006 21362 39058
rect 21362 39006 21364 39058
rect 21308 39004 21364 39006
rect 21420 36428 21476 36484
rect 20636 35532 20692 35588
rect 21308 35586 21364 35588
rect 21308 35534 21310 35586
rect 21310 35534 21362 35586
rect 21362 35534 21364 35586
rect 21308 35532 21364 35534
rect 21420 35420 21476 35476
rect 21196 35308 21252 35364
rect 21308 34802 21364 34804
rect 21308 34750 21310 34802
rect 21310 34750 21362 34802
rect 21362 34750 21364 34802
rect 21308 34748 21364 34750
rect 21420 34354 21476 34356
rect 21420 34302 21422 34354
rect 21422 34302 21474 34354
rect 21474 34302 21476 34354
rect 21420 34300 21476 34302
rect 20524 33180 20580 33236
rect 21084 33964 21140 34020
rect 20300 33068 20356 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19964 32674 20020 32676
rect 19964 32622 19966 32674
rect 19966 32622 20018 32674
rect 20018 32622 20020 32674
rect 19964 32620 20020 32622
rect 20412 32674 20468 32676
rect 20412 32622 20414 32674
rect 20414 32622 20466 32674
rect 20466 32622 20468 32674
rect 20412 32620 20468 32622
rect 20972 32620 21028 32676
rect 20748 32508 20804 32564
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20076 30994 20132 30996
rect 20076 30942 20078 30994
rect 20078 30942 20130 30994
rect 20130 30942 20132 30994
rect 20076 30940 20132 30942
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20188 29596 20244 29652
rect 19852 28700 19908 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18284 26684 18340 26740
rect 18508 26796 18564 26852
rect 18284 26124 18340 26180
rect 20524 30882 20580 30884
rect 20524 30830 20526 30882
rect 20526 30830 20578 30882
rect 20578 30830 20580 30882
rect 20524 30828 20580 30830
rect 20748 30156 20804 30212
rect 20636 29650 20692 29652
rect 20636 29598 20638 29650
rect 20638 29598 20690 29650
rect 20690 29598 20692 29650
rect 20636 29596 20692 29598
rect 20524 28028 20580 28084
rect 20524 27746 20580 27748
rect 20524 27694 20526 27746
rect 20526 27694 20578 27746
rect 20578 27694 20580 27746
rect 20524 27692 20580 27694
rect 20412 27244 20468 27300
rect 20636 27244 20692 27300
rect 20748 27074 20804 27076
rect 20748 27022 20750 27074
rect 20750 27022 20802 27074
rect 20802 27022 20804 27074
rect 20748 27020 20804 27022
rect 18284 25506 18340 25508
rect 18284 25454 18286 25506
rect 18286 25454 18338 25506
rect 18338 25454 18340 25506
rect 18284 25452 18340 25454
rect 18060 24722 18116 24724
rect 18060 24670 18062 24722
rect 18062 24670 18114 24722
rect 18114 24670 18116 24722
rect 18060 24668 18116 24670
rect 17948 21756 18004 21812
rect 17612 21586 17668 21588
rect 17612 21534 17614 21586
rect 17614 21534 17666 21586
rect 17666 21534 17668 21586
rect 17612 21532 17668 21534
rect 17724 21362 17780 21364
rect 17724 21310 17726 21362
rect 17726 21310 17778 21362
rect 17778 21310 17780 21362
rect 17724 21308 17780 21310
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18508 25228 18564 25284
rect 18732 25788 18788 25844
rect 18508 23772 18564 23828
rect 18172 22092 18228 22148
rect 18284 21756 18340 21812
rect 18732 25564 18788 25620
rect 18732 23436 18788 23492
rect 18956 25116 19012 25172
rect 20076 25228 20132 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19964 24780 20020 24836
rect 19292 23660 19348 23716
rect 20300 24722 20356 24724
rect 20300 24670 20302 24722
rect 20302 24670 20354 24722
rect 20354 24670 20356 24722
rect 20300 24668 20356 24670
rect 20188 23826 20244 23828
rect 20188 23774 20190 23826
rect 20190 23774 20242 23826
rect 20242 23774 20244 23826
rect 20188 23772 20244 23774
rect 19852 23660 19908 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19404 22652 19460 22708
rect 20188 22652 20244 22708
rect 19740 22482 19796 22484
rect 19740 22430 19742 22482
rect 19742 22430 19794 22482
rect 19794 22430 19796 22482
rect 19740 22428 19796 22430
rect 18732 22204 18788 22260
rect 18060 21532 18116 21588
rect 17948 21196 18004 21252
rect 17836 20860 17892 20916
rect 17276 20412 17332 20468
rect 17724 20748 17780 20804
rect 17164 20076 17220 20132
rect 17948 20130 18004 20132
rect 17948 20078 17950 20130
rect 17950 20078 18002 20130
rect 18002 20078 18004 20130
rect 17948 20076 18004 20078
rect 17276 20018 17332 20020
rect 17276 19966 17278 20018
rect 17278 19966 17330 20018
rect 17330 19966 17332 20018
rect 17276 19964 17332 19966
rect 17164 18508 17220 18564
rect 18844 21868 18900 21924
rect 20076 22092 20132 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20748 25564 20804 25620
rect 20636 25452 20692 25508
rect 22316 41916 22372 41972
rect 23548 45836 23604 45892
rect 23436 45778 23492 45780
rect 23436 45726 23438 45778
rect 23438 45726 23490 45778
rect 23490 45726 23492 45778
rect 23436 45724 23492 45726
rect 23324 45276 23380 45332
rect 23772 46732 23828 46788
rect 23100 44546 23156 44548
rect 23100 44494 23102 44546
rect 23102 44494 23154 44546
rect 23154 44494 23156 44546
rect 23100 44492 23156 44494
rect 22988 44098 23044 44100
rect 22988 44046 22990 44098
rect 22990 44046 23042 44098
rect 23042 44046 23044 44098
rect 22988 44044 23044 44046
rect 22764 43932 22820 43988
rect 22652 41916 22708 41972
rect 22764 43596 22820 43652
rect 22092 41580 22148 41636
rect 21980 41132 22036 41188
rect 21868 36988 21924 37044
rect 21644 35644 21700 35700
rect 21756 35420 21812 35476
rect 21308 33346 21364 33348
rect 21308 33294 21310 33346
rect 21310 33294 21362 33346
rect 21362 33294 21364 33346
rect 21308 33292 21364 33294
rect 21532 33234 21588 33236
rect 21532 33182 21534 33234
rect 21534 33182 21586 33234
rect 21586 33182 21588 33234
rect 21532 33180 21588 33182
rect 21308 33068 21364 33124
rect 21196 30156 21252 30212
rect 21084 28700 21140 28756
rect 21196 25282 21252 25284
rect 21196 25230 21198 25282
rect 21198 25230 21250 25282
rect 21250 25230 21252 25282
rect 21196 25228 21252 25230
rect 23660 44940 23716 44996
rect 23548 44434 23604 44436
rect 23548 44382 23550 44434
rect 23550 44382 23602 44434
rect 23602 44382 23604 44434
rect 23548 44380 23604 44382
rect 23324 43932 23380 43988
rect 23548 44044 23604 44100
rect 23884 45890 23940 45892
rect 23884 45838 23886 45890
rect 23886 45838 23938 45890
rect 23938 45838 23940 45890
rect 23884 45836 23940 45838
rect 23996 44380 24052 44436
rect 23884 44156 23940 44212
rect 23772 43820 23828 43876
rect 25228 56924 25284 56980
rect 25340 56364 25396 56420
rect 25676 56812 25732 56868
rect 25452 55298 25508 55300
rect 25452 55246 25454 55298
rect 25454 55246 25506 55298
rect 25506 55246 25508 55298
rect 25452 55244 25508 55246
rect 25564 55132 25620 55188
rect 25340 55020 25396 55076
rect 26124 56642 26180 56644
rect 26124 56590 26126 56642
rect 26126 56590 26178 56642
rect 26178 56590 26180 56642
rect 26124 56588 26180 56590
rect 26124 56364 26180 56420
rect 26460 56812 26516 56868
rect 26460 56588 26516 56644
rect 26124 55970 26180 55972
rect 26124 55918 26126 55970
rect 26126 55918 26178 55970
rect 26178 55918 26180 55970
rect 26124 55916 26180 55918
rect 26124 55132 26180 55188
rect 26124 54572 26180 54628
rect 25788 54514 25844 54516
rect 25788 54462 25790 54514
rect 25790 54462 25842 54514
rect 25842 54462 25844 54514
rect 25788 54460 25844 54462
rect 26236 54460 26292 54516
rect 26012 54236 26068 54292
rect 25676 53676 25732 53732
rect 25452 53564 25508 53620
rect 25340 53506 25396 53508
rect 25340 53454 25342 53506
rect 25342 53454 25394 53506
rect 25394 53454 25396 53506
rect 25340 53452 25396 53454
rect 24668 52108 24724 52164
rect 24444 51996 24500 52052
rect 24220 51602 24276 51604
rect 24220 51550 24222 51602
rect 24222 51550 24274 51602
rect 24274 51550 24276 51602
rect 24220 51548 24276 51550
rect 24332 48860 24388 48916
rect 24668 49698 24724 49700
rect 24668 49646 24670 49698
rect 24670 49646 24722 49698
rect 24722 49646 24724 49698
rect 24668 49644 24724 49646
rect 24668 49084 24724 49140
rect 24556 48076 24612 48132
rect 24556 47516 24612 47572
rect 24220 46786 24276 46788
rect 24220 46734 24222 46786
rect 24222 46734 24274 46786
rect 24274 46734 24276 46786
rect 24220 46732 24276 46734
rect 24556 46674 24612 46676
rect 24556 46622 24558 46674
rect 24558 46622 24610 46674
rect 24610 46622 24612 46674
rect 24556 46620 24612 46622
rect 24332 46060 24388 46116
rect 24444 45890 24500 45892
rect 24444 45838 24446 45890
rect 24446 45838 24498 45890
rect 24498 45838 24500 45890
rect 24444 45836 24500 45838
rect 24444 45164 24500 45220
rect 24108 44044 24164 44100
rect 24108 43820 24164 43876
rect 24220 43596 24276 43652
rect 22988 41916 23044 41972
rect 22764 41692 22820 41748
rect 22428 41074 22484 41076
rect 22428 41022 22430 41074
rect 22430 41022 22482 41074
rect 22482 41022 22484 41074
rect 22428 41020 22484 41022
rect 23436 41132 23492 41188
rect 22876 40962 22932 40964
rect 22876 40910 22878 40962
rect 22878 40910 22930 40962
rect 22930 40910 22932 40962
rect 22876 40908 22932 40910
rect 22428 40796 22484 40852
rect 22652 40402 22708 40404
rect 22652 40350 22654 40402
rect 22654 40350 22706 40402
rect 22706 40350 22708 40402
rect 22652 40348 22708 40350
rect 22988 40514 23044 40516
rect 22988 40462 22990 40514
rect 22990 40462 23042 40514
rect 23042 40462 23044 40514
rect 22988 40460 23044 40462
rect 23324 40514 23380 40516
rect 23324 40462 23326 40514
rect 23326 40462 23378 40514
rect 23378 40462 23380 40514
rect 23324 40460 23380 40462
rect 23660 41692 23716 41748
rect 24332 41916 24388 41972
rect 24444 42924 24500 42980
rect 24220 41804 24276 41860
rect 23772 41244 23828 41300
rect 23660 40908 23716 40964
rect 23884 41020 23940 41076
rect 23548 40796 23604 40852
rect 23660 40178 23716 40180
rect 23660 40126 23662 40178
rect 23662 40126 23714 40178
rect 23714 40126 23716 40178
rect 23660 40124 23716 40126
rect 22316 39058 22372 39060
rect 22316 39006 22318 39058
rect 22318 39006 22370 39058
rect 22370 39006 22372 39058
rect 22316 39004 22372 39006
rect 22764 38780 22820 38836
rect 23212 39618 23268 39620
rect 23212 39566 23214 39618
rect 23214 39566 23266 39618
rect 23266 39566 23268 39618
rect 23212 39564 23268 39566
rect 22092 35308 22148 35364
rect 21980 34914 22036 34916
rect 21980 34862 21982 34914
rect 21982 34862 22034 34914
rect 22034 34862 22036 34914
rect 21980 34860 22036 34862
rect 21868 34748 21924 34804
rect 22316 36594 22372 36596
rect 22316 36542 22318 36594
rect 22318 36542 22370 36594
rect 22370 36542 22372 36594
rect 22316 36540 22372 36542
rect 22204 34300 22260 34356
rect 21980 33234 22036 33236
rect 21980 33182 21982 33234
rect 21982 33182 22034 33234
rect 22034 33182 22036 33234
rect 21980 33180 22036 33182
rect 21868 32562 21924 32564
rect 21868 32510 21870 32562
rect 21870 32510 21922 32562
rect 21922 32510 21924 32562
rect 21868 32508 21924 32510
rect 21756 31388 21812 31444
rect 22316 31500 22372 31556
rect 21868 31276 21924 31332
rect 21644 29596 21700 29652
rect 21868 29986 21924 29988
rect 21868 29934 21870 29986
rect 21870 29934 21922 29986
rect 21922 29934 21924 29986
rect 21868 29932 21924 29934
rect 21532 28642 21588 28644
rect 21532 28590 21534 28642
rect 21534 28590 21586 28642
rect 21586 28590 21588 28642
rect 21532 28588 21588 28590
rect 21644 28476 21700 28532
rect 21532 27970 21588 27972
rect 21532 27918 21534 27970
rect 21534 27918 21586 27970
rect 21586 27918 21588 27970
rect 21532 27916 21588 27918
rect 22652 37378 22708 37380
rect 22652 37326 22654 37378
rect 22654 37326 22706 37378
rect 22706 37326 22708 37378
rect 22652 37324 22708 37326
rect 22652 36652 22708 36708
rect 22764 35868 22820 35924
rect 23548 39618 23604 39620
rect 23548 39566 23550 39618
rect 23550 39566 23602 39618
rect 23602 39566 23604 39618
rect 23548 39564 23604 39566
rect 23548 38834 23604 38836
rect 23548 38782 23550 38834
rect 23550 38782 23602 38834
rect 23602 38782 23604 38834
rect 23548 38780 23604 38782
rect 23100 36594 23156 36596
rect 23100 36542 23102 36594
rect 23102 36542 23154 36594
rect 23154 36542 23156 36594
rect 23100 36540 23156 36542
rect 22988 34860 23044 34916
rect 23100 35308 23156 35364
rect 22764 32562 22820 32564
rect 22764 32510 22766 32562
rect 22766 32510 22818 32562
rect 22818 32510 22820 32562
rect 22764 32508 22820 32510
rect 24668 45388 24724 45444
rect 26236 53506 26292 53508
rect 26236 53454 26238 53506
rect 26238 53454 26290 53506
rect 26290 53454 26292 53506
rect 26236 53452 26292 53454
rect 25900 52780 25956 52836
rect 25004 51884 25060 51940
rect 24892 51324 24948 51380
rect 25340 51996 25396 52052
rect 26236 52722 26292 52724
rect 26236 52670 26238 52722
rect 26238 52670 26290 52722
rect 26290 52670 26292 52722
rect 26236 52668 26292 52670
rect 25452 51548 25508 51604
rect 25788 51884 25844 51940
rect 25788 50204 25844 50260
rect 25900 50428 25956 50484
rect 25340 49980 25396 50036
rect 26236 51884 26292 51940
rect 26236 50764 26292 50820
rect 25340 49644 25396 49700
rect 26124 49868 26180 49924
rect 26012 49308 26068 49364
rect 26012 48972 26068 49028
rect 27132 61682 27188 61684
rect 27132 61630 27134 61682
rect 27134 61630 27186 61682
rect 27186 61630 27188 61682
rect 27132 61628 27188 61630
rect 26908 58658 26964 58660
rect 26908 58606 26910 58658
rect 26910 58606 26962 58658
rect 26962 58606 26964 58658
rect 26908 58604 26964 58606
rect 27020 58380 27076 58436
rect 26908 57372 26964 57428
rect 27804 60620 27860 60676
rect 27804 59106 27860 59108
rect 27804 59054 27806 59106
rect 27806 59054 27858 59106
rect 27858 59054 27860 59106
rect 27804 59052 27860 59054
rect 28028 63084 28084 63140
rect 28028 62466 28084 62468
rect 28028 62414 28030 62466
rect 28030 62414 28082 62466
rect 28082 62414 28084 62466
rect 28028 62412 28084 62414
rect 29148 76412 29204 76468
rect 31164 76636 31220 76692
rect 32620 76690 32676 76692
rect 32620 76638 32622 76690
rect 32622 76638 32674 76690
rect 32674 76638 32676 76690
rect 32620 76636 32676 76638
rect 31164 76466 31220 76468
rect 31164 76414 31166 76466
rect 31166 76414 31218 76466
rect 31218 76414 31220 76466
rect 31164 76412 31220 76414
rect 32396 76412 32452 76468
rect 29260 75682 29316 75684
rect 29260 75630 29262 75682
rect 29262 75630 29314 75682
rect 29314 75630 29316 75682
rect 29260 75628 29316 75630
rect 29596 75628 29652 75684
rect 31500 75682 31556 75684
rect 31500 75630 31502 75682
rect 31502 75630 31554 75682
rect 31554 75630 31556 75682
rect 31500 75628 31556 75630
rect 31948 75682 32004 75684
rect 31948 75630 31950 75682
rect 31950 75630 32002 75682
rect 32002 75630 32004 75682
rect 31948 75628 32004 75630
rect 29596 74844 29652 74900
rect 31276 74786 31332 74788
rect 31276 74734 31278 74786
rect 31278 74734 31330 74786
rect 31330 74734 31332 74786
rect 31276 74732 31332 74734
rect 36876 76636 36932 76692
rect 35084 76524 35140 76580
rect 33404 76466 33460 76468
rect 33404 76414 33406 76466
rect 33406 76414 33458 76466
rect 33458 76414 33460 76466
rect 33404 76412 33460 76414
rect 34748 76412 34804 76468
rect 28364 72044 28420 72100
rect 33964 73612 34020 73668
rect 36092 76578 36148 76580
rect 36092 76526 36094 76578
rect 36094 76526 36146 76578
rect 36146 76526 36148 76578
rect 36092 76524 36148 76526
rect 37548 76690 37604 76692
rect 37548 76638 37550 76690
rect 37550 76638 37602 76690
rect 37602 76638 37604 76690
rect 37548 76636 37604 76638
rect 42364 76636 42420 76692
rect 40124 76524 40180 76580
rect 40796 76524 40852 76580
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 38332 75852 38388 75908
rect 41468 76578 41524 76580
rect 41468 76526 41470 76578
rect 41470 76526 41522 76578
rect 41522 76526 41524 76578
rect 41468 76524 41524 76526
rect 42924 76690 42980 76692
rect 42924 76638 42926 76690
rect 42926 76638 42978 76690
rect 42978 76638 42980 76690
rect 42924 76636 42980 76638
rect 43708 76466 43764 76468
rect 43708 76414 43710 76466
rect 43710 76414 43762 76466
rect 43762 76414 43764 76466
rect 43708 76412 43764 76414
rect 40012 75740 40068 75796
rect 36540 73164 36596 73220
rect 40348 73948 40404 74004
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 34300 72604 34356 72660
rect 31164 71986 31220 71988
rect 31164 71934 31166 71986
rect 31166 71934 31218 71986
rect 31218 71934 31220 71986
rect 31164 71932 31220 71934
rect 28476 71820 28532 71876
rect 29820 71874 29876 71876
rect 29820 71822 29822 71874
rect 29822 71822 29874 71874
rect 29874 71822 29876 71874
rect 29820 71820 29876 71822
rect 28252 70476 28308 70532
rect 29148 70476 29204 70532
rect 29036 70364 29092 70420
rect 28364 67058 28420 67060
rect 28364 67006 28366 67058
rect 28366 67006 28418 67058
rect 28418 67006 28420 67058
rect 28364 67004 28420 67006
rect 29260 67116 29316 67172
rect 28588 66780 28644 66836
rect 29148 65996 29204 66052
rect 29596 70588 29652 70644
rect 30492 71874 30548 71876
rect 30492 71822 30494 71874
rect 30494 71822 30546 71874
rect 30546 71822 30548 71874
rect 30492 71820 30548 71822
rect 31948 71986 32004 71988
rect 31948 71934 31950 71986
rect 31950 71934 32002 71986
rect 32002 71934 32004 71986
rect 31948 71932 32004 71934
rect 29932 70978 29988 70980
rect 29932 70926 29934 70978
rect 29934 70926 29986 70978
rect 29986 70926 29988 70978
rect 29932 70924 29988 70926
rect 33852 72268 33908 72324
rect 30268 70588 30324 70644
rect 30492 70924 30548 70980
rect 30940 70812 30996 70868
rect 29820 69804 29876 69860
rect 29820 67842 29876 67844
rect 29820 67790 29822 67842
rect 29822 67790 29874 67842
rect 29874 67790 29876 67842
rect 29820 67788 29876 67790
rect 29596 67116 29652 67172
rect 29484 67004 29540 67060
rect 29484 66274 29540 66276
rect 29484 66222 29486 66274
rect 29486 66222 29538 66274
rect 29538 66222 29540 66274
rect 29484 66220 29540 66222
rect 29596 66780 29652 66836
rect 29820 66220 29876 66276
rect 28924 62972 28980 63028
rect 27916 57036 27972 57092
rect 27244 55132 27300 55188
rect 27580 56588 27636 56644
rect 28924 60674 28980 60676
rect 28924 60622 28926 60674
rect 28926 60622 28978 60674
rect 28978 60622 28980 60674
rect 28924 60620 28980 60622
rect 28140 58492 28196 58548
rect 28364 57596 28420 57652
rect 28140 57372 28196 57428
rect 28252 56866 28308 56868
rect 28252 56814 28254 56866
rect 28254 56814 28306 56866
rect 28306 56814 28308 56866
rect 28252 56812 28308 56814
rect 28588 58210 28644 58212
rect 28588 58158 28590 58210
rect 28590 58158 28642 58210
rect 28642 58158 28644 58210
rect 28588 58156 28644 58158
rect 27132 54626 27188 54628
rect 27132 54574 27134 54626
rect 27134 54574 27186 54626
rect 27186 54574 27188 54626
rect 27132 54572 27188 54574
rect 26572 54514 26628 54516
rect 26572 54462 26574 54514
rect 26574 54462 26626 54514
rect 26626 54462 26628 54514
rect 26572 54460 26628 54462
rect 26796 54460 26852 54516
rect 26908 54514 26964 54516
rect 26908 54462 26910 54514
rect 26910 54462 26962 54514
rect 26962 54462 26964 54514
rect 26908 54460 26964 54462
rect 26796 54012 26852 54068
rect 27244 54124 27300 54180
rect 27580 55356 27636 55412
rect 27580 54460 27636 54516
rect 27580 54290 27636 54292
rect 27580 54238 27582 54290
rect 27582 54238 27634 54290
rect 27634 54238 27636 54290
rect 27580 54236 27636 54238
rect 27468 54124 27524 54180
rect 27132 53676 27188 53732
rect 26796 53564 26852 53620
rect 26684 52162 26740 52164
rect 26684 52110 26686 52162
rect 26686 52110 26738 52162
rect 26738 52110 26740 52162
rect 26684 52108 26740 52110
rect 26796 51772 26852 51828
rect 27020 51660 27076 51716
rect 26796 50876 26852 50932
rect 26684 50652 26740 50708
rect 26572 49922 26628 49924
rect 26572 49870 26574 49922
rect 26574 49870 26626 49922
rect 26626 49870 26628 49922
rect 26572 49868 26628 49870
rect 26460 49084 26516 49140
rect 25116 47516 25172 47572
rect 24892 46956 24948 47012
rect 25228 47404 25284 47460
rect 25788 48076 25844 48132
rect 25676 47570 25732 47572
rect 25676 47518 25678 47570
rect 25678 47518 25730 47570
rect 25730 47518 25732 47570
rect 25676 47516 25732 47518
rect 26236 47516 26292 47572
rect 26124 47234 26180 47236
rect 26124 47182 26126 47234
rect 26126 47182 26178 47234
rect 26178 47182 26180 47234
rect 26124 47180 26180 47182
rect 25116 46674 25172 46676
rect 25116 46622 25118 46674
rect 25118 46622 25170 46674
rect 25170 46622 25172 46674
rect 25116 46620 25172 46622
rect 25340 46562 25396 46564
rect 25340 46510 25342 46562
rect 25342 46510 25394 46562
rect 25394 46510 25396 46562
rect 25340 46508 25396 46510
rect 25564 46396 25620 46452
rect 24892 46060 24948 46116
rect 25676 45836 25732 45892
rect 24668 44268 24724 44324
rect 24892 44322 24948 44324
rect 24892 44270 24894 44322
rect 24894 44270 24946 44322
rect 24946 44270 24948 44322
rect 24892 44268 24948 44270
rect 24556 42364 24612 42420
rect 24668 43708 24724 43764
rect 25452 45276 25508 45332
rect 25228 45164 25284 45220
rect 25564 44940 25620 44996
rect 25116 44546 25172 44548
rect 25116 44494 25118 44546
rect 25118 44494 25170 44546
rect 25170 44494 25172 44546
rect 25116 44492 25172 44494
rect 25900 45218 25956 45220
rect 25900 45166 25902 45218
rect 25902 45166 25954 45218
rect 25954 45166 25956 45218
rect 25900 45164 25956 45166
rect 25788 45106 25844 45108
rect 25788 45054 25790 45106
rect 25790 45054 25842 45106
rect 25842 45054 25844 45106
rect 25788 45052 25844 45054
rect 26236 46450 26292 46452
rect 26236 46398 26238 46450
rect 26238 46398 26290 46450
rect 26290 46398 26292 46450
rect 26236 46396 26292 46398
rect 26572 47570 26628 47572
rect 26572 47518 26574 47570
rect 26574 47518 26626 47570
rect 26626 47518 26628 47570
rect 26572 47516 26628 47518
rect 27020 50428 27076 50484
rect 27132 51436 27188 51492
rect 27580 53618 27636 53620
rect 27580 53566 27582 53618
rect 27582 53566 27634 53618
rect 27634 53566 27636 53618
rect 27580 53564 27636 53566
rect 27468 53228 27524 53284
rect 27468 50540 27524 50596
rect 27132 49810 27188 49812
rect 27132 49758 27134 49810
rect 27134 49758 27186 49810
rect 27186 49758 27188 49810
rect 27132 49756 27188 49758
rect 27132 49308 27188 49364
rect 27356 49084 27412 49140
rect 27020 48972 27076 49028
rect 26684 46844 26740 46900
rect 26012 44940 26068 44996
rect 25340 43708 25396 43764
rect 25116 43596 25172 43652
rect 25564 43538 25620 43540
rect 25564 43486 25566 43538
rect 25566 43486 25618 43538
rect 25618 43486 25620 43538
rect 25564 43484 25620 43486
rect 25340 43426 25396 43428
rect 25340 43374 25342 43426
rect 25342 43374 25394 43426
rect 25394 43374 25396 43426
rect 25340 43372 25396 43374
rect 24892 42476 24948 42532
rect 25116 41970 25172 41972
rect 25116 41918 25118 41970
rect 25118 41918 25170 41970
rect 25170 41918 25172 41970
rect 25116 41916 25172 41918
rect 24668 41858 24724 41860
rect 24668 41806 24670 41858
rect 24670 41806 24722 41858
rect 24722 41806 24724 41858
rect 24668 41804 24724 41806
rect 24556 40962 24612 40964
rect 24556 40910 24558 40962
rect 24558 40910 24610 40962
rect 24610 40910 24612 40962
rect 24556 40908 24612 40910
rect 24444 39564 24500 39620
rect 24556 40684 24612 40740
rect 24780 41356 24836 41412
rect 25340 41858 25396 41860
rect 25340 41806 25342 41858
rect 25342 41806 25394 41858
rect 25394 41806 25396 41858
rect 25340 41804 25396 41806
rect 25452 41356 25508 41412
rect 25340 40348 25396 40404
rect 25116 40124 25172 40180
rect 24332 38892 24388 38948
rect 23996 38332 24052 38388
rect 23884 36764 23940 36820
rect 23772 36540 23828 36596
rect 23436 36370 23492 36372
rect 23436 36318 23438 36370
rect 23438 36318 23490 36370
rect 23490 36318 23492 36370
rect 23436 36316 23492 36318
rect 23548 35698 23604 35700
rect 23548 35646 23550 35698
rect 23550 35646 23602 35698
rect 23602 35646 23604 35698
rect 23548 35644 23604 35646
rect 23996 36652 24052 36708
rect 24780 39116 24836 39172
rect 24668 38892 24724 38948
rect 24556 38668 24612 38724
rect 23884 35644 23940 35700
rect 24220 35980 24276 36036
rect 24220 35532 24276 35588
rect 23324 32844 23380 32900
rect 22540 31724 22596 31780
rect 22540 31500 22596 31556
rect 23324 31890 23380 31892
rect 23324 31838 23326 31890
rect 23326 31838 23378 31890
rect 23378 31838 23380 31890
rect 23324 31836 23380 31838
rect 22876 31388 22932 31444
rect 22540 30940 22596 30996
rect 23212 30828 23268 30884
rect 22092 28530 22148 28532
rect 22092 28478 22094 28530
rect 22094 28478 22146 28530
rect 22146 28478 22148 28530
rect 22092 28476 22148 28478
rect 21980 27804 22036 27860
rect 21644 27132 21700 27188
rect 21868 27298 21924 27300
rect 21868 27246 21870 27298
rect 21870 27246 21922 27298
rect 21922 27246 21924 27298
rect 21868 27244 21924 27246
rect 21868 26908 21924 26964
rect 21532 25564 21588 25620
rect 21420 25394 21476 25396
rect 21420 25342 21422 25394
rect 21422 25342 21474 25394
rect 21474 25342 21476 25394
rect 21420 25340 21476 25342
rect 20860 24834 20916 24836
rect 20860 24782 20862 24834
rect 20862 24782 20914 24834
rect 20914 24782 20916 24834
rect 20860 24780 20916 24782
rect 20524 22316 20580 22372
rect 21420 23660 21476 23716
rect 21308 22316 21364 22372
rect 21084 22204 21140 22260
rect 20188 21532 20244 21588
rect 20636 21586 20692 21588
rect 20636 21534 20638 21586
rect 20638 21534 20690 21586
rect 20690 21534 20692 21586
rect 20636 21532 20692 21534
rect 19516 21308 19572 21364
rect 19292 20802 19348 20804
rect 19292 20750 19294 20802
rect 19294 20750 19346 20802
rect 19346 20750 19348 20802
rect 19292 20748 19348 20750
rect 18844 20300 18900 20356
rect 18732 19740 18788 19796
rect 17836 18396 17892 18452
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 16716 17500 16772 17556
rect 15708 16828 15764 16884
rect 16268 16828 16324 16884
rect 15708 15484 15764 15540
rect 16156 15484 16212 15540
rect 15708 14588 15764 14644
rect 18732 16882 18788 16884
rect 18732 16830 18734 16882
rect 18734 16830 18786 16882
rect 18786 16830 18788 16882
rect 18732 16828 18788 16830
rect 18732 16604 18788 16660
rect 15372 14418 15428 14420
rect 15372 14366 15374 14418
rect 15374 14366 15426 14418
rect 15426 14366 15428 14418
rect 15372 14364 15428 14366
rect 16716 14588 16772 14644
rect 16604 14418 16660 14420
rect 16604 14366 16606 14418
rect 16606 14366 16658 14418
rect 16658 14366 16660 14418
rect 16604 14364 16660 14366
rect 15484 13804 15540 13860
rect 15372 12850 15428 12852
rect 15372 12798 15374 12850
rect 15374 12798 15426 12850
rect 15426 12798 15428 12850
rect 15372 12796 15428 12798
rect 15372 12348 15428 12404
rect 15148 12178 15204 12180
rect 15148 12126 15150 12178
rect 15150 12126 15202 12178
rect 15202 12126 15204 12178
rect 15148 12124 15204 12126
rect 15596 13244 15652 13300
rect 15036 11788 15092 11844
rect 17836 14530 17892 14532
rect 17836 14478 17838 14530
rect 17838 14478 17890 14530
rect 17890 14478 17892 14530
rect 17836 14476 17892 14478
rect 16716 13916 16772 13972
rect 17052 14364 17108 14420
rect 15932 13634 15988 13636
rect 15932 13582 15934 13634
rect 15934 13582 15986 13634
rect 15986 13582 15988 13634
rect 15932 13580 15988 13582
rect 15820 13356 15876 13412
rect 15932 13244 15988 13300
rect 15932 13074 15988 13076
rect 15932 13022 15934 13074
rect 15934 13022 15986 13074
rect 15986 13022 15988 13074
rect 15932 13020 15988 13022
rect 17388 14306 17444 14308
rect 17388 14254 17390 14306
rect 17390 14254 17442 14306
rect 17442 14254 17444 14306
rect 17388 14252 17444 14254
rect 17612 13468 17668 13524
rect 15820 12124 15876 12180
rect 16604 12402 16660 12404
rect 16604 12350 16606 12402
rect 16606 12350 16658 12402
rect 16658 12350 16660 12402
rect 16604 12348 16660 12350
rect 15596 11788 15652 11844
rect 14364 9548 14420 9604
rect 14924 9154 14980 9156
rect 14924 9102 14926 9154
rect 14926 9102 14978 9154
rect 14978 9102 14980 9154
rect 14924 9100 14980 9102
rect 15708 9996 15764 10052
rect 15596 9826 15652 9828
rect 15596 9774 15598 9826
rect 15598 9774 15650 9826
rect 15650 9774 15652 9826
rect 15596 9772 15652 9774
rect 15820 9884 15876 9940
rect 15484 8316 15540 8372
rect 15708 8258 15764 8260
rect 15708 8206 15710 8258
rect 15710 8206 15762 8258
rect 15762 8206 15764 8258
rect 15708 8204 15764 8206
rect 13468 5906 13524 5908
rect 13468 5854 13470 5906
rect 13470 5854 13522 5906
rect 13522 5854 13524 5906
rect 13468 5852 13524 5854
rect 14364 5852 14420 5908
rect 14588 5682 14644 5684
rect 14588 5630 14590 5682
rect 14590 5630 14642 5682
rect 14642 5630 14644 5682
rect 14588 5628 14644 5630
rect 15036 5740 15092 5796
rect 15708 5740 15764 5796
rect 16604 9996 16660 10052
rect 16268 9938 16324 9940
rect 16268 9886 16270 9938
rect 16270 9886 16322 9938
rect 16322 9886 16324 9938
rect 16268 9884 16324 9886
rect 17164 9938 17220 9940
rect 17164 9886 17166 9938
rect 17166 9886 17218 9938
rect 17218 9886 17220 9938
rect 17164 9884 17220 9886
rect 16492 8316 16548 8372
rect 16604 8204 16660 8260
rect 17388 8146 17444 8148
rect 17388 8094 17390 8146
rect 17390 8094 17442 8146
rect 17442 8094 17444 8146
rect 17388 8092 17444 8094
rect 16268 5906 16324 5908
rect 16268 5854 16270 5906
rect 16270 5854 16322 5906
rect 16322 5854 16324 5906
rect 16268 5852 16324 5854
rect 18732 13970 18788 13972
rect 18732 13918 18734 13970
rect 18734 13918 18786 13970
rect 18786 13918 18788 13970
rect 18732 13916 18788 13918
rect 18620 12684 18676 12740
rect 18172 11116 18228 11172
rect 17724 9548 17780 9604
rect 18396 9548 18452 9604
rect 19180 18338 19236 18340
rect 19180 18286 19182 18338
rect 19182 18286 19234 18338
rect 19234 18286 19236 18338
rect 19180 18284 19236 18286
rect 19068 17554 19124 17556
rect 19068 17502 19070 17554
rect 19070 17502 19122 17554
rect 19122 17502 19124 17554
rect 19068 17500 19124 17502
rect 19180 16044 19236 16100
rect 19292 15986 19348 15988
rect 19292 15934 19294 15986
rect 19294 15934 19346 15986
rect 19346 15934 19348 15986
rect 19292 15932 19348 15934
rect 20524 21362 20580 21364
rect 20524 21310 20526 21362
rect 20526 21310 20578 21362
rect 20578 21310 20580 21362
rect 20524 21308 20580 21310
rect 20300 21196 20356 21252
rect 20188 20636 20244 20692
rect 20076 20524 20132 20580
rect 20748 20636 20804 20692
rect 20972 21756 21028 21812
rect 20412 20524 20468 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 20018 19796 20020
rect 19740 19966 19742 20018
rect 19742 19966 19794 20018
rect 19794 19966 19796 20018
rect 19740 19964 19796 19966
rect 19628 19740 19684 19796
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20076 18338 20132 18340
rect 20076 18286 20078 18338
rect 20078 18286 20130 18338
rect 20130 18286 20132 18338
rect 20076 18284 20132 18286
rect 21532 22092 21588 22148
rect 21420 20748 21476 20804
rect 21196 20636 21252 20692
rect 21532 20130 21588 20132
rect 21532 20078 21534 20130
rect 21534 20078 21586 20130
rect 21586 20078 21588 20130
rect 21532 20076 21588 20078
rect 21868 20018 21924 20020
rect 21868 19966 21870 20018
rect 21870 19966 21922 20018
rect 21922 19966 21924 20018
rect 21868 19964 21924 19966
rect 22652 28642 22708 28644
rect 22652 28590 22654 28642
rect 22654 28590 22706 28642
rect 22706 28590 22708 28642
rect 22652 28588 22708 28590
rect 22764 27916 22820 27972
rect 22764 27186 22820 27188
rect 22764 27134 22766 27186
rect 22766 27134 22818 27186
rect 22818 27134 22820 27186
rect 22764 27132 22820 27134
rect 22764 26908 22820 26964
rect 22092 26514 22148 26516
rect 22092 26462 22094 26514
rect 22094 26462 22146 26514
rect 22146 26462 22148 26514
rect 22092 26460 22148 26462
rect 22092 22482 22148 22484
rect 22092 22430 22094 22482
rect 22094 22430 22146 22482
rect 22146 22430 22148 22482
rect 22092 22428 22148 22430
rect 22204 22370 22260 22372
rect 22204 22318 22206 22370
rect 22206 22318 22258 22370
rect 22258 22318 22260 22370
rect 22204 22316 22260 22318
rect 22204 22092 22260 22148
rect 23548 31778 23604 31780
rect 23548 31726 23550 31778
rect 23550 31726 23602 31778
rect 23602 31726 23604 31778
rect 23548 31724 23604 31726
rect 23772 31554 23828 31556
rect 23772 31502 23774 31554
rect 23774 31502 23826 31554
rect 23826 31502 23828 31554
rect 23772 31500 23828 31502
rect 23884 30828 23940 30884
rect 23996 32284 24052 32340
rect 23548 30210 23604 30212
rect 23548 30158 23550 30210
rect 23550 30158 23602 30210
rect 23602 30158 23604 30210
rect 23548 30156 23604 30158
rect 23996 30156 24052 30212
rect 24220 28754 24276 28756
rect 24220 28702 24222 28754
rect 24222 28702 24274 28754
rect 24274 28702 24276 28754
rect 24220 28700 24276 28702
rect 23436 27916 23492 27972
rect 23100 27580 23156 27636
rect 23100 26908 23156 26964
rect 23996 27634 24052 27636
rect 23996 27582 23998 27634
rect 23998 27582 24050 27634
rect 24050 27582 24052 27634
rect 23996 27580 24052 27582
rect 23772 27132 23828 27188
rect 24220 27074 24276 27076
rect 24220 27022 24222 27074
rect 24222 27022 24274 27074
rect 24274 27022 24276 27074
rect 24220 27020 24276 27022
rect 23772 26290 23828 26292
rect 23772 26238 23774 26290
rect 23774 26238 23826 26290
rect 23826 26238 23828 26290
rect 23772 26236 23828 26238
rect 24556 35980 24612 36036
rect 24556 35196 24612 35252
rect 24892 38332 24948 38388
rect 25004 38050 25060 38052
rect 25004 37998 25006 38050
rect 25006 37998 25058 38050
rect 25058 37998 25060 38050
rect 25004 37996 25060 37998
rect 24892 37826 24948 37828
rect 24892 37774 24894 37826
rect 24894 37774 24946 37826
rect 24946 37774 24948 37826
rect 24892 37772 24948 37774
rect 24892 34300 24948 34356
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 24780 31276 24836 31332
rect 24668 29650 24724 29652
rect 24668 29598 24670 29650
rect 24670 29598 24722 29650
rect 24722 29598 24724 29650
rect 24668 29596 24724 29598
rect 23436 24556 23492 24612
rect 23212 23938 23268 23940
rect 23212 23886 23214 23938
rect 23214 23886 23266 23938
rect 23266 23886 23268 23938
rect 23212 23884 23268 23886
rect 22876 23826 22932 23828
rect 22876 23774 22878 23826
rect 22878 23774 22930 23826
rect 22930 23774 22932 23826
rect 22876 23772 22932 23774
rect 22988 23548 23044 23604
rect 22092 20242 22148 20244
rect 22092 20190 22094 20242
rect 22094 20190 22146 20242
rect 22146 20190 22148 20242
rect 22092 20188 22148 20190
rect 21980 19516 22036 19572
rect 21868 18956 21924 19012
rect 20524 18284 20580 18340
rect 19964 17554 20020 17556
rect 19964 17502 19966 17554
rect 19966 17502 20018 17554
rect 20018 17502 20020 17554
rect 19964 17500 20020 17502
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20188 16210 20244 16212
rect 20188 16158 20190 16210
rect 20190 16158 20242 16210
rect 20242 16158 20244 16210
rect 20188 16156 20244 16158
rect 19964 16098 20020 16100
rect 19964 16046 19966 16098
rect 19966 16046 20018 16098
rect 20018 16046 20020 16098
rect 19964 16044 20020 16046
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20860 16210 20916 16212
rect 20860 16158 20862 16210
rect 20862 16158 20914 16210
rect 20914 16158 20916 16210
rect 20860 16156 20916 16158
rect 19628 15036 19684 15092
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19628 13916 19684 13972
rect 21420 18060 21476 18116
rect 21420 16994 21476 16996
rect 21420 16942 21422 16994
rect 21422 16942 21474 16994
rect 21474 16942 21476 16994
rect 21420 16940 21476 16942
rect 21084 16882 21140 16884
rect 21084 16830 21086 16882
rect 21086 16830 21138 16882
rect 21138 16830 21140 16882
rect 21084 16828 21140 16830
rect 22540 20188 22596 20244
rect 22316 20130 22372 20132
rect 22316 20078 22318 20130
rect 22318 20078 22370 20130
rect 22370 20078 22372 20130
rect 22316 20076 22372 20078
rect 23212 20076 23268 20132
rect 22204 19010 22260 19012
rect 22204 18958 22206 19010
rect 22206 18958 22258 19010
rect 22258 18958 22260 19010
rect 22204 18956 22260 18958
rect 22652 18284 22708 18340
rect 22204 16994 22260 16996
rect 22204 16942 22206 16994
rect 22206 16942 22258 16994
rect 22258 16942 22260 16994
rect 22204 16940 22260 16942
rect 22092 16210 22148 16212
rect 22092 16158 22094 16210
rect 22094 16158 22146 16210
rect 22146 16158 22148 16210
rect 22092 16156 22148 16158
rect 21980 16098 22036 16100
rect 21980 16046 21982 16098
rect 21982 16046 22034 16098
rect 22034 16046 22036 16098
rect 21980 16044 22036 16046
rect 21532 15538 21588 15540
rect 21532 15486 21534 15538
rect 21534 15486 21586 15538
rect 21586 15486 21588 15538
rect 21532 15484 21588 15486
rect 22316 15820 22372 15876
rect 22316 15484 22372 15540
rect 21196 15036 21252 15092
rect 20636 13746 20692 13748
rect 20636 13694 20638 13746
rect 20638 13694 20690 13746
rect 20690 13694 20692 13746
rect 20636 13692 20692 13694
rect 19292 13522 19348 13524
rect 19292 13470 19294 13522
rect 19294 13470 19346 13522
rect 19346 13470 19348 13522
rect 19292 13468 19348 13470
rect 19628 13020 19684 13076
rect 19068 12850 19124 12852
rect 19068 12798 19070 12850
rect 19070 12798 19122 12850
rect 19122 12798 19124 12850
rect 19068 12796 19124 12798
rect 20076 13074 20132 13076
rect 20076 13022 20078 13074
rect 20078 13022 20130 13074
rect 20130 13022 20132 13074
rect 20076 13020 20132 13022
rect 20412 13020 20468 13076
rect 19628 12796 19684 12852
rect 19068 11788 19124 11844
rect 18620 10610 18676 10612
rect 18620 10558 18622 10610
rect 18622 10558 18674 10610
rect 18674 10558 18676 10610
rect 18620 10556 18676 10558
rect 18956 11170 19012 11172
rect 18956 11118 18958 11170
rect 18958 11118 19010 11170
rect 19010 11118 19012 11170
rect 18956 11116 19012 11118
rect 18732 9714 18788 9716
rect 18732 9662 18734 9714
rect 18734 9662 18786 9714
rect 18786 9662 18788 9714
rect 18732 9660 18788 9662
rect 17948 8316 18004 8372
rect 17724 8258 17780 8260
rect 17724 8206 17726 8258
rect 17726 8206 17778 8258
rect 17778 8206 17780 8258
rect 17724 8204 17780 8206
rect 18620 8092 18676 8148
rect 19740 12738 19796 12740
rect 19740 12686 19742 12738
rect 19742 12686 19794 12738
rect 19794 12686 19796 12738
rect 19740 12684 19796 12686
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19628 10610 19684 10612
rect 19628 10558 19630 10610
rect 19630 10558 19682 10610
rect 19682 10558 19684 10610
rect 19628 10556 19684 10558
rect 19180 9772 19236 9828
rect 20076 10610 20132 10612
rect 20076 10558 20078 10610
rect 20078 10558 20130 10610
rect 20130 10558 20132 10610
rect 20076 10556 20132 10558
rect 20748 10556 20804 10612
rect 21084 13580 21140 13636
rect 20188 9826 20244 9828
rect 20188 9774 20190 9826
rect 20190 9774 20242 9826
rect 20242 9774 20244 9826
rect 20188 9772 20244 9774
rect 19628 9714 19684 9716
rect 19628 9662 19630 9714
rect 19630 9662 19682 9714
rect 19682 9662 19684 9714
rect 19628 9660 19684 9662
rect 21532 14530 21588 14532
rect 21532 14478 21534 14530
rect 21534 14478 21586 14530
rect 21586 14478 21588 14530
rect 21532 14476 21588 14478
rect 22540 15372 22596 15428
rect 22876 15426 22932 15428
rect 22876 15374 22878 15426
rect 22878 15374 22930 15426
rect 22930 15374 22932 15426
rect 22876 15372 22932 15374
rect 22092 14306 22148 14308
rect 22092 14254 22094 14306
rect 22094 14254 22146 14306
rect 22146 14254 22148 14306
rect 22092 14252 22148 14254
rect 22652 14418 22708 14420
rect 22652 14366 22654 14418
rect 22654 14366 22706 14418
rect 22706 14366 22708 14418
rect 22652 14364 22708 14366
rect 22204 13746 22260 13748
rect 22204 13694 22206 13746
rect 22206 13694 22258 13746
rect 22258 13694 22260 13746
rect 22204 13692 22260 13694
rect 21756 13580 21812 13636
rect 21532 10722 21588 10724
rect 21532 10670 21534 10722
rect 21534 10670 21586 10722
rect 21586 10670 21588 10722
rect 21532 10668 21588 10670
rect 21868 10556 21924 10612
rect 20860 9660 20916 9716
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 8146 19572 8148
rect 19516 8094 19518 8146
rect 19518 8094 19570 8146
rect 19570 8094 19572 8146
rect 19516 8092 19572 8094
rect 20412 8146 20468 8148
rect 20412 8094 20414 8146
rect 20414 8094 20466 8146
rect 20466 8094 20468 8146
rect 20412 8092 20468 8094
rect 20076 7980 20132 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20636 8034 20692 8036
rect 20636 7982 20638 8034
rect 20638 7982 20690 8034
rect 20690 7982 20692 8034
rect 20636 7980 20692 7982
rect 20972 7586 21028 7588
rect 20972 7534 20974 7586
rect 20974 7534 21026 7586
rect 21026 7534 21028 7586
rect 20972 7532 21028 7534
rect 16716 5852 16772 5908
rect 18396 6018 18452 6020
rect 18396 5966 18398 6018
rect 18398 5966 18450 6018
rect 18450 5966 18452 6018
rect 18396 5964 18452 5966
rect 17724 5906 17780 5908
rect 17724 5854 17726 5906
rect 17726 5854 17778 5906
rect 17778 5854 17780 5906
rect 17724 5852 17780 5854
rect 18844 6076 18900 6132
rect 17276 5628 17332 5684
rect 17948 5180 18004 5236
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19068 5852 19124 5908
rect 19180 5964 19236 6020
rect 19404 5292 19460 5348
rect 20300 6130 20356 6132
rect 20300 6078 20302 6130
rect 20302 6078 20354 6130
rect 20354 6078 20356 6130
rect 20300 6076 20356 6078
rect 19852 5852 19908 5908
rect 20860 5852 20916 5908
rect 20300 5682 20356 5684
rect 20300 5630 20302 5682
rect 20302 5630 20354 5682
rect 20354 5630 20356 5682
rect 20300 5628 20356 5630
rect 20524 5292 20580 5348
rect 20748 5122 20804 5124
rect 20748 5070 20750 5122
rect 20750 5070 20802 5122
rect 20802 5070 20804 5122
rect 20748 5068 20804 5070
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 14700 4450 14756 4452
rect 14700 4398 14702 4450
rect 14702 4398 14754 4450
rect 14754 4398 14756 4450
rect 14700 4396 14756 4398
rect 11340 4172 11396 4228
rect 8764 3388 8820 3444
rect 13468 4226 13524 4228
rect 13468 4174 13470 4226
rect 13470 4174 13522 4226
rect 13522 4174 13524 4226
rect 13468 4172 13524 4174
rect 14812 3442 14868 3444
rect 14812 3390 14814 3442
rect 14814 3390 14866 3442
rect 14866 3390 14868 3442
rect 14812 3388 14868 3390
rect 18956 4060 19012 4116
rect 15372 3442 15428 3444
rect 15372 3390 15374 3442
rect 15374 3390 15426 3442
rect 15426 3390 15428 3442
rect 15372 3388 15428 3390
rect 19404 4114 19460 4116
rect 19404 4062 19406 4114
rect 19406 4062 19458 4114
rect 19458 4062 19460 4114
rect 19404 4060 19460 4062
rect 21644 9714 21700 9716
rect 21644 9662 21646 9714
rect 21646 9662 21698 9714
rect 21698 9662 21700 9714
rect 21644 9660 21700 9662
rect 21756 8316 21812 8372
rect 22540 12684 22596 12740
rect 23100 16210 23156 16212
rect 23100 16158 23102 16210
rect 23102 16158 23154 16210
rect 23154 16158 23156 16210
rect 23100 16156 23156 16158
rect 22764 11676 22820 11732
rect 24108 24332 24164 24388
rect 23548 23772 23604 23828
rect 23996 23660 24052 23716
rect 24220 23548 24276 23604
rect 24220 20130 24276 20132
rect 24220 20078 24222 20130
rect 24222 20078 24274 20130
rect 24274 20078 24276 20130
rect 24220 20076 24276 20078
rect 23996 19346 24052 19348
rect 23996 19294 23998 19346
rect 23998 19294 24050 19346
rect 24050 19294 24052 19346
rect 23996 19292 24052 19294
rect 23436 18844 23492 18900
rect 23436 15874 23492 15876
rect 23436 15822 23438 15874
rect 23438 15822 23490 15874
rect 23490 15822 23492 15874
rect 23436 15820 23492 15822
rect 23324 15260 23380 15316
rect 24332 18396 24388 18452
rect 24444 17612 24500 17668
rect 24668 16268 24724 16324
rect 24444 15484 24500 15540
rect 24108 15314 24164 15316
rect 24108 15262 24110 15314
rect 24110 15262 24162 15314
rect 24162 15262 24164 15314
rect 24108 15260 24164 15262
rect 23548 14476 23604 14532
rect 24668 14252 24724 14308
rect 23996 13804 24052 13860
rect 23436 13692 23492 13748
rect 23436 13522 23492 13524
rect 23436 13470 23438 13522
rect 23438 13470 23490 13522
rect 23490 13470 23492 13522
rect 23436 13468 23492 13470
rect 24108 13746 24164 13748
rect 24108 13694 24110 13746
rect 24110 13694 24162 13746
rect 24162 13694 24164 13746
rect 24108 13692 24164 13694
rect 24556 13692 24612 13748
rect 23772 11788 23828 11844
rect 22764 10668 22820 10724
rect 23660 11676 23716 11732
rect 24556 11116 24612 11172
rect 24892 29596 24948 29652
rect 25004 26124 25060 26180
rect 25676 42364 25732 42420
rect 26236 45778 26292 45780
rect 26236 45726 26238 45778
rect 26238 45726 26290 45778
rect 26290 45726 26292 45778
rect 26236 45724 26292 45726
rect 27580 47292 27636 47348
rect 26684 46396 26740 46452
rect 26236 43708 26292 43764
rect 26236 42754 26292 42756
rect 26236 42702 26238 42754
rect 26238 42702 26290 42754
rect 26290 42702 26292 42754
rect 26236 42700 26292 42702
rect 25564 40460 25620 40516
rect 25788 39116 25844 39172
rect 25788 38946 25844 38948
rect 25788 38894 25790 38946
rect 25790 38894 25842 38946
rect 25842 38894 25844 38946
rect 25788 38892 25844 38894
rect 25676 38780 25732 38836
rect 25564 37826 25620 37828
rect 25564 37774 25566 37826
rect 25566 37774 25618 37826
rect 25618 37774 25620 37826
rect 25564 37772 25620 37774
rect 25676 36482 25732 36484
rect 25676 36430 25678 36482
rect 25678 36430 25730 36482
rect 25730 36430 25732 36482
rect 25676 36428 25732 36430
rect 25452 34130 25508 34132
rect 25452 34078 25454 34130
rect 25454 34078 25506 34130
rect 25506 34078 25508 34130
rect 25452 34076 25508 34078
rect 25900 34860 25956 34916
rect 25228 32396 25284 32452
rect 25452 29596 25508 29652
rect 25900 33906 25956 33908
rect 25900 33854 25902 33906
rect 25902 33854 25954 33906
rect 25954 33854 25956 33906
rect 25900 33852 25956 33854
rect 26236 38946 26292 38948
rect 26236 38894 26238 38946
rect 26238 38894 26290 38946
rect 26290 38894 26292 38946
rect 26236 38892 26292 38894
rect 26124 37996 26180 38052
rect 26124 37154 26180 37156
rect 26124 37102 26126 37154
rect 26126 37102 26178 37154
rect 26178 37102 26180 37154
rect 26124 37100 26180 37102
rect 26684 42700 26740 42756
rect 26908 45948 26964 46004
rect 27132 45218 27188 45220
rect 27132 45166 27134 45218
rect 27134 45166 27186 45218
rect 27186 45166 27188 45218
rect 27132 45164 27188 45166
rect 27020 43484 27076 43540
rect 26908 42924 26964 42980
rect 27244 43426 27300 43428
rect 27244 43374 27246 43426
rect 27246 43374 27298 43426
rect 27298 43374 27300 43426
rect 27244 43372 27300 43374
rect 27468 46562 27524 46564
rect 27468 46510 27470 46562
rect 27470 46510 27522 46562
rect 27522 46510 27524 46562
rect 27468 46508 27524 46510
rect 28028 55410 28084 55412
rect 28028 55358 28030 55410
rect 28030 55358 28082 55410
rect 28082 55358 28084 55410
rect 28028 55356 28084 55358
rect 27916 55132 27972 55188
rect 28476 56306 28532 56308
rect 28476 56254 28478 56306
rect 28478 56254 28530 56306
rect 28530 56254 28532 56306
rect 28476 56252 28532 56254
rect 27916 53788 27972 53844
rect 27916 53228 27972 53284
rect 28476 55132 28532 55188
rect 28140 54460 28196 54516
rect 28140 54012 28196 54068
rect 28252 53564 28308 53620
rect 28140 53452 28196 53508
rect 28028 50428 28084 50484
rect 28476 52220 28532 52276
rect 28252 50764 28308 50820
rect 28476 51212 28532 51268
rect 28700 57596 28756 57652
rect 28700 52668 28756 52724
rect 28924 57538 28980 57540
rect 28924 57486 28926 57538
rect 28926 57486 28978 57538
rect 28978 57486 28980 57538
rect 28924 57484 28980 57486
rect 29260 63810 29316 63812
rect 29260 63758 29262 63810
rect 29262 63758 29314 63810
rect 29314 63758 29316 63810
rect 29260 63756 29316 63758
rect 29932 65996 29988 66052
rect 30940 67788 30996 67844
rect 30604 66780 30660 66836
rect 31724 67618 31780 67620
rect 31724 67566 31726 67618
rect 31726 67566 31778 67618
rect 31778 67566 31780 67618
rect 31724 67564 31780 67566
rect 31052 67452 31108 67508
rect 30604 66274 30660 66276
rect 30604 66222 30606 66274
rect 30606 66222 30658 66274
rect 30658 66222 30660 66274
rect 30604 66220 30660 66222
rect 32732 72156 32788 72212
rect 33852 70588 33908 70644
rect 34972 71596 35028 71652
rect 34076 71036 34132 71092
rect 34860 71036 34916 71092
rect 34076 70588 34132 70644
rect 33404 68684 33460 68740
rect 33068 68572 33124 68628
rect 32396 68460 32452 68516
rect 32956 67676 33012 67732
rect 33404 67730 33460 67732
rect 33404 67678 33406 67730
rect 33406 67678 33458 67730
rect 33458 67678 33460 67730
rect 33404 67676 33460 67678
rect 32396 67564 32452 67620
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35532 71036 35588 71092
rect 35644 70812 35700 70868
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35644 69522 35700 69524
rect 35644 69470 35646 69522
rect 35646 69470 35698 69522
rect 35698 69470 35700 69522
rect 35644 69468 35700 69470
rect 35196 69186 35252 69188
rect 35196 69134 35198 69186
rect 35198 69134 35250 69186
rect 35250 69134 35252 69186
rect 35196 69132 35252 69134
rect 35868 71202 35924 71204
rect 35868 71150 35870 71202
rect 35870 71150 35922 71202
rect 35922 71150 35924 71202
rect 35868 71148 35924 71150
rect 36988 70866 37044 70868
rect 36988 70814 36990 70866
rect 36990 70814 37042 70866
rect 37042 70814 37044 70866
rect 36988 70812 37044 70814
rect 35980 70588 36036 70644
rect 37324 71650 37380 71652
rect 37324 71598 37326 71650
rect 37326 71598 37378 71650
rect 37378 71598 37380 71650
rect 37324 71596 37380 71598
rect 37996 71596 38052 71652
rect 37772 70476 37828 70532
rect 38892 70476 38948 70532
rect 36428 70028 36484 70084
rect 34300 68738 34356 68740
rect 34300 68686 34302 68738
rect 34302 68686 34354 68738
rect 34354 68686 34356 68738
rect 34300 68684 34356 68686
rect 34188 68626 34244 68628
rect 34188 68574 34190 68626
rect 34190 68574 34242 68626
rect 34242 68574 34244 68626
rect 34188 68572 34244 68574
rect 31836 66332 31892 66388
rect 31052 66050 31108 66052
rect 31052 65998 31054 66050
rect 31054 65998 31106 66050
rect 31106 65998 31108 66050
rect 31052 65996 31108 65998
rect 31276 66220 31332 66276
rect 29932 63756 29988 63812
rect 29484 63026 29540 63028
rect 29484 62974 29486 63026
rect 29486 62974 29538 63026
rect 29538 62974 29540 63026
rect 29484 62972 29540 62974
rect 29372 62860 29428 62916
rect 29372 62130 29428 62132
rect 29372 62078 29374 62130
rect 29374 62078 29426 62130
rect 29426 62078 29428 62130
rect 29372 62076 29428 62078
rect 29260 60674 29316 60676
rect 29260 60622 29262 60674
rect 29262 60622 29314 60674
rect 29314 60622 29316 60674
rect 29260 60620 29316 60622
rect 29148 58156 29204 58212
rect 29260 56866 29316 56868
rect 29260 56814 29262 56866
rect 29262 56814 29314 56866
rect 29314 56814 29316 56866
rect 29260 56812 29316 56814
rect 29036 56364 29092 56420
rect 29260 54402 29316 54404
rect 29260 54350 29262 54402
rect 29262 54350 29314 54402
rect 29314 54350 29316 54402
rect 29260 54348 29316 54350
rect 29148 53788 29204 53844
rect 30044 62860 30100 62916
rect 30380 63756 30436 63812
rect 29932 61682 29988 61684
rect 29932 61630 29934 61682
rect 29934 61630 29986 61682
rect 29986 61630 29988 61682
rect 29932 61628 29988 61630
rect 29596 58156 29652 58212
rect 28812 51436 28868 51492
rect 29036 51660 29092 51716
rect 28812 51154 28868 51156
rect 28812 51102 28814 51154
rect 28814 51102 28866 51154
rect 28866 51102 28868 51154
rect 28812 51100 28868 51102
rect 28364 50594 28420 50596
rect 28364 50542 28366 50594
rect 28366 50542 28418 50594
rect 28418 50542 28420 50594
rect 28364 50540 28420 50542
rect 27804 48972 27860 49028
rect 27804 48802 27860 48804
rect 27804 48750 27806 48802
rect 27806 48750 27858 48802
rect 27858 48750 27860 48802
rect 27804 48748 27860 48750
rect 26460 41916 26516 41972
rect 26684 41970 26740 41972
rect 26684 41918 26686 41970
rect 26686 41918 26738 41970
rect 26738 41918 26740 41970
rect 26684 41916 26740 41918
rect 27356 41916 27412 41972
rect 27468 41858 27524 41860
rect 27468 41806 27470 41858
rect 27470 41806 27522 41858
rect 27522 41806 27524 41858
rect 27468 41804 27524 41806
rect 26908 41020 26964 41076
rect 26460 40684 26516 40740
rect 26460 40460 26516 40516
rect 26796 38946 26852 38948
rect 26796 38894 26798 38946
rect 26798 38894 26850 38946
rect 26850 38894 26852 38946
rect 26796 38892 26852 38894
rect 26460 38834 26516 38836
rect 26460 38782 26462 38834
rect 26462 38782 26514 38834
rect 26514 38782 26516 38834
rect 26460 38780 26516 38782
rect 26236 35420 26292 35476
rect 26348 36876 26404 36932
rect 25564 29484 25620 29540
rect 25452 28812 25508 28868
rect 26572 37490 26628 37492
rect 26572 37438 26574 37490
rect 26574 37438 26626 37490
rect 26626 37438 26628 37490
rect 26572 37436 26628 37438
rect 26684 37378 26740 37380
rect 26684 37326 26686 37378
rect 26686 37326 26738 37378
rect 26738 37326 26740 37378
rect 26684 37324 26740 37326
rect 27468 38050 27524 38052
rect 27468 37998 27470 38050
rect 27470 37998 27522 38050
rect 27522 37998 27524 38050
rect 27468 37996 27524 37998
rect 27244 37490 27300 37492
rect 27244 37438 27246 37490
rect 27246 37438 27298 37490
rect 27298 37438 27300 37490
rect 27244 37436 27300 37438
rect 27020 37324 27076 37380
rect 27356 37100 27412 37156
rect 26572 35308 26628 35364
rect 26684 36988 26740 37044
rect 26236 29596 26292 29652
rect 26460 34300 26516 34356
rect 26348 29148 26404 29204
rect 26012 28812 26068 28868
rect 25564 27186 25620 27188
rect 25564 27134 25566 27186
rect 25566 27134 25618 27186
rect 25618 27134 25620 27186
rect 25564 27132 25620 27134
rect 25228 25004 25284 25060
rect 25452 24722 25508 24724
rect 25452 24670 25454 24722
rect 25454 24670 25506 24722
rect 25506 24670 25508 24722
rect 25452 24668 25508 24670
rect 25900 25004 25956 25060
rect 24892 20076 24948 20132
rect 25676 24332 25732 24388
rect 25452 23938 25508 23940
rect 25452 23886 25454 23938
rect 25454 23886 25506 23938
rect 25506 23886 25508 23938
rect 25452 23884 25508 23886
rect 25116 23826 25172 23828
rect 25116 23774 25118 23826
rect 25118 23774 25170 23826
rect 25170 23774 25172 23826
rect 25116 23772 25172 23774
rect 25788 23042 25844 23044
rect 25788 22990 25790 23042
rect 25790 22990 25842 23042
rect 25842 22990 25844 23042
rect 25788 22988 25844 22990
rect 26124 23996 26180 24052
rect 25900 22540 25956 22596
rect 26908 35644 26964 35700
rect 27356 36428 27412 36484
rect 26796 35586 26852 35588
rect 26796 35534 26798 35586
rect 26798 35534 26850 35586
rect 26850 35534 26852 35586
rect 26796 35532 26852 35534
rect 26796 29426 26852 29428
rect 26796 29374 26798 29426
rect 26798 29374 26850 29426
rect 26850 29374 26852 29426
rect 26796 29372 26852 29374
rect 26796 29036 26852 29092
rect 26348 24892 26404 24948
rect 26460 24780 26516 24836
rect 26460 23996 26516 24052
rect 26348 23660 26404 23716
rect 26124 22540 26180 22596
rect 26236 22316 26292 22372
rect 25228 20914 25284 20916
rect 25228 20862 25230 20914
rect 25230 20862 25282 20914
rect 25282 20862 25284 20914
rect 25228 20860 25284 20862
rect 25228 19906 25284 19908
rect 25228 19854 25230 19906
rect 25230 19854 25282 19906
rect 25282 19854 25284 19906
rect 25228 19852 25284 19854
rect 25788 20860 25844 20916
rect 26124 21698 26180 21700
rect 26124 21646 26126 21698
rect 26126 21646 26178 21698
rect 26178 21646 26180 21698
rect 26124 21644 26180 21646
rect 26236 20972 26292 21028
rect 26124 20802 26180 20804
rect 26124 20750 26126 20802
rect 26126 20750 26178 20802
rect 26178 20750 26180 20802
rect 26124 20748 26180 20750
rect 25676 20578 25732 20580
rect 25676 20526 25678 20578
rect 25678 20526 25730 20578
rect 25730 20526 25732 20578
rect 25676 20524 25732 20526
rect 25564 20076 25620 20132
rect 26684 23154 26740 23156
rect 26684 23102 26686 23154
rect 26686 23102 26738 23154
rect 26738 23102 26740 23154
rect 26684 23100 26740 23102
rect 26572 20972 26628 21028
rect 25452 19234 25508 19236
rect 25452 19182 25454 19234
rect 25454 19182 25506 19234
rect 25506 19182 25508 19234
rect 25452 19180 25508 19182
rect 26124 19234 26180 19236
rect 26124 19182 26126 19234
rect 26126 19182 26178 19234
rect 26178 19182 26180 19234
rect 26124 19180 26180 19182
rect 25228 18396 25284 18452
rect 26236 18396 26292 18452
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 25004 17724 25060 17780
rect 25116 17666 25172 17668
rect 25116 17614 25118 17666
rect 25118 17614 25170 17666
rect 25170 17614 25172 17666
rect 25116 17612 25172 17614
rect 24892 16210 24948 16212
rect 24892 16158 24894 16210
rect 24894 16158 24946 16210
rect 24946 16158 24948 16210
rect 24892 16156 24948 16158
rect 25564 17666 25620 17668
rect 25564 17614 25566 17666
rect 25566 17614 25618 17666
rect 25618 17614 25620 17666
rect 25564 17612 25620 17614
rect 26236 17052 26292 17108
rect 25788 16268 25844 16324
rect 25340 15538 25396 15540
rect 25340 15486 25342 15538
rect 25342 15486 25394 15538
rect 25394 15486 25396 15538
rect 25340 15484 25396 15486
rect 25900 16210 25956 16212
rect 25900 16158 25902 16210
rect 25902 16158 25954 16210
rect 25954 16158 25956 16210
rect 25900 16156 25956 16158
rect 25788 15260 25844 15316
rect 25900 15036 25956 15092
rect 25564 14476 25620 14532
rect 25228 13804 25284 13860
rect 25676 14364 25732 14420
rect 25340 12684 25396 12740
rect 26460 15092 26516 15148
rect 25452 12402 25508 12404
rect 25452 12350 25454 12402
rect 25454 12350 25506 12402
rect 25506 12350 25508 12402
rect 25452 12348 25508 12350
rect 25004 11788 25060 11844
rect 25116 11116 25172 11172
rect 24780 10834 24836 10836
rect 24780 10782 24782 10834
rect 24782 10782 24834 10834
rect 24834 10782 24836 10834
rect 24780 10780 24836 10782
rect 22428 8316 22484 8372
rect 22316 8258 22372 8260
rect 22316 8206 22318 8258
rect 22318 8206 22370 8258
rect 22370 8206 22372 8258
rect 22316 8204 22372 8206
rect 21868 7586 21924 7588
rect 21868 7534 21870 7586
rect 21870 7534 21922 7586
rect 21922 7534 21924 7586
rect 21868 7532 21924 7534
rect 22876 7980 22932 8036
rect 21532 5068 21588 5124
rect 23772 8258 23828 8260
rect 23772 8206 23774 8258
rect 23774 8206 23826 8258
rect 23826 8206 23828 8258
rect 23772 8204 23828 8206
rect 23660 7980 23716 8036
rect 24108 7420 24164 7476
rect 24332 6860 24388 6916
rect 24556 5852 24612 5908
rect 22316 5628 22372 5684
rect 24332 5180 24388 5236
rect 22316 5068 22372 5124
rect 22652 5068 22708 5124
rect 23772 4956 23828 5012
rect 23548 4338 23604 4340
rect 23548 4286 23550 4338
rect 23550 4286 23602 4338
rect 23602 4286 23604 4338
rect 23548 4284 23604 4286
rect 22988 3666 23044 3668
rect 22988 3614 22990 3666
rect 22990 3614 23042 3666
rect 23042 3614 23044 3666
rect 22988 3612 23044 3614
rect 27132 34972 27188 35028
rect 27020 34748 27076 34804
rect 27020 31612 27076 31668
rect 27356 35308 27412 35364
rect 27020 30156 27076 30212
rect 27020 28588 27076 28644
rect 27020 28364 27076 28420
rect 27244 31612 27300 31668
rect 27244 30210 27300 30212
rect 27244 30158 27246 30210
rect 27246 30158 27298 30210
rect 27298 30158 27300 30210
rect 27244 30156 27300 30158
rect 27468 32284 27524 32340
rect 27468 31612 27524 31668
rect 27692 42754 27748 42756
rect 27692 42702 27694 42754
rect 27694 42702 27746 42754
rect 27746 42702 27748 42754
rect 27692 42700 27748 42702
rect 27804 37548 27860 37604
rect 27804 36428 27860 36484
rect 27804 35698 27860 35700
rect 27804 35646 27806 35698
rect 27806 35646 27858 35698
rect 27858 35646 27860 35698
rect 27804 35644 27860 35646
rect 28252 50204 28308 50260
rect 28028 49868 28084 49924
rect 28028 48748 28084 48804
rect 28588 50370 28644 50372
rect 28588 50318 28590 50370
rect 28590 50318 28642 50370
rect 28642 50318 28644 50370
rect 28588 50316 28644 50318
rect 28364 49756 28420 49812
rect 28588 49698 28644 49700
rect 28588 49646 28590 49698
rect 28590 49646 28642 49698
rect 28642 49646 28644 49698
rect 28588 49644 28644 49646
rect 28252 47068 28308 47124
rect 28140 45276 28196 45332
rect 28028 42364 28084 42420
rect 28028 37266 28084 37268
rect 28028 37214 28030 37266
rect 28030 37214 28082 37266
rect 28082 37214 28084 37266
rect 28028 37212 28084 37214
rect 28588 47068 28644 47124
rect 29036 50482 29092 50484
rect 29036 50430 29038 50482
rect 29038 50430 29090 50482
rect 29090 50430 29092 50482
rect 29036 50428 29092 50430
rect 28924 50316 28980 50372
rect 29484 52780 29540 52836
rect 29260 52162 29316 52164
rect 29260 52110 29262 52162
rect 29262 52110 29314 52162
rect 29314 52110 29316 52162
rect 29260 52108 29316 52110
rect 29372 51660 29428 51716
rect 29260 50316 29316 50372
rect 29148 49026 29204 49028
rect 29148 48974 29150 49026
rect 29150 48974 29202 49026
rect 29202 48974 29204 49026
rect 29148 48972 29204 48974
rect 28252 37548 28308 37604
rect 29148 46732 29204 46788
rect 28700 45388 28756 45444
rect 28700 40572 28756 40628
rect 28700 40348 28756 40404
rect 28700 40012 28756 40068
rect 28700 38444 28756 38500
rect 29260 45612 29316 45668
rect 29708 56642 29764 56644
rect 29708 56590 29710 56642
rect 29710 56590 29762 56642
rect 29762 56590 29764 56642
rect 29708 56588 29764 56590
rect 29708 55692 29764 55748
rect 29596 46732 29652 46788
rect 29708 52108 29764 52164
rect 29596 46562 29652 46564
rect 29596 46510 29598 46562
rect 29598 46510 29650 46562
rect 29650 46510 29652 46562
rect 29596 46508 29652 46510
rect 29484 45388 29540 45444
rect 29484 45052 29540 45108
rect 30492 63698 30548 63700
rect 30492 63646 30494 63698
rect 30494 63646 30546 63698
rect 30546 63646 30548 63698
rect 30492 63644 30548 63646
rect 31164 63644 31220 63700
rect 30940 63308 30996 63364
rect 30492 62300 30548 62356
rect 31164 62188 31220 62244
rect 32172 66386 32228 66388
rect 32172 66334 32174 66386
rect 32174 66334 32226 66386
rect 32226 66334 32228 66386
rect 32172 66332 32228 66334
rect 32060 66274 32116 66276
rect 32060 66222 32062 66274
rect 32062 66222 32114 66274
rect 32114 66222 32116 66274
rect 32060 66220 32116 66222
rect 34076 67676 34132 67732
rect 36316 69298 36372 69300
rect 36316 69246 36318 69298
rect 36318 69246 36370 69298
rect 36370 69246 36372 69298
rect 36316 69244 36372 69246
rect 35196 68514 35252 68516
rect 35196 68462 35198 68514
rect 35198 68462 35250 68514
rect 35250 68462 35252 68514
rect 35196 68460 35252 68462
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 37660 70028 37716 70084
rect 37772 70140 37828 70196
rect 37324 69244 37380 69300
rect 35756 68514 35812 68516
rect 35756 68462 35758 68514
rect 35758 68462 35810 68514
rect 35810 68462 35812 68514
rect 35756 68460 35812 68462
rect 35644 67452 35700 67508
rect 32844 66274 32900 66276
rect 32844 66222 32846 66274
rect 32846 66222 32898 66274
rect 32898 66222 32900 66274
rect 32844 66220 32900 66222
rect 31836 65548 31892 65604
rect 31948 63362 32004 63364
rect 31948 63310 31950 63362
rect 31950 63310 32002 63362
rect 32002 63310 32004 63362
rect 31948 63308 32004 63310
rect 31388 62354 31444 62356
rect 31388 62302 31390 62354
rect 31390 62302 31442 62354
rect 31442 62302 31444 62354
rect 31388 62300 31444 62302
rect 31724 62076 31780 62132
rect 32396 65660 32452 65716
rect 32284 65436 32340 65492
rect 32508 65324 32564 65380
rect 32284 63532 32340 63588
rect 32060 62188 32116 62244
rect 31612 61628 31668 61684
rect 31500 61404 31556 61460
rect 31388 61010 31444 61012
rect 31388 60958 31390 61010
rect 31390 60958 31442 61010
rect 31442 60958 31444 61010
rect 31388 60956 31444 60958
rect 31948 60898 32004 60900
rect 31948 60846 31950 60898
rect 31950 60846 32002 60898
rect 32002 60846 32004 60898
rect 31948 60844 32004 60846
rect 31052 59052 31108 59108
rect 31612 60562 31668 60564
rect 31612 60510 31614 60562
rect 31614 60510 31666 60562
rect 31666 60510 31668 60562
rect 31612 60508 31668 60510
rect 31836 60620 31892 60676
rect 31724 59890 31780 59892
rect 31724 59838 31726 59890
rect 31726 59838 31778 59890
rect 31778 59838 31780 59890
rect 31724 59836 31780 59838
rect 31276 59778 31332 59780
rect 31276 59726 31278 59778
rect 31278 59726 31330 59778
rect 31330 59726 31332 59778
rect 31276 59724 31332 59726
rect 31612 59778 31668 59780
rect 31612 59726 31614 59778
rect 31614 59726 31666 59778
rect 31666 59726 31668 59778
rect 31612 59724 31668 59726
rect 31388 59612 31444 59668
rect 31276 59330 31332 59332
rect 31276 59278 31278 59330
rect 31278 59278 31330 59330
rect 31330 59278 31332 59330
rect 31276 59276 31332 59278
rect 30268 57148 30324 57204
rect 30492 57260 30548 57316
rect 30156 57036 30212 57092
rect 30716 57148 30772 57204
rect 29932 53730 29988 53732
rect 29932 53678 29934 53730
rect 29934 53678 29986 53730
rect 29986 53678 29988 53730
rect 29932 53676 29988 53678
rect 29820 51548 29876 51604
rect 29820 50706 29876 50708
rect 29820 50654 29822 50706
rect 29822 50654 29874 50706
rect 29874 50654 29876 50706
rect 29820 50652 29876 50654
rect 29932 48914 29988 48916
rect 29932 48862 29934 48914
rect 29934 48862 29986 48914
rect 29986 48862 29988 48914
rect 29932 48860 29988 48862
rect 31052 57260 31108 57316
rect 31276 57036 31332 57092
rect 31612 56588 31668 56644
rect 31724 59052 31780 59108
rect 35308 67058 35364 67060
rect 35308 67006 35310 67058
rect 35310 67006 35362 67058
rect 35362 67006 35364 67058
rect 35308 67004 35364 67006
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 34300 66332 34356 66388
rect 33404 66274 33460 66276
rect 33404 66222 33406 66274
rect 33406 66222 33458 66274
rect 33458 66222 33460 66274
rect 33404 66220 33460 66222
rect 34412 66220 34468 66276
rect 33740 65660 33796 65716
rect 34524 65548 34580 65604
rect 33628 65490 33684 65492
rect 33628 65438 33630 65490
rect 33630 65438 33682 65490
rect 33682 65438 33684 65490
rect 33628 65436 33684 65438
rect 33180 65378 33236 65380
rect 33180 65326 33182 65378
rect 33182 65326 33234 65378
rect 33234 65326 33236 65378
rect 33180 65324 33236 65326
rect 34412 64818 34468 64820
rect 34412 64766 34414 64818
rect 34414 64766 34466 64818
rect 34466 64766 34468 64818
rect 34412 64764 34468 64766
rect 34188 62972 34244 63028
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 36316 67004 36372 67060
rect 35420 64818 35476 64820
rect 35420 64766 35422 64818
rect 35422 64766 35474 64818
rect 35474 64766 35476 64818
rect 35420 64764 35476 64766
rect 34300 63084 34356 63140
rect 33180 62354 33236 62356
rect 33180 62302 33182 62354
rect 33182 62302 33234 62354
rect 33234 62302 33236 62354
rect 33180 62300 33236 62302
rect 32620 61458 32676 61460
rect 32620 61406 32622 61458
rect 32622 61406 32674 61458
rect 32674 61406 32676 61458
rect 32620 61404 32676 61406
rect 32620 60732 32676 60788
rect 32172 60674 32228 60676
rect 32172 60622 32174 60674
rect 32174 60622 32226 60674
rect 32226 60622 32228 60674
rect 32172 60620 32228 60622
rect 32508 60508 32564 60564
rect 32172 59890 32228 59892
rect 32172 59838 32174 59890
rect 32174 59838 32226 59890
rect 32226 59838 32228 59890
rect 32172 59836 32228 59838
rect 32396 59778 32452 59780
rect 32396 59726 32398 59778
rect 32398 59726 32450 59778
rect 32450 59726 32452 59778
rect 32396 59724 32452 59726
rect 33180 60956 33236 61012
rect 33628 60844 33684 60900
rect 32956 60508 33012 60564
rect 33404 60508 33460 60564
rect 33180 60284 33236 60340
rect 32172 59052 32228 59108
rect 30716 56140 30772 56196
rect 30604 55970 30660 55972
rect 30604 55918 30606 55970
rect 30606 55918 30658 55970
rect 30658 55918 30660 55970
rect 30604 55916 30660 55918
rect 30604 55692 30660 55748
rect 30156 52780 30212 52836
rect 30268 52332 30324 52388
rect 30268 51266 30324 51268
rect 30268 51214 30270 51266
rect 30270 51214 30322 51266
rect 30322 51214 30324 51266
rect 30268 51212 30324 51214
rect 30268 50594 30324 50596
rect 30268 50542 30270 50594
rect 30270 50542 30322 50594
rect 30322 50542 30324 50594
rect 30268 50540 30324 50542
rect 30044 48524 30100 48580
rect 30380 50204 30436 50260
rect 30268 47292 30324 47348
rect 29708 45500 29764 45556
rect 30268 45388 30324 45444
rect 29932 45052 29988 45108
rect 30044 45164 30100 45220
rect 29708 44828 29764 44884
rect 29708 44492 29764 44548
rect 30156 45106 30212 45108
rect 30156 45054 30158 45106
rect 30158 45054 30210 45106
rect 30210 45054 30212 45106
rect 30156 45052 30212 45054
rect 29708 43596 29764 43652
rect 29820 41916 29876 41972
rect 29596 41858 29652 41860
rect 29596 41806 29598 41858
rect 29598 41806 29650 41858
rect 29650 41806 29652 41858
rect 29596 41804 29652 41806
rect 28588 38220 28644 38276
rect 28476 38162 28532 38164
rect 28476 38110 28478 38162
rect 28478 38110 28530 38162
rect 28530 38110 28532 38162
rect 28476 38108 28532 38110
rect 29596 38946 29652 38948
rect 29596 38894 29598 38946
rect 29598 38894 29650 38946
rect 29650 38894 29652 38946
rect 29596 38892 29652 38894
rect 30716 52834 30772 52836
rect 30716 52782 30718 52834
rect 30718 52782 30770 52834
rect 30770 52782 30772 52834
rect 30716 52780 30772 52782
rect 31052 50316 31108 50372
rect 30604 48860 30660 48916
rect 30716 48748 30772 48804
rect 30716 47292 30772 47348
rect 30492 45276 30548 45332
rect 30156 40684 30212 40740
rect 30380 40236 30436 40292
rect 30380 40012 30436 40068
rect 30828 45778 30884 45780
rect 30828 45726 30830 45778
rect 30830 45726 30882 45778
rect 30882 45726 30884 45778
rect 30828 45724 30884 45726
rect 30828 45164 30884 45220
rect 30716 45052 30772 45108
rect 30716 44322 30772 44324
rect 30716 44270 30718 44322
rect 30718 44270 30770 44322
rect 30770 44270 30772 44322
rect 30716 44268 30772 44270
rect 31500 56140 31556 56196
rect 31388 53228 31444 53284
rect 31388 52780 31444 52836
rect 31612 56028 31668 56084
rect 32172 55356 32228 55412
rect 32060 54348 32116 54404
rect 31612 53564 31668 53620
rect 31836 53452 31892 53508
rect 31724 52162 31780 52164
rect 31724 52110 31726 52162
rect 31726 52110 31778 52162
rect 31778 52110 31780 52162
rect 31724 52108 31780 52110
rect 31500 51100 31556 51156
rect 31612 51996 31668 52052
rect 32172 52780 32228 52836
rect 32284 52274 32340 52276
rect 32284 52222 32286 52274
rect 32286 52222 32338 52274
rect 32338 52222 32340 52274
rect 32284 52220 32340 52222
rect 32172 52108 32228 52164
rect 32620 59276 32676 59332
rect 32956 59052 33012 59108
rect 33180 59724 33236 59780
rect 33740 60284 33796 60340
rect 33852 60620 33908 60676
rect 33516 59106 33572 59108
rect 33516 59054 33518 59106
rect 33518 59054 33570 59106
rect 33570 59054 33572 59106
rect 33516 59052 33572 59054
rect 34076 59778 34132 59780
rect 34076 59726 34078 59778
rect 34078 59726 34130 59778
rect 34130 59726 34132 59778
rect 34076 59724 34132 59726
rect 33964 59052 34020 59108
rect 34188 59052 34244 59108
rect 33516 57596 33572 57652
rect 32844 55916 32900 55972
rect 32508 55244 32564 55300
rect 32956 53788 33012 53844
rect 33516 55298 33572 55300
rect 33516 55246 33518 55298
rect 33518 55246 33570 55298
rect 33570 55246 33572 55298
rect 33516 55244 33572 55246
rect 33292 55132 33348 55188
rect 33516 54908 33572 54964
rect 33740 54796 33796 54852
rect 34076 57650 34132 57652
rect 34076 57598 34078 57650
rect 34078 57598 34130 57650
rect 34130 57598 34132 57650
rect 34076 57596 34132 57598
rect 34188 55186 34244 55188
rect 34188 55134 34190 55186
rect 34190 55134 34242 55186
rect 34242 55134 34244 55186
rect 34188 55132 34244 55134
rect 33964 54908 34020 54964
rect 34076 55020 34132 55076
rect 34188 54796 34244 54852
rect 33516 53788 33572 53844
rect 33404 53506 33460 53508
rect 33404 53454 33406 53506
rect 33406 53454 33458 53506
rect 33458 53454 33460 53506
rect 33404 53452 33460 53454
rect 32620 52050 32676 52052
rect 32620 51998 32622 52050
rect 32622 51998 32674 52050
rect 32674 51998 32676 52050
rect 32620 51996 32676 51998
rect 32732 51884 32788 51940
rect 32508 51324 32564 51380
rect 31724 50316 31780 50372
rect 31500 49644 31556 49700
rect 31388 49084 31444 49140
rect 31724 48860 31780 48916
rect 31500 46508 31556 46564
rect 31164 45500 31220 45556
rect 31388 45276 31444 45332
rect 31052 41020 31108 41076
rect 30940 40684 30996 40740
rect 31836 48636 31892 48692
rect 31724 47516 31780 47572
rect 30828 40402 30884 40404
rect 30828 40350 30830 40402
rect 30830 40350 30882 40402
rect 30882 40350 30884 40402
rect 30828 40348 30884 40350
rect 29036 38332 29092 38388
rect 28812 37996 28868 38052
rect 28924 38220 28980 38276
rect 28588 37212 28644 37268
rect 28364 37100 28420 37156
rect 28476 35756 28532 35812
rect 27692 34972 27748 35028
rect 27916 34524 27972 34580
rect 27356 29538 27412 29540
rect 27356 29486 27358 29538
rect 27358 29486 27410 29538
rect 27410 29486 27412 29538
rect 27356 29484 27412 29486
rect 28700 36316 28756 36372
rect 28252 35308 28308 35364
rect 28364 34748 28420 34804
rect 28476 34524 28532 34580
rect 28252 32786 28308 32788
rect 28252 32734 28254 32786
rect 28254 32734 28306 32786
rect 28306 32734 28308 32786
rect 28252 32732 28308 32734
rect 27580 28866 27636 28868
rect 27580 28814 27582 28866
rect 27582 28814 27634 28866
rect 27634 28814 27636 28866
rect 27580 28812 27636 28814
rect 27580 28642 27636 28644
rect 27580 28590 27582 28642
rect 27582 28590 27634 28642
rect 27634 28590 27636 28642
rect 27580 28588 27636 28590
rect 26908 22092 26964 22148
rect 27020 26684 27076 26740
rect 27132 25452 27188 25508
rect 27132 24834 27188 24836
rect 27132 24782 27134 24834
rect 27134 24782 27186 24834
rect 27186 24782 27188 24834
rect 27132 24780 27188 24782
rect 27468 26066 27524 26068
rect 27468 26014 27470 26066
rect 27470 26014 27522 26066
rect 27522 26014 27524 26066
rect 27468 26012 27524 26014
rect 27692 26850 27748 26852
rect 27692 26798 27694 26850
rect 27694 26798 27746 26850
rect 27746 26798 27748 26850
rect 27692 26796 27748 26798
rect 27468 25452 27524 25508
rect 27692 24892 27748 24948
rect 26908 21084 26964 21140
rect 27020 21026 27076 21028
rect 27020 20974 27022 21026
rect 27022 20974 27074 21026
rect 27074 20974 27076 21026
rect 27020 20972 27076 20974
rect 26796 18396 26852 18452
rect 26572 14418 26628 14420
rect 26572 14366 26574 14418
rect 26574 14366 26626 14418
rect 26626 14366 26628 14418
rect 26572 14364 26628 14366
rect 26908 14418 26964 14420
rect 26908 14366 26910 14418
rect 26910 14366 26962 14418
rect 26962 14366 26964 14418
rect 26908 14364 26964 14366
rect 27580 23324 27636 23380
rect 27580 23154 27636 23156
rect 27580 23102 27582 23154
rect 27582 23102 27634 23154
rect 27634 23102 27636 23154
rect 27580 23100 27636 23102
rect 27244 22370 27300 22372
rect 27244 22318 27246 22370
rect 27246 22318 27298 22370
rect 27298 22318 27300 22370
rect 27244 22316 27300 22318
rect 27244 22092 27300 22148
rect 27244 21084 27300 21140
rect 27356 20636 27412 20692
rect 27244 20130 27300 20132
rect 27244 20078 27246 20130
rect 27246 20078 27298 20130
rect 27298 20078 27300 20130
rect 27244 20076 27300 20078
rect 27468 18620 27524 18676
rect 27468 18284 27524 18340
rect 28252 30210 28308 30212
rect 28252 30158 28254 30210
rect 28254 30158 28306 30210
rect 28306 30158 28308 30210
rect 28252 30156 28308 30158
rect 28028 30044 28084 30100
rect 28028 28364 28084 28420
rect 28252 28588 28308 28644
rect 28588 31666 28644 31668
rect 28588 31614 28590 31666
rect 28590 31614 28642 31666
rect 28642 31614 28644 31666
rect 28588 31612 28644 31614
rect 28476 30828 28532 30884
rect 28476 30044 28532 30100
rect 28476 27916 28532 27972
rect 28812 31164 28868 31220
rect 29148 37884 29204 37940
rect 29596 38050 29652 38052
rect 29596 37998 29598 38050
rect 29598 37998 29650 38050
rect 29650 37998 29652 38050
rect 29596 37996 29652 37998
rect 30716 39676 30772 39732
rect 29260 37154 29316 37156
rect 29260 37102 29262 37154
rect 29262 37102 29314 37154
rect 29314 37102 29316 37154
rect 29260 37100 29316 37102
rect 29932 37884 29988 37940
rect 30044 37996 30100 38052
rect 29596 37772 29652 37828
rect 29596 37266 29652 37268
rect 29596 37214 29598 37266
rect 29598 37214 29650 37266
rect 29650 37214 29652 37266
rect 29596 37212 29652 37214
rect 29484 37100 29540 37156
rect 30156 36988 30212 37044
rect 30044 36876 30100 36932
rect 29932 35810 29988 35812
rect 29932 35758 29934 35810
rect 29934 35758 29986 35810
rect 29986 35758 29988 35810
rect 29932 35756 29988 35758
rect 29484 35644 29540 35700
rect 30044 35644 30100 35700
rect 30156 36652 30212 36708
rect 29036 34972 29092 35028
rect 29484 34748 29540 34804
rect 29036 34524 29092 34580
rect 29260 34524 29316 34580
rect 29260 32508 29316 32564
rect 29484 31666 29540 31668
rect 29484 31614 29486 31666
rect 29486 31614 29538 31666
rect 29538 31614 29540 31666
rect 29484 31612 29540 31614
rect 29036 30994 29092 30996
rect 29036 30942 29038 30994
rect 29038 30942 29090 30994
rect 29090 30942 29092 30994
rect 29036 30940 29092 30942
rect 28700 30380 28756 30436
rect 29260 30156 29316 30212
rect 29372 30098 29428 30100
rect 29372 30046 29374 30098
rect 29374 30046 29426 30098
rect 29426 30046 29428 30098
rect 29372 30044 29428 30046
rect 30044 35420 30100 35476
rect 29596 29820 29652 29876
rect 29708 35308 29764 35364
rect 29932 35084 29988 35140
rect 29820 34802 29876 34804
rect 29820 34750 29822 34802
rect 29822 34750 29874 34802
rect 29874 34750 29876 34802
rect 29820 34748 29876 34750
rect 30492 37826 30548 37828
rect 30492 37774 30494 37826
rect 30494 37774 30546 37826
rect 30546 37774 30548 37826
rect 30492 37772 30548 37774
rect 30492 35084 30548 35140
rect 30156 33964 30212 34020
rect 30940 38946 30996 38948
rect 30940 38894 30942 38946
rect 30942 38894 30994 38946
rect 30994 38894 30996 38946
rect 30940 38892 30996 38894
rect 31164 40348 31220 40404
rect 30828 37212 30884 37268
rect 30716 35644 30772 35700
rect 31052 37100 31108 37156
rect 31500 41970 31556 41972
rect 31500 41918 31502 41970
rect 31502 41918 31554 41970
rect 31554 41918 31556 41970
rect 31500 41916 31556 41918
rect 31388 41074 31444 41076
rect 31388 41022 31390 41074
rect 31390 41022 31442 41074
rect 31442 41022 31444 41074
rect 31388 41020 31444 41022
rect 31388 40796 31444 40852
rect 31612 40684 31668 40740
rect 31500 39676 31556 39732
rect 32060 49138 32116 49140
rect 32060 49086 32062 49138
rect 32062 49086 32114 49138
rect 32114 49086 32116 49138
rect 32060 49084 32116 49086
rect 32844 51324 32900 51380
rect 32732 49756 32788 49812
rect 32620 48972 32676 49028
rect 32396 48914 32452 48916
rect 32396 48862 32398 48914
rect 32398 48862 32450 48914
rect 32450 48862 32452 48914
rect 32396 48860 32452 48862
rect 32284 47292 32340 47348
rect 32060 45778 32116 45780
rect 32060 45726 32062 45778
rect 32062 45726 32114 45778
rect 32114 45726 32116 45778
rect 32060 45724 32116 45726
rect 32060 45218 32116 45220
rect 32060 45166 32062 45218
rect 32062 45166 32114 45218
rect 32114 45166 32116 45218
rect 32060 45164 32116 45166
rect 31836 45106 31892 45108
rect 31836 45054 31838 45106
rect 31838 45054 31890 45106
rect 31890 45054 31892 45106
rect 31836 45052 31892 45054
rect 31948 44268 32004 44324
rect 32284 45500 32340 45556
rect 31948 42028 32004 42084
rect 31948 41804 32004 41860
rect 31948 40626 32004 40628
rect 31948 40574 31950 40626
rect 31950 40574 32002 40626
rect 32002 40574 32004 40626
rect 31948 40572 32004 40574
rect 32396 44434 32452 44436
rect 32396 44382 32398 44434
rect 32398 44382 32450 44434
rect 32450 44382 32452 44434
rect 32396 44380 32452 44382
rect 32396 41916 32452 41972
rect 32396 41244 32452 41300
rect 32396 40684 32452 40740
rect 32396 40348 32452 40404
rect 32732 48748 32788 48804
rect 32732 45612 32788 45668
rect 33404 53004 33460 53060
rect 33404 52220 33460 52276
rect 34636 63756 34692 63812
rect 34860 60898 34916 60900
rect 34860 60846 34862 60898
rect 34862 60846 34914 60898
rect 34914 60846 34916 60898
rect 34860 60844 34916 60846
rect 34748 60786 34804 60788
rect 34748 60734 34750 60786
rect 34750 60734 34802 60786
rect 34802 60734 34804 60786
rect 34748 60732 34804 60734
rect 34972 60786 35028 60788
rect 34972 60734 34974 60786
rect 34974 60734 35026 60786
rect 35026 60734 35028 60786
rect 34972 60732 35028 60734
rect 34860 60002 34916 60004
rect 34860 59950 34862 60002
rect 34862 59950 34914 60002
rect 34914 59950 34916 60002
rect 34860 59948 34916 59950
rect 34972 59500 35028 59556
rect 34412 55298 34468 55300
rect 34412 55246 34414 55298
rect 34414 55246 34466 55298
rect 34466 55246 34468 55298
rect 34412 55244 34468 55246
rect 33740 53058 33796 53060
rect 33740 53006 33742 53058
rect 33742 53006 33794 53058
rect 33794 53006 33796 53058
rect 33740 53004 33796 53006
rect 33628 52668 33684 52724
rect 33292 50652 33348 50708
rect 34300 52668 34356 52724
rect 34412 51324 34468 51380
rect 33964 50706 34020 50708
rect 33964 50654 33966 50706
rect 33966 50654 34018 50706
rect 34018 50654 34020 50706
rect 33964 50652 34020 50654
rect 33180 50316 33236 50372
rect 33404 50316 33460 50372
rect 33068 49810 33124 49812
rect 33068 49758 33070 49810
rect 33070 49758 33122 49810
rect 33122 49758 33124 49810
rect 33068 49756 33124 49758
rect 32956 48914 33012 48916
rect 32956 48862 32958 48914
rect 32958 48862 33010 48914
rect 33010 48862 33012 48914
rect 32956 48860 33012 48862
rect 33068 47740 33124 47796
rect 33180 49644 33236 49700
rect 32956 47516 33012 47572
rect 32956 47346 33012 47348
rect 32956 47294 32958 47346
rect 32958 47294 33010 47346
rect 33010 47294 33012 47346
rect 32956 47292 33012 47294
rect 33404 49922 33460 49924
rect 33404 49870 33406 49922
rect 33406 49870 33458 49922
rect 33458 49870 33460 49922
rect 33404 49868 33460 49870
rect 33740 49810 33796 49812
rect 33740 49758 33742 49810
rect 33742 49758 33794 49810
rect 33794 49758 33796 49810
rect 33740 49756 33796 49758
rect 33292 48802 33348 48804
rect 33292 48750 33294 48802
rect 33294 48750 33346 48802
rect 33346 48750 33348 48802
rect 33292 48748 33348 48750
rect 33180 46732 33236 46788
rect 33628 48914 33684 48916
rect 33628 48862 33630 48914
rect 33630 48862 33682 48914
rect 33682 48862 33684 48914
rect 33628 48860 33684 48862
rect 33852 48300 33908 48356
rect 34188 50316 34244 50372
rect 33628 47570 33684 47572
rect 33628 47518 33630 47570
rect 33630 47518 33682 47570
rect 33682 47518 33684 47570
rect 33628 47516 33684 47518
rect 33852 47458 33908 47460
rect 33852 47406 33854 47458
rect 33854 47406 33906 47458
rect 33906 47406 33908 47458
rect 33852 47404 33908 47406
rect 33852 47068 33908 47124
rect 33628 46732 33684 46788
rect 33068 45052 33124 45108
rect 33404 45612 33460 45668
rect 34300 49922 34356 49924
rect 34300 49870 34302 49922
rect 34302 49870 34354 49922
rect 34354 49870 34356 49922
rect 34300 49868 34356 49870
rect 34300 48748 34356 48804
rect 34636 55244 34692 55300
rect 35756 63980 35812 64036
rect 35196 63810 35252 63812
rect 35196 63758 35198 63810
rect 35198 63758 35250 63810
rect 35250 63758 35252 63810
rect 35196 63756 35252 63758
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35420 63138 35476 63140
rect 35420 63086 35422 63138
rect 35422 63086 35474 63138
rect 35474 63086 35476 63138
rect 35420 63084 35476 63086
rect 35196 63026 35252 63028
rect 35196 62974 35198 63026
rect 35198 62974 35250 63026
rect 35250 62974 35252 63026
rect 35196 62972 35252 62974
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35756 60732 35812 60788
rect 35308 60508 35364 60564
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 60172 35252 60228
rect 39004 70140 39060 70196
rect 37996 69916 38052 69972
rect 38780 69970 38836 69972
rect 38780 69918 38782 69970
rect 38782 69918 38834 69970
rect 38834 69918 38836 69970
rect 38780 69916 38836 69918
rect 42028 72268 42084 72324
rect 44380 74956 44436 75012
rect 40348 70700 40404 70756
rect 41804 70252 41860 70308
rect 39564 70194 39620 70196
rect 39564 70142 39566 70194
rect 39566 70142 39618 70194
rect 39618 70142 39620 70194
rect 39564 70140 39620 70142
rect 41692 70140 41748 70196
rect 38444 69634 38500 69636
rect 38444 69582 38446 69634
rect 38446 69582 38498 69634
rect 38498 69582 38500 69634
rect 38444 69580 38500 69582
rect 39004 69468 39060 69524
rect 37772 69132 37828 69188
rect 38668 68626 38724 68628
rect 38668 68574 38670 68626
rect 38670 68574 38722 68626
rect 38722 68574 38724 68626
rect 38668 68572 38724 68574
rect 37436 68460 37492 68516
rect 38780 68402 38836 68404
rect 38780 68350 38782 68402
rect 38782 68350 38834 68402
rect 38834 68350 38836 68402
rect 38780 68348 38836 68350
rect 39228 68572 39284 68628
rect 39564 68626 39620 68628
rect 39564 68574 39566 68626
rect 39566 68574 39618 68626
rect 39618 68574 39620 68626
rect 39564 68572 39620 68574
rect 40572 68348 40628 68404
rect 40908 67730 40964 67732
rect 40908 67678 40910 67730
rect 40910 67678 40962 67730
rect 40962 67678 40964 67730
rect 40908 67676 40964 67678
rect 42252 67676 42308 67732
rect 43596 67730 43652 67732
rect 43596 67678 43598 67730
rect 43598 67678 43650 67730
rect 43650 67678 43652 67730
rect 43596 67676 43652 67678
rect 37548 66332 37604 66388
rect 37436 66220 37492 66276
rect 38332 66220 38388 66276
rect 37548 66162 37604 66164
rect 37548 66110 37550 66162
rect 37550 66110 37602 66162
rect 37602 66110 37604 66162
rect 37548 66108 37604 66110
rect 36428 63810 36484 63812
rect 36428 63758 36430 63810
rect 36430 63758 36482 63810
rect 36482 63758 36484 63810
rect 36428 63756 36484 63758
rect 36316 60732 36372 60788
rect 36316 60562 36372 60564
rect 36316 60510 36318 60562
rect 36318 60510 36370 60562
rect 36370 60510 36372 60562
rect 36316 60508 36372 60510
rect 35980 59500 36036 59556
rect 35644 59218 35700 59220
rect 35644 59166 35646 59218
rect 35646 59166 35698 59218
rect 35698 59166 35700 59218
rect 35644 59164 35700 59166
rect 35980 59106 36036 59108
rect 35980 59054 35982 59106
rect 35982 59054 36034 59106
rect 36034 59054 36036 59106
rect 35980 59052 36036 59054
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35644 56252 35700 56308
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35532 55356 35588 55412
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35756 56588 35812 56644
rect 35756 55074 35812 55076
rect 35756 55022 35758 55074
rect 35758 55022 35810 55074
rect 35810 55022 35812 55074
rect 35756 55020 35812 55022
rect 35532 53340 35588 53396
rect 35644 52892 35700 52948
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34524 50876 34580 50932
rect 34524 50652 34580 50708
rect 34412 48076 34468 48132
rect 34300 47964 34356 48020
rect 34524 46620 34580 46676
rect 34972 51938 35028 51940
rect 34972 51886 34974 51938
rect 34974 51886 35026 51938
rect 35026 51886 35028 51938
rect 34972 51884 35028 51886
rect 35532 51884 35588 51940
rect 35420 51378 35476 51380
rect 35420 51326 35422 51378
rect 35422 51326 35474 51378
rect 35474 51326 35476 51378
rect 35420 51324 35476 51326
rect 35756 51212 35812 51268
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 36428 59218 36484 59220
rect 36428 59166 36430 59218
rect 36430 59166 36482 59218
rect 36482 59166 36484 59218
rect 36428 59164 36484 59166
rect 36316 58940 36372 58996
rect 36652 64034 36708 64036
rect 36652 63982 36654 64034
rect 36654 63982 36706 64034
rect 36706 63982 36708 64034
rect 36652 63980 36708 63982
rect 36876 65436 36932 65492
rect 37660 65490 37716 65492
rect 37660 65438 37662 65490
rect 37662 65438 37714 65490
rect 37714 65438 37716 65490
rect 37660 65436 37716 65438
rect 37548 65324 37604 65380
rect 38444 66108 38500 66164
rect 37884 64818 37940 64820
rect 37884 64766 37886 64818
rect 37886 64766 37938 64818
rect 37938 64766 37940 64818
rect 37884 64764 37940 64766
rect 38668 64764 38724 64820
rect 37884 63756 37940 63812
rect 36764 60898 36820 60900
rect 36764 60846 36766 60898
rect 36766 60846 36818 60898
rect 36818 60846 36820 60898
rect 36764 60844 36820 60846
rect 38780 63922 38836 63924
rect 38780 63870 38782 63922
rect 38782 63870 38834 63922
rect 38834 63870 38836 63922
rect 38780 63868 38836 63870
rect 38220 63644 38276 63700
rect 36876 60956 36932 61012
rect 37772 61458 37828 61460
rect 37772 61406 37774 61458
rect 37774 61406 37826 61458
rect 37826 61406 37828 61458
rect 37772 61404 37828 61406
rect 37100 61180 37156 61236
rect 37212 60732 37268 60788
rect 37100 59836 37156 59892
rect 37324 60508 37380 60564
rect 36764 59052 36820 59108
rect 36652 56194 36708 56196
rect 36652 56142 36654 56194
rect 36654 56142 36706 56194
rect 36706 56142 36708 56194
rect 36652 56140 36708 56142
rect 36876 59218 36932 59220
rect 36876 59166 36878 59218
rect 36878 59166 36930 59218
rect 36930 59166 36932 59218
rect 36876 59164 36932 59166
rect 37212 59218 37268 59220
rect 37212 59166 37214 59218
rect 37214 59166 37266 59218
rect 37266 59166 37268 59218
rect 37212 59164 37268 59166
rect 39004 67058 39060 67060
rect 39004 67006 39006 67058
rect 39006 67006 39058 67058
rect 39058 67006 39060 67058
rect 39004 67004 39060 67006
rect 39116 66332 39172 66388
rect 39228 66274 39284 66276
rect 39228 66222 39230 66274
rect 39230 66222 39282 66274
rect 39282 66222 39284 66274
rect 39228 66220 39284 66222
rect 39564 67004 39620 67060
rect 41356 66386 41412 66388
rect 41356 66334 41358 66386
rect 41358 66334 41410 66386
rect 41410 66334 41412 66386
rect 41356 66332 41412 66334
rect 40124 65996 40180 66052
rect 40012 65212 40068 65268
rect 39788 64146 39844 64148
rect 39788 64094 39790 64146
rect 39790 64094 39842 64146
rect 39842 64094 39844 64146
rect 39788 64092 39844 64094
rect 41020 66050 41076 66052
rect 41020 65998 41022 66050
rect 41022 65998 41074 66050
rect 41074 65998 41076 66050
rect 41020 65996 41076 65998
rect 40572 65324 40628 65380
rect 41916 65772 41972 65828
rect 41020 65324 41076 65380
rect 40348 65212 40404 65268
rect 40908 65266 40964 65268
rect 40908 65214 40910 65266
rect 40910 65214 40962 65266
rect 40962 65214 40964 65266
rect 40908 65212 40964 65214
rect 42252 66332 42308 66388
rect 42588 67004 42644 67060
rect 43372 67058 43428 67060
rect 43372 67006 43374 67058
rect 43374 67006 43426 67058
rect 43426 67006 43428 67058
rect 43372 67004 43428 67006
rect 43260 66780 43316 66836
rect 42364 65772 42420 65828
rect 41356 65324 41412 65380
rect 39900 63868 39956 63924
rect 39004 63810 39060 63812
rect 39004 63758 39006 63810
rect 39006 63758 39058 63810
rect 39058 63758 39060 63810
rect 39004 63756 39060 63758
rect 39676 63698 39732 63700
rect 39676 63646 39678 63698
rect 39678 63646 39730 63698
rect 39730 63646 39732 63698
rect 39676 63644 39732 63646
rect 38668 60284 38724 60340
rect 37884 59948 37940 60004
rect 37660 59890 37716 59892
rect 37660 59838 37662 59890
rect 37662 59838 37714 59890
rect 37714 59838 37716 59890
rect 37660 59836 37716 59838
rect 39116 60060 39172 60116
rect 38108 59218 38164 59220
rect 38108 59166 38110 59218
rect 38110 59166 38162 59218
rect 38162 59166 38164 59218
rect 38108 59164 38164 59166
rect 36988 58940 37044 58996
rect 36988 58156 37044 58212
rect 38556 59052 38612 59108
rect 37996 58156 38052 58212
rect 37324 57372 37380 57428
rect 38332 57372 38388 57428
rect 36204 55020 36260 55076
rect 36316 52946 36372 52948
rect 36316 52894 36318 52946
rect 36318 52894 36370 52946
rect 36370 52894 36372 52946
rect 36316 52892 36372 52894
rect 36316 51266 36372 51268
rect 36316 51214 36318 51266
rect 36318 51214 36370 51266
rect 36370 51214 36372 51266
rect 36316 51212 36372 51214
rect 36316 50652 36372 50708
rect 34860 49586 34916 49588
rect 34860 49534 34862 49586
rect 34862 49534 34914 49586
rect 34914 49534 34916 49586
rect 34860 49532 34916 49534
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34972 48860 35028 48916
rect 34860 48802 34916 48804
rect 34860 48750 34862 48802
rect 34862 48750 34914 48802
rect 34914 48750 34916 48802
rect 34860 48748 34916 48750
rect 35868 49532 35924 49588
rect 35532 48914 35588 48916
rect 35532 48862 35534 48914
rect 35534 48862 35586 48914
rect 35586 48862 35588 48914
rect 35532 48860 35588 48862
rect 35308 48802 35364 48804
rect 35308 48750 35310 48802
rect 35310 48750 35362 48802
rect 35362 48750 35364 48802
rect 35308 48748 35364 48750
rect 35756 48636 35812 48692
rect 34972 48130 35028 48132
rect 34972 48078 34974 48130
rect 34974 48078 35026 48130
rect 35026 48078 35028 48130
rect 34972 48076 35028 48078
rect 34748 47516 34804 47572
rect 34972 47458 35028 47460
rect 34972 47406 34974 47458
rect 34974 47406 35026 47458
rect 35026 47406 35028 47458
rect 34972 47404 35028 47406
rect 35196 47964 35252 48020
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 34748 46674 34804 46676
rect 34748 46622 34750 46674
rect 34750 46622 34802 46674
rect 34802 46622 34804 46674
rect 34748 46620 34804 46622
rect 34636 46396 34692 46452
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 33628 45388 33684 45444
rect 34300 44994 34356 44996
rect 34300 44942 34302 44994
rect 34302 44942 34354 44994
rect 34354 44942 34356 44994
rect 34300 44940 34356 44942
rect 34300 44380 34356 44436
rect 34748 45164 34804 45220
rect 35308 45276 35364 45332
rect 35644 45218 35700 45220
rect 35644 45166 35646 45218
rect 35646 45166 35698 45218
rect 35698 45166 35700 45218
rect 35644 45164 35700 45166
rect 35532 44940 35588 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34412 44322 34468 44324
rect 34412 44270 34414 44322
rect 34414 44270 34466 44322
rect 34466 44270 34468 44322
rect 34412 44268 34468 44270
rect 34972 44322 35028 44324
rect 34972 44270 34974 44322
rect 34974 44270 35026 44322
rect 35026 44270 35028 44322
rect 34972 44268 35028 44270
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 33516 42588 33572 42644
rect 33404 42140 33460 42196
rect 33180 42028 33236 42084
rect 32844 41916 32900 41972
rect 33292 41916 33348 41972
rect 33180 41804 33236 41860
rect 32956 41186 33012 41188
rect 32956 41134 32958 41186
rect 32958 41134 33010 41186
rect 33010 41134 33012 41186
rect 32956 41132 33012 41134
rect 31724 38892 31780 38948
rect 32284 40124 32340 40180
rect 31276 38108 31332 38164
rect 31500 36988 31556 37044
rect 31276 36876 31332 36932
rect 32732 40348 32788 40404
rect 32396 40012 32452 40068
rect 32396 39228 32452 39284
rect 31948 37100 32004 37156
rect 32060 37042 32116 37044
rect 32060 36990 32062 37042
rect 32062 36990 32114 37042
rect 32114 36990 32116 37042
rect 32060 36988 32116 36990
rect 31836 36876 31892 36932
rect 30940 35196 30996 35252
rect 31052 34860 31108 34916
rect 29932 31724 29988 31780
rect 29820 30940 29876 30996
rect 29932 30828 29988 30884
rect 29708 29596 29764 29652
rect 30044 30044 30100 30100
rect 29484 29372 29540 29428
rect 28028 26796 28084 26852
rect 28700 26348 28756 26404
rect 27916 26236 27972 26292
rect 28028 25506 28084 25508
rect 28028 25454 28030 25506
rect 28030 25454 28082 25506
rect 28082 25454 28084 25506
rect 28028 25452 28084 25454
rect 28924 26402 28980 26404
rect 28924 26350 28926 26402
rect 28926 26350 28978 26402
rect 28978 26350 28980 26402
rect 28924 26348 28980 26350
rect 28140 23436 28196 23492
rect 28028 21084 28084 21140
rect 28140 20690 28196 20692
rect 28140 20638 28142 20690
rect 28142 20638 28194 20690
rect 28194 20638 28196 20690
rect 28140 20636 28196 20638
rect 27804 20578 27860 20580
rect 27804 20526 27806 20578
rect 27806 20526 27858 20578
rect 27858 20526 27860 20578
rect 27804 20524 27860 20526
rect 27916 19906 27972 19908
rect 27916 19854 27918 19906
rect 27918 19854 27970 19906
rect 27970 19854 27972 19906
rect 27916 19852 27972 19854
rect 27916 15484 27972 15540
rect 27132 13580 27188 13636
rect 26348 12402 26404 12404
rect 26348 12350 26350 12402
rect 26350 12350 26402 12402
rect 26402 12350 26404 12402
rect 26348 12348 26404 12350
rect 26236 12178 26292 12180
rect 26236 12126 26238 12178
rect 26238 12126 26290 12178
rect 26290 12126 26292 12178
rect 26236 12124 26292 12126
rect 26236 11788 26292 11844
rect 26012 10780 26068 10836
rect 25564 9884 25620 9940
rect 28588 24556 28644 24612
rect 28476 23154 28532 23156
rect 28476 23102 28478 23154
rect 28478 23102 28530 23154
rect 28530 23102 28532 23154
rect 28476 23100 28532 23102
rect 28812 23324 28868 23380
rect 28812 22428 28868 22484
rect 28588 21084 28644 21140
rect 28588 20636 28644 20692
rect 28700 19292 28756 19348
rect 28812 18450 28868 18452
rect 28812 18398 28814 18450
rect 28814 18398 28866 18450
rect 28866 18398 28868 18450
rect 28812 18396 28868 18398
rect 28588 17106 28644 17108
rect 28588 17054 28590 17106
rect 28590 17054 28642 17106
rect 28642 17054 28644 17106
rect 28588 17052 28644 17054
rect 27804 12290 27860 12292
rect 27804 12238 27806 12290
rect 27806 12238 27858 12290
rect 27858 12238 27860 12290
rect 27804 12236 27860 12238
rect 27468 12178 27524 12180
rect 27468 12126 27470 12178
rect 27470 12126 27522 12178
rect 27522 12126 27524 12178
rect 27468 12124 27524 12126
rect 26236 7756 26292 7812
rect 25788 7474 25844 7476
rect 25788 7422 25790 7474
rect 25790 7422 25842 7474
rect 25842 7422 25844 7474
rect 25788 7420 25844 7422
rect 25228 6860 25284 6916
rect 26460 10108 26516 10164
rect 27020 10332 27076 10388
rect 27020 9714 27076 9716
rect 27020 9662 27022 9714
rect 27022 9662 27074 9714
rect 27074 9662 27076 9714
rect 27020 9660 27076 9662
rect 26908 7868 26964 7924
rect 26908 6860 26964 6916
rect 26572 6076 26628 6132
rect 25004 5346 25060 5348
rect 25004 5294 25006 5346
rect 25006 5294 25058 5346
rect 25058 5294 25060 5346
rect 25004 5292 25060 5294
rect 25340 5180 25396 5236
rect 26012 5234 26068 5236
rect 26012 5182 26014 5234
rect 26014 5182 26066 5234
rect 26066 5182 26068 5234
rect 26012 5180 26068 5182
rect 25340 4956 25396 5012
rect 25900 4284 25956 4340
rect 27356 10108 27412 10164
rect 27692 10332 27748 10388
rect 27580 9714 27636 9716
rect 27580 9662 27582 9714
rect 27582 9662 27634 9714
rect 27634 9662 27636 9714
rect 27580 9660 27636 9662
rect 28252 12348 28308 12404
rect 29148 26290 29204 26292
rect 29148 26238 29150 26290
rect 29150 26238 29202 26290
rect 29202 26238 29204 26290
rect 29148 26236 29204 26238
rect 29036 25452 29092 25508
rect 29596 29260 29652 29316
rect 29148 24668 29204 24724
rect 30156 29260 30212 29316
rect 29708 27970 29764 27972
rect 29708 27918 29710 27970
rect 29710 27918 29762 27970
rect 29762 27918 29764 27970
rect 29708 27916 29764 27918
rect 29148 23154 29204 23156
rect 29148 23102 29150 23154
rect 29150 23102 29202 23154
rect 29202 23102 29204 23154
rect 29148 23100 29204 23102
rect 29708 27692 29764 27748
rect 30268 27580 30324 27636
rect 29708 24220 29764 24276
rect 30716 31778 30772 31780
rect 30716 31726 30718 31778
rect 30718 31726 30770 31778
rect 30770 31726 30772 31778
rect 30716 31724 30772 31726
rect 30828 30994 30884 30996
rect 30828 30942 30830 30994
rect 30830 30942 30882 30994
rect 30882 30942 30884 30994
rect 30828 30940 30884 30942
rect 30828 28364 30884 28420
rect 30604 27746 30660 27748
rect 30604 27694 30606 27746
rect 30606 27694 30658 27746
rect 30658 27694 30660 27746
rect 30604 27692 30660 27694
rect 29596 23660 29652 23716
rect 29372 22652 29428 22708
rect 29260 22482 29316 22484
rect 29260 22430 29262 22482
rect 29262 22430 29314 22482
rect 29314 22430 29316 22482
rect 29260 22428 29316 22430
rect 29036 19906 29092 19908
rect 29036 19854 29038 19906
rect 29038 19854 29090 19906
rect 29090 19854 29092 19906
rect 29036 19852 29092 19854
rect 28924 14588 28980 14644
rect 29372 17778 29428 17780
rect 29372 17726 29374 17778
rect 29374 17726 29426 17778
rect 29426 17726 29428 17778
rect 29372 17724 29428 17726
rect 29372 16828 29428 16884
rect 29932 23324 29988 23380
rect 29708 21586 29764 21588
rect 29708 21534 29710 21586
rect 29710 21534 29762 21586
rect 29762 21534 29764 21586
rect 29708 21532 29764 21534
rect 30268 21586 30324 21588
rect 30268 21534 30270 21586
rect 30270 21534 30322 21586
rect 30322 21534 30324 21586
rect 30268 21532 30324 21534
rect 30828 26852 30884 26908
rect 31052 32562 31108 32564
rect 31052 32510 31054 32562
rect 31054 32510 31106 32562
rect 31106 32510 31108 32562
rect 31052 32508 31108 32510
rect 30940 26684 30996 26740
rect 31164 26572 31220 26628
rect 31836 35084 31892 35140
rect 32060 35196 32116 35252
rect 31836 34914 31892 34916
rect 31836 34862 31838 34914
rect 31838 34862 31890 34914
rect 31890 34862 31892 34914
rect 31836 34860 31892 34862
rect 32060 33068 32116 33124
rect 32060 32562 32116 32564
rect 32060 32510 32062 32562
rect 32062 32510 32114 32562
rect 32114 32510 32116 32562
rect 32060 32508 32116 32510
rect 31724 31890 31780 31892
rect 31724 31838 31726 31890
rect 31726 31838 31778 31890
rect 31778 31838 31780 31890
rect 31724 31836 31780 31838
rect 31612 31724 31668 31780
rect 31500 31276 31556 31332
rect 31948 31164 32004 31220
rect 31388 30940 31444 30996
rect 31948 30828 32004 30884
rect 32060 30716 32116 30772
rect 31948 29426 32004 29428
rect 31948 29374 31950 29426
rect 31950 29374 32002 29426
rect 32002 29374 32004 29426
rect 31948 29372 32004 29374
rect 31612 28476 31668 28532
rect 31948 28476 32004 28532
rect 31276 26348 31332 26404
rect 31388 27692 31444 27748
rect 31612 27580 31668 27636
rect 32060 28364 32116 28420
rect 32060 28028 32116 28084
rect 31500 26908 31556 26964
rect 31724 26796 31780 26852
rect 31612 26236 31668 26292
rect 30044 20748 30100 20804
rect 30716 20748 30772 20804
rect 30156 19964 30212 20020
rect 30828 20076 30884 20132
rect 29932 18338 29988 18340
rect 29932 18286 29934 18338
rect 29934 18286 29986 18338
rect 29986 18286 29988 18338
rect 29932 18284 29988 18286
rect 29932 17442 29988 17444
rect 29932 17390 29934 17442
rect 29934 17390 29986 17442
rect 29986 17390 29988 17442
rect 29932 17388 29988 17390
rect 29932 16882 29988 16884
rect 29932 16830 29934 16882
rect 29934 16830 29986 16882
rect 29986 16830 29988 16882
rect 29932 16828 29988 16830
rect 30492 17442 30548 17444
rect 30492 17390 30494 17442
rect 30494 17390 30546 17442
rect 30546 17390 30548 17442
rect 30492 17388 30548 17390
rect 29708 16156 29764 16212
rect 29820 16098 29876 16100
rect 29820 16046 29822 16098
rect 29822 16046 29874 16098
rect 29874 16046 29876 16098
rect 29820 16044 29876 16046
rect 29820 15596 29876 15652
rect 29596 15036 29652 15092
rect 29260 14588 29316 14644
rect 29148 14028 29204 14084
rect 28476 12124 28532 12180
rect 28252 11340 28308 11396
rect 29148 11452 29204 11508
rect 28028 11282 28084 11284
rect 28028 11230 28030 11282
rect 28030 11230 28082 11282
rect 28082 11230 28084 11282
rect 28028 11228 28084 11230
rect 28588 11282 28644 11284
rect 28588 11230 28590 11282
rect 28590 11230 28642 11282
rect 28642 11230 28644 11282
rect 28588 11228 28644 11230
rect 29708 14642 29764 14644
rect 29708 14590 29710 14642
rect 29710 14590 29762 14642
rect 29762 14590 29764 14642
rect 29708 14588 29764 14590
rect 29932 15372 29988 15428
rect 29820 11506 29876 11508
rect 29820 11454 29822 11506
rect 29822 11454 29874 11506
rect 29874 11454 29876 11506
rect 29820 11452 29876 11454
rect 29260 11282 29316 11284
rect 29260 11230 29262 11282
rect 29262 11230 29314 11282
rect 29314 11230 29316 11282
rect 29260 11228 29316 11230
rect 30156 15036 30212 15092
rect 30716 16156 30772 16212
rect 30380 16098 30436 16100
rect 30380 16046 30382 16098
rect 30382 16046 30434 16098
rect 30434 16046 30436 16098
rect 30380 16044 30436 16046
rect 30492 15036 30548 15092
rect 30492 14700 30548 14756
rect 30604 14588 30660 14644
rect 30492 13858 30548 13860
rect 30492 13806 30494 13858
rect 30494 13806 30546 13858
rect 30546 13806 30548 13858
rect 30492 13804 30548 13806
rect 29484 9996 29540 10052
rect 28476 8988 28532 9044
rect 27132 7756 27188 7812
rect 27468 7868 27524 7924
rect 27916 8034 27972 8036
rect 27916 7982 27918 8034
rect 27918 7982 27970 8034
rect 27970 7982 27972 8034
rect 27916 7980 27972 7982
rect 27804 7756 27860 7812
rect 28028 7644 28084 7700
rect 28252 7868 28308 7924
rect 27356 6860 27412 6916
rect 28700 7698 28756 7700
rect 28700 7646 28702 7698
rect 28702 7646 28754 7698
rect 28754 7646 28756 7698
rect 28700 7644 28756 7646
rect 30940 19852 30996 19908
rect 30940 17836 30996 17892
rect 30828 12962 30884 12964
rect 30828 12910 30830 12962
rect 30830 12910 30882 12962
rect 30882 12910 30884 12962
rect 30828 12908 30884 12910
rect 30268 11282 30324 11284
rect 30268 11230 30270 11282
rect 30270 11230 30322 11282
rect 30322 11230 30324 11282
rect 30268 11228 30324 11230
rect 29820 7084 29876 7140
rect 28700 5292 28756 5348
rect 29820 6300 29876 6356
rect 30268 7084 30324 7140
rect 29372 5068 29428 5124
rect 30044 5068 30100 5124
rect 28028 4844 28084 4900
rect 29932 4450 29988 4452
rect 29932 4398 29934 4450
rect 29934 4398 29986 4450
rect 29986 4398 29988 4450
rect 29932 4396 29988 4398
rect 27468 4338 27524 4340
rect 27468 4286 27470 4338
rect 27470 4286 27522 4338
rect 27522 4286 27524 4338
rect 27468 4284 27524 4286
rect 30380 6300 30436 6356
rect 30716 9996 30772 10052
rect 31612 23884 31668 23940
rect 32060 27020 32116 27076
rect 32620 39618 32676 39620
rect 32620 39566 32622 39618
rect 32622 39566 32674 39618
rect 32674 39566 32676 39618
rect 32620 39564 32676 39566
rect 32620 36988 32676 37044
rect 32732 35644 32788 35700
rect 32732 29372 32788 29428
rect 32620 28530 32676 28532
rect 32620 28478 32622 28530
rect 32622 28478 32674 28530
rect 32674 28478 32676 28530
rect 32620 28476 32676 28478
rect 33180 40572 33236 40628
rect 33180 40348 33236 40404
rect 32956 36540 33012 36596
rect 33964 42642 34020 42644
rect 33964 42590 33966 42642
rect 33966 42590 34018 42642
rect 34018 42590 34020 42642
rect 33964 42588 34020 42590
rect 33852 42082 33908 42084
rect 33852 42030 33854 42082
rect 33854 42030 33906 42082
rect 33906 42030 33908 42082
rect 33852 42028 33908 42030
rect 34412 42082 34468 42084
rect 34412 42030 34414 42082
rect 34414 42030 34466 42082
rect 34466 42030 34468 42082
rect 34412 42028 34468 42030
rect 35420 41970 35476 41972
rect 35420 41918 35422 41970
rect 35422 41918 35474 41970
rect 35474 41918 35476 41970
rect 35420 41916 35476 41918
rect 34300 41804 34356 41860
rect 34412 41746 34468 41748
rect 34412 41694 34414 41746
rect 34414 41694 34466 41746
rect 34466 41694 34468 41746
rect 34412 41692 34468 41694
rect 35532 41692 35588 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 33964 41186 34020 41188
rect 33964 41134 33966 41186
rect 33966 41134 34018 41186
rect 34018 41134 34020 41186
rect 33964 41132 34020 41134
rect 33516 40796 33572 40852
rect 33740 41074 33796 41076
rect 33740 41022 33742 41074
rect 33742 41022 33794 41074
rect 33794 41022 33796 41074
rect 33740 41020 33796 41022
rect 33516 39618 33572 39620
rect 33516 39566 33518 39618
rect 33518 39566 33570 39618
rect 33570 39566 33572 39618
rect 33516 39564 33572 39566
rect 33292 35756 33348 35812
rect 35084 41356 35140 41412
rect 34972 41244 35028 41300
rect 34524 41132 34580 41188
rect 34748 40962 34804 40964
rect 34748 40910 34750 40962
rect 34750 40910 34802 40962
rect 34802 40910 34804 40962
rect 34748 40908 34804 40910
rect 33740 34188 33796 34244
rect 34188 38892 34244 38948
rect 34188 34860 34244 34916
rect 35868 48130 35924 48132
rect 35868 48078 35870 48130
rect 35870 48078 35922 48130
rect 35922 48078 35924 48130
rect 35868 48076 35924 48078
rect 35868 45218 35924 45220
rect 35868 45166 35870 45218
rect 35870 45166 35922 45218
rect 35922 45166 35924 45218
rect 35868 45164 35924 45166
rect 36428 48300 36484 48356
rect 36204 45218 36260 45220
rect 36204 45166 36206 45218
rect 36206 45166 36258 45218
rect 36258 45166 36260 45218
rect 36204 45164 36260 45166
rect 36092 43932 36148 43988
rect 36092 41970 36148 41972
rect 36092 41918 36094 41970
rect 36094 41918 36146 41970
rect 36146 41918 36148 41970
rect 36092 41916 36148 41918
rect 37100 56642 37156 56644
rect 37100 56590 37102 56642
rect 37102 56590 37154 56642
rect 37154 56590 37156 56642
rect 37100 56588 37156 56590
rect 37100 56306 37156 56308
rect 37100 56254 37102 56306
rect 37102 56254 37154 56306
rect 37154 56254 37156 56306
rect 37100 56252 37156 56254
rect 37212 56194 37268 56196
rect 37212 56142 37214 56194
rect 37214 56142 37266 56194
rect 37266 56142 37268 56194
rect 37212 56140 37268 56142
rect 37436 54012 37492 54068
rect 37436 52892 37492 52948
rect 37212 52220 37268 52276
rect 37884 54012 37940 54068
rect 38332 54012 38388 54068
rect 37996 52274 38052 52276
rect 37996 52222 37998 52274
rect 37998 52222 38050 52274
rect 38050 52222 38052 52274
rect 37996 52220 38052 52222
rect 36876 48748 36932 48804
rect 37212 48300 37268 48356
rect 37100 48130 37156 48132
rect 37100 48078 37102 48130
rect 37102 48078 37154 48130
rect 37154 48078 37156 48130
rect 37100 48076 37156 48078
rect 36876 45612 36932 45668
rect 36764 45388 36820 45444
rect 37324 45276 37380 45332
rect 36428 44268 36484 44324
rect 36316 42252 36372 42308
rect 35084 40572 35140 40628
rect 35420 41020 35476 41076
rect 34412 40236 34468 40292
rect 34636 40236 34692 40292
rect 35532 40348 35588 40404
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34412 39228 34468 39284
rect 35084 39676 35140 39732
rect 35084 39228 35140 39284
rect 34748 38780 34804 38836
rect 34972 38892 35028 38948
rect 34972 37378 35028 37380
rect 34972 37326 34974 37378
rect 34974 37326 35026 37378
rect 35026 37326 35028 37378
rect 34972 37324 35028 37326
rect 34748 37266 34804 37268
rect 34748 37214 34750 37266
rect 34750 37214 34802 37266
rect 34802 37214 34804 37266
rect 34748 37212 34804 37214
rect 34412 35756 34468 35812
rect 34860 35644 34916 35700
rect 34748 34690 34804 34692
rect 34748 34638 34750 34690
rect 34750 34638 34802 34690
rect 34802 34638 34804 34690
rect 34748 34636 34804 34638
rect 34188 32732 34244 32788
rect 32956 31836 33012 31892
rect 33292 30716 33348 30772
rect 33852 29932 33908 29988
rect 33180 27634 33236 27636
rect 33180 27582 33182 27634
rect 33182 27582 33234 27634
rect 33234 27582 33236 27634
rect 33180 27580 33236 27582
rect 32732 27244 32788 27300
rect 31836 24892 31892 24948
rect 31948 23938 32004 23940
rect 31948 23886 31950 23938
rect 31950 23886 32002 23938
rect 32002 23886 32004 23938
rect 31948 23884 32004 23886
rect 31724 20860 31780 20916
rect 31612 20188 31668 20244
rect 31164 20076 31220 20132
rect 31500 20130 31556 20132
rect 31500 20078 31502 20130
rect 31502 20078 31554 20130
rect 31554 20078 31556 20130
rect 31500 20076 31556 20078
rect 31388 20018 31444 20020
rect 31388 19966 31390 20018
rect 31390 19966 31442 20018
rect 31442 19966 31444 20018
rect 31388 19964 31444 19966
rect 31948 20188 32004 20244
rect 32284 20860 32340 20916
rect 32396 20188 32452 20244
rect 32620 26236 32676 26292
rect 32844 27020 32900 27076
rect 33068 27020 33124 27076
rect 33628 27020 33684 27076
rect 33964 29820 34020 29876
rect 33516 26460 33572 26516
rect 32620 20914 32676 20916
rect 32620 20862 32622 20914
rect 32622 20862 32674 20914
rect 32674 20862 32676 20914
rect 32620 20860 32676 20862
rect 31164 18732 31220 18788
rect 31948 18732 32004 18788
rect 31164 17724 31220 17780
rect 31724 18562 31780 18564
rect 31724 18510 31726 18562
rect 31726 18510 31778 18562
rect 31778 18510 31780 18562
rect 31724 18508 31780 18510
rect 31724 17778 31780 17780
rect 31724 17726 31726 17778
rect 31726 17726 31778 17778
rect 31778 17726 31780 17778
rect 31724 17724 31780 17726
rect 31164 17442 31220 17444
rect 31164 17390 31166 17442
rect 31166 17390 31218 17442
rect 31218 17390 31220 17442
rect 31164 17388 31220 17390
rect 31164 16828 31220 16884
rect 31276 16210 31332 16212
rect 31276 16158 31278 16210
rect 31278 16158 31330 16210
rect 31330 16158 31332 16210
rect 31276 16156 31332 16158
rect 32060 16882 32116 16884
rect 32060 16830 32062 16882
rect 32062 16830 32114 16882
rect 32114 16830 32116 16882
rect 32060 16828 32116 16830
rect 32284 17724 32340 17780
rect 32060 16098 32116 16100
rect 32060 16046 32062 16098
rect 32062 16046 32114 16098
rect 32114 16046 32116 16098
rect 32060 16044 32116 16046
rect 31052 14588 31108 14644
rect 31052 13804 31108 13860
rect 31836 13916 31892 13972
rect 32060 14700 32116 14756
rect 33068 23714 33124 23716
rect 33068 23662 33070 23714
rect 33070 23662 33122 23714
rect 33122 23662 33124 23714
rect 33068 23660 33124 23662
rect 33852 26236 33908 26292
rect 33964 24892 34020 24948
rect 33516 24668 33572 24724
rect 33292 20748 33348 20804
rect 33068 20076 33124 20132
rect 33068 19292 33124 19348
rect 33292 20188 33348 20244
rect 33964 24722 34020 24724
rect 33964 24670 33966 24722
rect 33966 24670 34018 24722
rect 34018 24670 34020 24722
rect 33964 24668 34020 24670
rect 33964 23660 34020 23716
rect 34076 23772 34132 23828
rect 33852 23212 33908 23268
rect 33852 22988 33908 23044
rect 34076 23042 34132 23044
rect 34076 22990 34078 23042
rect 34078 22990 34130 23042
rect 34130 22990 34132 23042
rect 34076 22988 34132 22990
rect 33740 20860 33796 20916
rect 33852 20972 33908 21028
rect 33740 19346 33796 19348
rect 33740 19294 33742 19346
rect 33742 19294 33794 19346
rect 33794 19294 33796 19346
rect 33740 19292 33796 19294
rect 33628 19234 33684 19236
rect 33628 19182 33630 19234
rect 33630 19182 33682 19234
rect 33682 19182 33684 19234
rect 33628 19180 33684 19182
rect 34412 33964 34468 34020
rect 34636 34242 34692 34244
rect 34636 34190 34638 34242
rect 34638 34190 34690 34242
rect 34690 34190 34692 34242
rect 34636 34188 34692 34190
rect 34860 33906 34916 33908
rect 34860 33854 34862 33906
rect 34862 33854 34914 33906
rect 34914 33854 34916 33906
rect 34860 33852 34916 33854
rect 34748 32508 34804 32564
rect 34972 32786 35028 32788
rect 34972 32734 34974 32786
rect 34974 32734 35026 32786
rect 35026 32734 35028 32786
rect 34972 32732 35028 32734
rect 34412 31836 34468 31892
rect 34524 31724 34580 31780
rect 34636 31612 34692 31668
rect 34748 30156 34804 30212
rect 34524 30044 34580 30100
rect 35756 41186 35812 41188
rect 35756 41134 35758 41186
rect 35758 41134 35810 41186
rect 35810 41134 35812 41186
rect 35756 41132 35812 41134
rect 35980 39730 36036 39732
rect 35980 39678 35982 39730
rect 35982 39678 36034 39730
rect 36034 39678 36036 39730
rect 35980 39676 36036 39678
rect 35868 39116 35924 39172
rect 35196 38834 35252 38836
rect 35196 38782 35198 38834
rect 35198 38782 35250 38834
rect 35250 38782 35252 38834
rect 35196 38780 35252 38782
rect 35868 38668 35924 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35532 35756 35588 35812
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36204 41356 36260 41412
rect 36316 41074 36372 41076
rect 36316 41022 36318 41074
rect 36318 41022 36370 41074
rect 36370 41022 36372 41074
rect 36316 41020 36372 41022
rect 36204 40962 36260 40964
rect 36204 40910 36206 40962
rect 36206 40910 36258 40962
rect 36258 40910 36260 40962
rect 36204 40908 36260 40910
rect 36092 38668 36148 38724
rect 36428 39116 36484 39172
rect 36092 38444 36148 38500
rect 35196 34860 35252 34916
rect 35308 34300 35364 34356
rect 35532 34412 35588 34468
rect 35532 34188 35588 34244
rect 35868 34242 35924 34244
rect 35868 34190 35870 34242
rect 35870 34190 35922 34242
rect 35922 34190 35924 34242
rect 35868 34188 35924 34190
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35756 33852 35812 33908
rect 36204 34636 36260 34692
rect 35644 31890 35700 31892
rect 35644 31838 35646 31890
rect 35646 31838 35698 31890
rect 35698 31838 35700 31890
rect 35644 31836 35700 31838
rect 35532 31778 35588 31780
rect 35532 31726 35534 31778
rect 35534 31726 35586 31778
rect 35586 31726 35588 31778
rect 35532 31724 35588 31726
rect 35980 31666 36036 31668
rect 35980 31614 35982 31666
rect 35982 31614 36034 31666
rect 36034 31614 36036 31666
rect 35980 31612 36036 31614
rect 35308 30770 35364 30772
rect 35308 30718 35310 30770
rect 35310 30718 35362 30770
rect 35362 30718 35364 30770
rect 35308 30716 35364 30718
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35420 30210 35476 30212
rect 35420 30158 35422 30210
rect 35422 30158 35474 30210
rect 35474 30158 35476 30210
rect 35420 30156 35476 30158
rect 36204 30156 36260 30212
rect 35084 29596 35140 29652
rect 35868 30098 35924 30100
rect 35868 30046 35870 30098
rect 35870 30046 35922 30098
rect 35922 30046 35924 30098
rect 35868 30044 35924 30046
rect 35980 29986 36036 29988
rect 35980 29934 35982 29986
rect 35982 29934 36034 29986
rect 36034 29934 36036 29986
rect 35980 29932 36036 29934
rect 36204 29932 36260 29988
rect 37100 44322 37156 44324
rect 37100 44270 37102 44322
rect 37102 44270 37154 44322
rect 37154 44270 37156 44322
rect 37100 44268 37156 44270
rect 37548 46172 37604 46228
rect 38108 50428 38164 50484
rect 37884 48354 37940 48356
rect 37884 48302 37886 48354
rect 37886 48302 37938 48354
rect 37938 48302 37940 48354
rect 37884 48300 37940 48302
rect 37996 48076 38052 48132
rect 39004 59106 39060 59108
rect 39004 59054 39006 59106
rect 39006 59054 39058 59106
rect 39058 59054 39060 59106
rect 39004 59052 39060 59054
rect 38668 58940 38724 58996
rect 39228 58210 39284 58212
rect 39228 58158 39230 58210
rect 39230 58158 39282 58210
rect 39282 58158 39284 58210
rect 39228 58156 39284 58158
rect 39228 57650 39284 57652
rect 39228 57598 39230 57650
rect 39230 57598 39282 57650
rect 39282 57598 39284 57650
rect 39228 57596 39284 57598
rect 38892 56140 38948 56196
rect 40684 64092 40740 64148
rect 41020 64540 41076 64596
rect 41020 63644 41076 63700
rect 42812 62914 42868 62916
rect 42812 62862 42814 62914
rect 42814 62862 42866 62914
rect 42866 62862 42868 62914
rect 42812 62860 42868 62862
rect 45500 73948 45556 74004
rect 44268 66834 44324 66836
rect 44268 66782 44270 66834
rect 44270 66782 44322 66834
rect 44322 66782 44324 66834
rect 44268 66780 44324 66782
rect 43484 63756 43540 63812
rect 44268 63698 44324 63700
rect 44268 63646 44270 63698
rect 44270 63646 44322 63698
rect 44322 63646 44324 63698
rect 44268 63644 44324 63646
rect 43260 62412 43316 62468
rect 41020 61570 41076 61572
rect 41020 61518 41022 61570
rect 41022 61518 41074 61570
rect 41074 61518 41076 61570
rect 41020 61516 41076 61518
rect 39452 61404 39508 61460
rect 41020 61010 41076 61012
rect 41020 60958 41022 61010
rect 41022 60958 41074 61010
rect 41074 60958 41076 61010
rect 41020 60956 41076 60958
rect 40012 60732 40068 60788
rect 39564 60114 39620 60116
rect 39564 60062 39566 60114
rect 39566 60062 39618 60114
rect 39618 60062 39620 60114
rect 39564 60060 39620 60062
rect 39788 60284 39844 60340
rect 41132 60786 41188 60788
rect 41132 60734 41134 60786
rect 41134 60734 41186 60786
rect 41186 60734 41188 60786
rect 41132 60732 41188 60734
rect 40348 60508 40404 60564
rect 39900 59106 39956 59108
rect 39900 59054 39902 59106
rect 39902 59054 39954 59106
rect 39954 59054 39956 59106
rect 39900 59052 39956 59054
rect 40124 58322 40180 58324
rect 40124 58270 40126 58322
rect 40126 58270 40178 58322
rect 40178 58270 40180 58322
rect 40124 58268 40180 58270
rect 39564 58156 39620 58212
rect 40012 58210 40068 58212
rect 40012 58158 40014 58210
rect 40014 58158 40066 58210
rect 40066 58158 40068 58210
rect 40012 58156 40068 58158
rect 39676 57650 39732 57652
rect 39676 57598 39678 57650
rect 39678 57598 39730 57650
rect 39730 57598 39732 57650
rect 39676 57596 39732 57598
rect 39788 56140 39844 56196
rect 39228 54236 39284 54292
rect 38780 54124 38836 54180
rect 39116 52780 39172 52836
rect 39564 52668 39620 52724
rect 38892 51602 38948 51604
rect 38892 51550 38894 51602
rect 38894 51550 38946 51602
rect 38946 51550 38948 51602
rect 38892 51548 38948 51550
rect 38668 51100 38724 51156
rect 38332 50594 38388 50596
rect 38332 50542 38334 50594
rect 38334 50542 38386 50594
rect 38386 50542 38388 50594
rect 38332 50540 38388 50542
rect 38892 50428 38948 50484
rect 39452 50652 39508 50708
rect 38668 48972 38724 49028
rect 38668 48300 38724 48356
rect 38556 48130 38612 48132
rect 38556 48078 38558 48130
rect 38558 48078 38610 48130
rect 38610 48078 38612 48130
rect 38556 48076 38612 48078
rect 37436 44940 37492 44996
rect 38108 47180 38164 47236
rect 37772 45500 37828 45556
rect 37772 44828 37828 44884
rect 37884 44940 37940 44996
rect 37772 44604 37828 44660
rect 37772 43708 37828 43764
rect 37996 44828 38052 44884
rect 38108 44604 38164 44660
rect 38444 47234 38500 47236
rect 38444 47182 38446 47234
rect 38446 47182 38498 47234
rect 38498 47182 38500 47234
rect 38444 47180 38500 47182
rect 38332 45052 38388 45108
rect 38444 44604 38500 44660
rect 37996 44492 38052 44548
rect 37884 44268 37940 44324
rect 37996 43708 38052 43764
rect 36652 42252 36708 42308
rect 36764 42082 36820 42084
rect 36764 42030 36766 42082
rect 36766 42030 36818 42082
rect 36818 42030 36820 42082
rect 36764 42028 36820 42030
rect 37436 42476 37492 42532
rect 37324 41244 37380 41300
rect 37436 41970 37492 41972
rect 37436 41918 37438 41970
rect 37438 41918 37490 41970
rect 37490 41918 37492 41970
rect 37436 41916 37492 41918
rect 37436 40402 37492 40404
rect 37436 40350 37438 40402
rect 37438 40350 37490 40402
rect 37490 40350 37492 40402
rect 37436 40348 37492 40350
rect 37548 40236 37604 40292
rect 37324 38780 37380 38836
rect 36428 36876 36484 36932
rect 36540 32620 36596 32676
rect 36428 32508 36484 32564
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28812 35140 28868
rect 35308 28812 35364 28868
rect 34972 28476 35028 28532
rect 35196 28530 35252 28532
rect 35196 28478 35198 28530
rect 35198 28478 35250 28530
rect 35250 28478 35252 28530
rect 35196 28476 35252 28478
rect 35420 28588 35476 28644
rect 35308 27916 35364 27972
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35308 27298 35364 27300
rect 35308 27246 35310 27298
rect 35310 27246 35362 27298
rect 35362 27246 35364 27298
rect 35308 27244 35364 27246
rect 35980 28588 36036 28644
rect 35868 28530 35924 28532
rect 35868 28478 35870 28530
rect 35870 28478 35922 28530
rect 35922 28478 35924 28530
rect 35868 28476 35924 28478
rect 35868 27916 35924 27972
rect 35644 27580 35700 27636
rect 34300 20300 34356 20356
rect 36092 27580 36148 27636
rect 32844 16098 32900 16100
rect 32844 16046 32846 16098
rect 32846 16046 32898 16098
rect 32898 16046 32900 16098
rect 32844 16044 32900 16046
rect 32396 14252 32452 14308
rect 32284 13970 32340 13972
rect 32284 13918 32286 13970
rect 32286 13918 32338 13970
rect 32338 13918 32340 13970
rect 32284 13916 32340 13918
rect 32060 12908 32116 12964
rect 33292 14588 33348 14644
rect 32732 14418 32788 14420
rect 32732 14366 32734 14418
rect 32734 14366 32786 14418
rect 32786 14366 32788 14418
rect 32732 14364 32788 14366
rect 32956 11394 33012 11396
rect 32956 11342 32958 11394
rect 32958 11342 33010 11394
rect 33010 11342 33012 11394
rect 32956 11340 33012 11342
rect 33292 11452 33348 11508
rect 34748 26572 34804 26628
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34972 22988 35028 23044
rect 35308 23042 35364 23044
rect 35308 22990 35310 23042
rect 35310 22990 35362 23042
rect 35362 22990 35364 23042
rect 35308 22988 35364 22990
rect 35532 23266 35588 23268
rect 35532 23214 35534 23266
rect 35534 23214 35586 23266
rect 35586 23214 35588 23266
rect 35532 23212 35588 23214
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34748 20188 34804 20244
rect 34860 20300 34916 20356
rect 33628 17106 33684 17108
rect 33628 17054 33630 17106
rect 33630 17054 33682 17106
rect 33682 17054 33684 17106
rect 33628 17052 33684 17054
rect 31164 9154 31220 9156
rect 31164 9102 31166 9154
rect 31166 9102 31218 9154
rect 31218 9102 31220 9154
rect 31164 9100 31220 9102
rect 31724 9100 31780 9156
rect 31612 7420 31668 7476
rect 31276 6690 31332 6692
rect 31276 6638 31278 6690
rect 31278 6638 31330 6690
rect 31330 6638 31332 6690
rect 31276 6636 31332 6638
rect 31388 6578 31444 6580
rect 31388 6526 31390 6578
rect 31390 6526 31442 6578
rect 31442 6526 31444 6578
rect 31388 6524 31444 6526
rect 30604 5122 30660 5124
rect 30604 5070 30606 5122
rect 30606 5070 30658 5122
rect 30658 5070 30660 5122
rect 30604 5068 30660 5070
rect 30492 4450 30548 4452
rect 30492 4398 30494 4450
rect 30494 4398 30546 4450
rect 30546 4398 30548 4450
rect 30492 4396 30548 4398
rect 30604 4338 30660 4340
rect 30604 4286 30606 4338
rect 30606 4286 30658 4338
rect 30658 4286 30660 4338
rect 30604 4284 30660 4286
rect 32956 7474 33012 7476
rect 32956 7422 32958 7474
rect 32958 7422 33010 7474
rect 33010 7422 33012 7474
rect 32956 7420 33012 7422
rect 32396 6690 32452 6692
rect 32396 6638 32398 6690
rect 32398 6638 32450 6690
rect 32450 6638 32452 6690
rect 32396 6636 32452 6638
rect 34188 17106 34244 17108
rect 34188 17054 34190 17106
rect 34190 17054 34242 17106
rect 34242 17054 34244 17106
rect 34188 17052 34244 17054
rect 34524 16940 34580 16996
rect 35196 20300 35252 20356
rect 35084 19852 35140 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35868 24610 35924 24612
rect 35868 24558 35870 24610
rect 35870 24558 35922 24610
rect 35922 24558 35924 24610
rect 35868 24556 35924 24558
rect 36092 20300 36148 20356
rect 36428 20188 36484 20244
rect 35084 19180 35140 19236
rect 35980 19234 36036 19236
rect 35980 19182 35982 19234
rect 35982 19182 36034 19234
rect 36034 19182 36036 19234
rect 35980 19180 36036 19182
rect 36316 19906 36372 19908
rect 36316 19854 36318 19906
rect 36318 19854 36370 19906
rect 36370 19854 36372 19906
rect 36316 19852 36372 19854
rect 36652 19852 36708 19908
rect 36204 19346 36260 19348
rect 36204 19294 36206 19346
rect 36206 19294 36258 19346
rect 36258 19294 36260 19346
rect 36204 19292 36260 19294
rect 36316 19180 36372 19236
rect 36652 18562 36708 18564
rect 36652 18510 36654 18562
rect 36654 18510 36706 18562
rect 36706 18510 36708 18562
rect 36652 18508 36708 18510
rect 36540 18396 36596 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36204 17554 36260 17556
rect 36204 17502 36206 17554
rect 36206 17502 36258 17554
rect 36258 17502 36260 17554
rect 36204 17500 36260 17502
rect 35980 16940 36036 16996
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35980 16492 36036 16548
rect 37100 34690 37156 34692
rect 37100 34638 37102 34690
rect 37102 34638 37154 34690
rect 37154 34638 37156 34690
rect 37100 34636 37156 34638
rect 37100 33458 37156 33460
rect 37100 33406 37102 33458
rect 37102 33406 37154 33458
rect 37154 33406 37156 33458
rect 37100 33404 37156 33406
rect 37436 35420 37492 35476
rect 39116 48748 39172 48804
rect 39004 47516 39060 47572
rect 38892 47292 38948 47348
rect 38780 47068 38836 47124
rect 38668 45388 38724 45444
rect 38668 44940 38724 44996
rect 38668 44604 38724 44660
rect 38668 44322 38724 44324
rect 38668 44270 38670 44322
rect 38670 44270 38722 44322
rect 38722 44270 38724 44322
rect 38668 44268 38724 44270
rect 38108 42476 38164 42532
rect 38220 40236 38276 40292
rect 37996 38780 38052 38836
rect 38668 43260 38724 43316
rect 38444 42028 38500 42084
rect 38556 41804 38612 41860
rect 38556 40908 38612 40964
rect 39004 43372 39060 43428
rect 39004 42530 39060 42532
rect 39004 42478 39006 42530
rect 39006 42478 39058 42530
rect 39058 42478 39060 42530
rect 39004 42476 39060 42478
rect 39340 48412 39396 48468
rect 39340 47292 39396 47348
rect 39228 45948 39284 46004
rect 39340 45164 39396 45220
rect 39564 49922 39620 49924
rect 39564 49870 39566 49922
rect 39566 49870 39618 49922
rect 39618 49870 39620 49922
rect 39564 49868 39620 49870
rect 39676 49084 39732 49140
rect 39564 48972 39620 49028
rect 39564 48300 39620 48356
rect 40124 56140 40180 56196
rect 40012 54124 40068 54180
rect 41468 60732 41524 60788
rect 41692 62354 41748 62356
rect 41692 62302 41694 62354
rect 41694 62302 41746 62354
rect 41746 62302 41748 62354
rect 41692 62300 41748 62302
rect 42924 62354 42980 62356
rect 42924 62302 42926 62354
rect 42926 62302 42978 62354
rect 42978 62302 42980 62354
rect 42924 62300 42980 62302
rect 41916 61628 41972 61684
rect 41916 61010 41972 61012
rect 41916 60958 41918 61010
rect 41918 60958 41970 61010
rect 41970 60958 41972 61010
rect 41916 60956 41972 60958
rect 42476 61682 42532 61684
rect 42476 61630 42478 61682
rect 42478 61630 42530 61682
rect 42530 61630 42532 61682
rect 42476 61628 42532 61630
rect 40684 60284 40740 60340
rect 40460 60114 40516 60116
rect 40460 60062 40462 60114
rect 40462 60062 40514 60114
rect 40514 60062 40516 60114
rect 40460 60060 40516 60062
rect 41132 58268 41188 58324
rect 40572 58210 40628 58212
rect 40572 58158 40574 58210
rect 40574 58158 40626 58210
rect 40626 58158 40628 58210
rect 40572 58156 40628 58158
rect 40796 56866 40852 56868
rect 40796 56814 40798 56866
rect 40798 56814 40850 56866
rect 40850 56814 40852 56866
rect 40796 56812 40852 56814
rect 41020 56194 41076 56196
rect 41020 56142 41022 56194
rect 41022 56142 41074 56194
rect 41074 56142 41076 56194
rect 41020 56140 41076 56142
rect 40908 55916 40964 55972
rect 41580 55970 41636 55972
rect 41580 55918 41582 55970
rect 41582 55918 41634 55970
rect 41634 55918 41636 55970
rect 41580 55916 41636 55918
rect 40236 53058 40292 53060
rect 40236 53006 40238 53058
rect 40238 53006 40290 53058
rect 40290 53006 40292 53058
rect 40236 53004 40292 53006
rect 40012 51548 40068 51604
rect 40348 50764 40404 50820
rect 40684 55074 40740 55076
rect 40684 55022 40686 55074
rect 40686 55022 40738 55074
rect 40738 55022 40740 55074
rect 40684 55020 40740 55022
rect 40796 54348 40852 54404
rect 40684 53842 40740 53844
rect 40684 53790 40686 53842
rect 40686 53790 40738 53842
rect 40738 53790 40740 53842
rect 40684 53788 40740 53790
rect 42028 60508 42084 60564
rect 42140 61516 42196 61572
rect 43036 61628 43092 61684
rect 43148 61570 43204 61572
rect 43148 61518 43150 61570
rect 43150 61518 43202 61570
rect 43202 61518 43204 61570
rect 43148 61516 43204 61518
rect 41916 59388 41972 59444
rect 41916 57036 41972 57092
rect 43260 59276 43316 59332
rect 44044 62578 44100 62580
rect 44044 62526 44046 62578
rect 44046 62526 44098 62578
rect 44098 62526 44100 62578
rect 44044 62524 44100 62526
rect 44268 62860 44324 62916
rect 44044 62354 44100 62356
rect 44044 62302 44046 62354
rect 44046 62302 44098 62354
rect 44098 62302 44100 62354
rect 44044 62300 44100 62302
rect 43932 61404 43988 61460
rect 44604 67058 44660 67060
rect 44604 67006 44606 67058
rect 44606 67006 44658 67058
rect 44658 67006 44660 67058
rect 44604 67004 44660 67006
rect 45836 63810 45892 63812
rect 45836 63758 45838 63810
rect 45838 63758 45890 63810
rect 45890 63758 45892 63810
rect 45836 63756 45892 63758
rect 44940 63084 44996 63140
rect 45948 63196 46004 63252
rect 46060 63756 46116 63812
rect 45612 63138 45668 63140
rect 45612 63086 45614 63138
rect 45614 63086 45666 63138
rect 45666 63086 45668 63138
rect 45612 63084 45668 63086
rect 44604 62524 44660 62580
rect 46844 63250 46900 63252
rect 46844 63198 46846 63250
rect 46846 63198 46898 63250
rect 46898 63198 46900 63250
rect 46844 63196 46900 63198
rect 46620 63138 46676 63140
rect 46620 63086 46622 63138
rect 46622 63086 46674 63138
rect 46674 63086 46676 63138
rect 46620 63084 46676 63086
rect 44940 61458 44996 61460
rect 44940 61406 44942 61458
rect 44942 61406 44994 61458
rect 44994 61406 44996 61458
rect 44940 61404 44996 61406
rect 43372 58156 43428 58212
rect 43148 56812 43204 56868
rect 43036 56754 43092 56756
rect 43036 56702 43038 56754
rect 43038 56702 43090 56754
rect 43090 56702 43092 56754
rect 43036 56700 43092 56702
rect 42028 56194 42084 56196
rect 42028 56142 42030 56194
rect 42030 56142 42082 56194
rect 42082 56142 42084 56194
rect 42028 56140 42084 56142
rect 41692 54684 41748 54740
rect 42140 55468 42196 55524
rect 42028 54572 42084 54628
rect 41020 54348 41076 54404
rect 41692 54348 41748 54404
rect 41244 54124 41300 54180
rect 43148 55020 43204 55076
rect 43036 54572 43092 54628
rect 43708 56812 43764 56868
rect 44044 58210 44100 58212
rect 44044 58158 44046 58210
rect 44046 58158 44098 58210
rect 44098 58158 44100 58210
rect 44044 58156 44100 58158
rect 44492 57820 44548 57876
rect 45836 59330 45892 59332
rect 45836 59278 45838 59330
rect 45838 59278 45890 59330
rect 45890 59278 45892 59330
rect 45836 59276 45892 59278
rect 44604 57596 44660 57652
rect 44268 57538 44324 57540
rect 44268 57486 44270 57538
rect 44270 57486 44322 57538
rect 44322 57486 44324 57538
rect 44268 57484 44324 57486
rect 43596 56588 43652 56644
rect 43484 55132 43540 55188
rect 42140 54124 42196 54180
rect 41916 53788 41972 53844
rect 41132 53564 41188 53620
rect 41468 53564 41524 53620
rect 41132 53340 41188 53396
rect 40908 52892 40964 52948
rect 41020 53228 41076 53284
rect 41132 52332 41188 52388
rect 41244 53058 41300 53060
rect 41244 53006 41246 53058
rect 41246 53006 41298 53058
rect 41298 53006 41300 53058
rect 41244 53004 41300 53006
rect 41020 52220 41076 52276
rect 43148 54348 43204 54404
rect 42924 54012 42980 54068
rect 42140 53564 42196 53620
rect 41916 53340 41972 53396
rect 42364 53340 42420 53396
rect 42028 53228 42084 53284
rect 41804 52668 41860 52724
rect 41692 52386 41748 52388
rect 41692 52334 41694 52386
rect 41694 52334 41746 52386
rect 41746 52334 41748 52386
rect 41692 52332 41748 52334
rect 41244 52220 41300 52276
rect 41804 52108 41860 52164
rect 41916 52220 41972 52276
rect 41020 51884 41076 51940
rect 40012 49026 40068 49028
rect 40012 48974 40014 49026
rect 40014 48974 40066 49026
rect 40066 48974 40068 49026
rect 40012 48972 40068 48974
rect 40124 48914 40180 48916
rect 40124 48862 40126 48914
rect 40126 48862 40178 48914
rect 40178 48862 40180 48914
rect 40124 48860 40180 48862
rect 39900 47516 39956 47572
rect 40012 48748 40068 48804
rect 39788 47404 39844 47460
rect 40124 48130 40180 48132
rect 40124 48078 40126 48130
rect 40126 48078 40178 48130
rect 40178 48078 40180 48130
rect 40124 48076 40180 48078
rect 39676 47234 39732 47236
rect 39676 47182 39678 47234
rect 39678 47182 39730 47234
rect 39730 47182 39732 47234
rect 39676 47180 39732 47182
rect 39564 47068 39620 47124
rect 40236 47628 40292 47684
rect 40908 51100 40964 51156
rect 41132 51660 41188 51716
rect 40908 49980 40964 50036
rect 41020 49922 41076 49924
rect 41020 49870 41022 49922
rect 41022 49870 41074 49922
rect 41074 49870 41076 49922
rect 41020 49868 41076 49870
rect 41020 49586 41076 49588
rect 41020 49534 41022 49586
rect 41022 49534 41074 49586
rect 41074 49534 41076 49586
rect 41020 49532 41076 49534
rect 41132 48972 41188 49028
rect 40684 48748 40740 48804
rect 40460 48300 40516 48356
rect 41356 48300 41412 48356
rect 40460 47346 40516 47348
rect 40460 47294 40462 47346
rect 40462 47294 40514 47346
rect 40514 47294 40516 47346
rect 40460 47292 40516 47294
rect 40236 47180 40292 47236
rect 39900 46002 39956 46004
rect 39900 45950 39902 46002
rect 39902 45950 39954 46002
rect 39954 45950 39956 46002
rect 39900 45948 39956 45950
rect 39676 44940 39732 44996
rect 38892 41132 38948 41188
rect 38556 40236 38612 40292
rect 38892 40402 38948 40404
rect 38892 40350 38894 40402
rect 38894 40350 38946 40402
rect 38946 40350 38948 40402
rect 38892 40348 38948 40350
rect 38668 38780 38724 38836
rect 37884 36652 37940 36708
rect 37772 35532 37828 35588
rect 37772 34914 37828 34916
rect 37772 34862 37774 34914
rect 37774 34862 37826 34914
rect 37826 34862 37828 34914
rect 37772 34860 37828 34862
rect 37884 36316 37940 36372
rect 39116 40962 39172 40964
rect 39116 40910 39118 40962
rect 39118 40910 39170 40962
rect 39170 40910 39172 40962
rect 39116 40908 39172 40910
rect 39116 40626 39172 40628
rect 39116 40574 39118 40626
rect 39118 40574 39170 40626
rect 39170 40574 39172 40626
rect 39116 40572 39172 40574
rect 39900 45218 39956 45220
rect 39900 45166 39902 45218
rect 39902 45166 39954 45218
rect 39954 45166 39956 45218
rect 39900 45164 39956 45166
rect 40572 47234 40628 47236
rect 40572 47182 40574 47234
rect 40574 47182 40626 47234
rect 40626 47182 40628 47234
rect 40572 47180 40628 47182
rect 40572 45948 40628 46004
rect 40460 45500 40516 45556
rect 40348 45276 40404 45332
rect 40124 45164 40180 45220
rect 40012 45052 40068 45108
rect 40908 47292 40964 47348
rect 41020 48076 41076 48132
rect 40796 47234 40852 47236
rect 40796 47182 40798 47234
rect 40798 47182 40850 47234
rect 40850 47182 40852 47234
rect 40796 47180 40852 47182
rect 41020 47068 41076 47124
rect 41020 45948 41076 46004
rect 40796 45890 40852 45892
rect 40796 45838 40798 45890
rect 40798 45838 40850 45890
rect 40850 45838 40852 45890
rect 40796 45836 40852 45838
rect 41244 45500 41300 45556
rect 41580 50034 41636 50036
rect 41580 49982 41582 50034
rect 41582 49982 41634 50034
rect 41634 49982 41636 50034
rect 41580 49980 41636 49982
rect 41580 48914 41636 48916
rect 41580 48862 41582 48914
rect 41582 48862 41634 48914
rect 41634 48862 41636 48914
rect 41580 48860 41636 48862
rect 39900 43932 39956 43988
rect 40348 43708 40404 43764
rect 39900 43372 39956 43428
rect 39340 42140 39396 42196
rect 39340 40572 39396 40628
rect 39452 41916 39508 41972
rect 39676 42476 39732 42532
rect 40012 41244 40068 41300
rect 39788 41186 39844 41188
rect 39788 41134 39790 41186
rect 39790 41134 39842 41186
rect 39842 41134 39844 41186
rect 39788 41132 39844 41134
rect 40684 44716 40740 44772
rect 40684 44210 40740 44212
rect 40684 44158 40686 44210
rect 40686 44158 40738 44210
rect 40738 44158 40740 44210
rect 40684 44156 40740 44158
rect 41020 44210 41076 44212
rect 41020 44158 41022 44210
rect 41022 44158 41074 44210
rect 41074 44158 41076 44210
rect 41020 44156 41076 44158
rect 40796 43932 40852 43988
rect 40684 43820 40740 43876
rect 41020 43762 41076 43764
rect 41020 43710 41022 43762
rect 41022 43710 41074 43762
rect 41074 43710 41076 43762
rect 41020 43708 41076 43710
rect 41580 48524 41636 48580
rect 41356 45106 41412 45108
rect 41356 45054 41358 45106
rect 41358 45054 41410 45106
rect 41410 45054 41412 45106
rect 41356 45052 41412 45054
rect 41468 44492 41524 44548
rect 42028 51324 42084 51380
rect 42028 50988 42084 51044
rect 44604 57372 44660 57428
rect 44604 56924 44660 56980
rect 45612 57874 45668 57876
rect 45612 57822 45614 57874
rect 45614 57822 45666 57874
rect 45666 57822 45668 57874
rect 45612 57820 45668 57822
rect 45500 57484 45556 57540
rect 45164 57148 45220 57204
rect 44604 55916 44660 55972
rect 43932 55186 43988 55188
rect 43932 55134 43934 55186
rect 43934 55134 43986 55186
rect 43986 55134 43988 55186
rect 43932 55132 43988 55134
rect 44044 55074 44100 55076
rect 44044 55022 44046 55074
rect 44046 55022 44098 55074
rect 44098 55022 44100 55074
rect 44044 55020 44100 55022
rect 43596 54626 43652 54628
rect 43596 54574 43598 54626
rect 43598 54574 43650 54626
rect 43650 54574 43652 54626
rect 43596 54572 43652 54574
rect 43484 54012 43540 54068
rect 43820 54402 43876 54404
rect 43820 54350 43822 54402
rect 43822 54350 43874 54402
rect 43874 54350 43876 54402
rect 43820 54348 43876 54350
rect 42700 51436 42756 51492
rect 42588 51378 42644 51380
rect 42588 51326 42590 51378
rect 42590 51326 42642 51378
rect 42642 51326 42644 51378
rect 42588 51324 42644 51326
rect 41804 47628 41860 47684
rect 41804 47068 41860 47124
rect 42252 47180 42308 47236
rect 43036 50706 43092 50708
rect 43036 50654 43038 50706
rect 43038 50654 43090 50706
rect 43090 50654 43092 50706
rect 43036 50652 43092 50654
rect 42812 49532 42868 49588
rect 43260 49196 43316 49252
rect 43260 48412 43316 48468
rect 42812 47628 42868 47684
rect 42812 47180 42868 47236
rect 42252 45890 42308 45892
rect 42252 45838 42254 45890
rect 42254 45838 42306 45890
rect 42306 45838 42308 45890
rect 42252 45836 42308 45838
rect 41580 44380 41636 44436
rect 41692 45164 41748 45220
rect 41356 44268 41412 44324
rect 41692 43932 41748 43988
rect 41580 43538 41636 43540
rect 41580 43486 41582 43538
rect 41582 43486 41634 43538
rect 41634 43486 41636 43538
rect 41580 43484 41636 43486
rect 41244 42866 41300 42868
rect 41244 42814 41246 42866
rect 41246 42814 41298 42866
rect 41298 42814 41300 42866
rect 41244 42812 41300 42814
rect 40684 42028 40740 42084
rect 40572 41244 40628 41300
rect 39788 40572 39844 40628
rect 39564 39564 39620 39620
rect 39340 39506 39396 39508
rect 39340 39454 39342 39506
rect 39342 39454 39394 39506
rect 39394 39454 39396 39506
rect 39340 39452 39396 39454
rect 39676 39506 39732 39508
rect 39676 39454 39678 39506
rect 39678 39454 39730 39506
rect 39730 39454 39732 39506
rect 39676 39452 39732 39454
rect 39340 38892 39396 38948
rect 38108 37378 38164 37380
rect 38108 37326 38110 37378
rect 38110 37326 38162 37378
rect 38162 37326 38164 37378
rect 38108 37324 38164 37326
rect 38780 38050 38836 38052
rect 38780 37998 38782 38050
rect 38782 37998 38834 38050
rect 38834 37998 38836 38050
rect 38780 37996 38836 37998
rect 38332 36428 38388 36484
rect 39116 36370 39172 36372
rect 39116 36318 39118 36370
rect 39118 36318 39170 36370
rect 39170 36318 39172 36370
rect 39116 36316 39172 36318
rect 37548 33628 37604 33684
rect 37212 33068 37268 33124
rect 37212 32674 37268 32676
rect 37212 32622 37214 32674
rect 37214 32622 37266 32674
rect 37266 32622 37268 32674
rect 37212 32620 37268 32622
rect 37436 32562 37492 32564
rect 37436 32510 37438 32562
rect 37438 32510 37490 32562
rect 37490 32510 37492 32562
rect 37436 32508 37492 32510
rect 36876 32284 36932 32340
rect 37436 31612 37492 31668
rect 36988 30210 37044 30212
rect 36988 30158 36990 30210
rect 36990 30158 37042 30210
rect 37042 30158 37044 30210
rect 36988 30156 37044 30158
rect 37884 33404 37940 33460
rect 38108 35420 38164 35476
rect 38444 35644 38500 35700
rect 39228 36204 39284 36260
rect 39564 37996 39620 38052
rect 39900 38050 39956 38052
rect 39900 37998 39902 38050
rect 39902 37998 39954 38050
rect 39954 37998 39956 38050
rect 39900 37996 39956 37998
rect 39788 37324 39844 37380
rect 39452 36482 39508 36484
rect 39452 36430 39454 36482
rect 39454 36430 39506 36482
rect 39506 36430 39508 36482
rect 39452 36428 39508 36430
rect 39004 35698 39060 35700
rect 39004 35646 39006 35698
rect 39006 35646 39058 35698
rect 39058 35646 39060 35698
rect 39004 35644 39060 35646
rect 40684 40572 40740 40628
rect 40236 40514 40292 40516
rect 40236 40462 40238 40514
rect 40238 40462 40290 40514
rect 40290 40462 40292 40514
rect 40236 40460 40292 40462
rect 40796 40460 40852 40516
rect 40236 39618 40292 39620
rect 40236 39566 40238 39618
rect 40238 39566 40290 39618
rect 40290 39566 40292 39618
rect 40236 39564 40292 39566
rect 40460 38780 40516 38836
rect 40124 36764 40180 36820
rect 40236 36876 40292 36932
rect 39900 36370 39956 36372
rect 39900 36318 39902 36370
rect 39902 36318 39954 36370
rect 39954 36318 39956 36370
rect 39900 36316 39956 36318
rect 39004 35474 39060 35476
rect 39004 35422 39006 35474
rect 39006 35422 39058 35474
rect 39058 35422 39060 35474
rect 39004 35420 39060 35422
rect 38556 35196 38612 35252
rect 38332 34860 38388 34916
rect 39340 35196 39396 35252
rect 39788 36204 39844 36260
rect 39788 35644 39844 35700
rect 39900 36092 39956 36148
rect 38332 33628 38388 33684
rect 38556 32508 38612 32564
rect 39676 34748 39732 34804
rect 39004 33964 39060 34020
rect 39676 34018 39732 34020
rect 39676 33966 39678 34018
rect 39678 33966 39730 34018
rect 39730 33966 39732 34018
rect 39676 33964 39732 33966
rect 40348 36092 40404 36148
rect 40236 35644 40292 35700
rect 40348 34188 40404 34244
rect 40572 35644 40628 35700
rect 41244 41132 41300 41188
rect 41244 40684 41300 40740
rect 41132 39564 41188 39620
rect 40796 39004 40852 39060
rect 41020 38892 41076 38948
rect 41244 39506 41300 39508
rect 41244 39454 41246 39506
rect 41246 39454 41298 39506
rect 41298 39454 41300 39506
rect 41244 39452 41300 39454
rect 41132 37266 41188 37268
rect 41132 37214 41134 37266
rect 41134 37214 41186 37266
rect 41186 37214 41188 37266
rect 41132 37212 41188 37214
rect 41132 36764 41188 36820
rect 41244 36482 41300 36484
rect 41244 36430 41246 36482
rect 41246 36430 41298 36482
rect 41298 36430 41300 36482
rect 41244 36428 41300 36430
rect 41132 35810 41188 35812
rect 41132 35758 41134 35810
rect 41134 35758 41186 35810
rect 41186 35758 41188 35810
rect 41132 35756 41188 35758
rect 41580 41298 41636 41300
rect 41580 41246 41582 41298
rect 41582 41246 41634 41298
rect 41634 41246 41636 41298
rect 41580 41244 41636 41246
rect 41580 41020 41636 41076
rect 41692 40626 41748 40628
rect 41692 40574 41694 40626
rect 41694 40574 41746 40626
rect 41746 40574 41748 40626
rect 41692 40572 41748 40574
rect 42028 45218 42084 45220
rect 42028 45166 42030 45218
rect 42030 45166 42082 45218
rect 42082 45166 42084 45218
rect 42028 45164 42084 45166
rect 42028 43708 42084 43764
rect 41916 42866 41972 42868
rect 41916 42814 41918 42866
rect 41918 42814 41970 42866
rect 41970 42814 41972 42866
rect 41916 42812 41972 42814
rect 41916 42476 41972 42532
rect 42028 41020 42084 41076
rect 41916 40684 41972 40740
rect 41580 40124 41636 40180
rect 41580 39618 41636 39620
rect 41580 39566 41582 39618
rect 41582 39566 41634 39618
rect 41634 39566 41636 39618
rect 41580 39564 41636 39566
rect 42252 40626 42308 40628
rect 42252 40574 42254 40626
rect 42254 40574 42306 40626
rect 42306 40574 42308 40626
rect 42252 40572 42308 40574
rect 41916 39618 41972 39620
rect 41916 39566 41918 39618
rect 41918 39566 41970 39618
rect 41970 39566 41972 39618
rect 41916 39564 41972 39566
rect 41804 39058 41860 39060
rect 41804 39006 41806 39058
rect 41806 39006 41858 39058
rect 41858 39006 41860 39058
rect 41804 39004 41860 39006
rect 42252 39452 42308 39508
rect 41692 38892 41748 38948
rect 41804 37266 41860 37268
rect 41804 37214 41806 37266
rect 41806 37214 41858 37266
rect 41858 37214 41860 37266
rect 41804 37212 41860 37214
rect 42140 37266 42196 37268
rect 42140 37214 42142 37266
rect 42142 37214 42194 37266
rect 42194 37214 42196 37266
rect 42140 37212 42196 37214
rect 41692 36482 41748 36484
rect 41692 36430 41694 36482
rect 41694 36430 41746 36482
rect 41746 36430 41748 36482
rect 41692 36428 41748 36430
rect 40460 33852 40516 33908
rect 40908 34802 40964 34804
rect 40908 34750 40910 34802
rect 40910 34750 40962 34802
rect 40962 34750 40964 34802
rect 40908 34748 40964 34750
rect 41244 34914 41300 34916
rect 41244 34862 41246 34914
rect 41246 34862 41298 34914
rect 41298 34862 41300 34914
rect 41244 34860 41300 34862
rect 41692 35474 41748 35476
rect 41692 35422 41694 35474
rect 41694 35422 41746 35474
rect 41746 35422 41748 35474
rect 41692 35420 41748 35422
rect 41692 35084 41748 35140
rect 40908 33852 40964 33908
rect 39788 33234 39844 33236
rect 39788 33182 39790 33234
rect 39790 33182 39842 33234
rect 39842 33182 39844 33234
rect 39788 33180 39844 33182
rect 39564 33068 39620 33124
rect 39788 32844 39844 32900
rect 38780 31612 38836 31668
rect 38556 31500 38612 31556
rect 37100 29932 37156 29988
rect 38444 29820 38500 29876
rect 38108 28700 38164 28756
rect 37660 28530 37716 28532
rect 37660 28478 37662 28530
rect 37662 28478 37714 28530
rect 37714 28478 37716 28530
rect 37660 28476 37716 28478
rect 37548 28028 37604 28084
rect 36988 27132 37044 27188
rect 37212 24892 37268 24948
rect 37436 23436 37492 23492
rect 37660 27298 37716 27300
rect 37660 27246 37662 27298
rect 37662 27246 37714 27298
rect 37714 27246 37716 27298
rect 37660 27244 37716 27246
rect 37996 27298 38052 27300
rect 37996 27246 37998 27298
rect 37998 27246 38050 27298
rect 38050 27246 38052 27298
rect 37996 27244 38052 27246
rect 37996 25004 38052 25060
rect 37884 24946 37940 24948
rect 37884 24894 37886 24946
rect 37886 24894 37938 24946
rect 37938 24894 37940 24946
rect 37884 24892 37940 24894
rect 37660 24556 37716 24612
rect 37660 23714 37716 23716
rect 37660 23662 37662 23714
rect 37662 23662 37714 23714
rect 37714 23662 37716 23714
rect 37660 23660 37716 23662
rect 37436 22204 37492 22260
rect 37436 21868 37492 21924
rect 37324 20076 37380 20132
rect 37100 19740 37156 19796
rect 36876 19516 36932 19572
rect 37212 19346 37268 19348
rect 37212 19294 37214 19346
rect 37214 19294 37266 19346
rect 37266 19294 37268 19346
rect 37212 19292 37268 19294
rect 36988 19234 37044 19236
rect 36988 19182 36990 19234
rect 36990 19182 37042 19234
rect 37042 19182 37044 19234
rect 36988 19180 37044 19182
rect 37100 18508 37156 18564
rect 37212 18172 37268 18228
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34188 11452 34244 11508
rect 33740 11394 33796 11396
rect 33740 11342 33742 11394
rect 33742 11342 33794 11394
rect 33794 11342 33796 11394
rect 33740 11340 33796 11342
rect 35420 14364 35476 14420
rect 35532 14252 35588 14308
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35868 15260 35924 15316
rect 36092 15314 36148 15316
rect 36092 15262 36094 15314
rect 36094 15262 36146 15314
rect 36146 15262 36148 15314
rect 36092 15260 36148 15262
rect 36764 15260 36820 15316
rect 35868 14642 35924 14644
rect 35868 14590 35870 14642
rect 35870 14590 35922 14642
rect 35922 14590 35924 14642
rect 35868 14588 35924 14590
rect 38668 28476 38724 28532
rect 38556 27858 38612 27860
rect 38556 27806 38558 27858
rect 38558 27806 38610 27858
rect 38610 27806 38612 27858
rect 38556 27804 38612 27806
rect 38332 27356 38388 27412
rect 38668 27020 38724 27076
rect 38780 28364 38836 28420
rect 38780 27244 38836 27300
rect 38444 25004 38500 25060
rect 38332 23212 38388 23268
rect 38780 25116 38836 25172
rect 39788 31666 39844 31668
rect 39788 31614 39790 31666
rect 39790 31614 39842 31666
rect 39842 31614 39844 31666
rect 39788 31612 39844 31614
rect 39116 29820 39172 29876
rect 39564 29820 39620 29876
rect 39564 29260 39620 29316
rect 39004 29202 39060 29204
rect 39004 29150 39006 29202
rect 39006 29150 39058 29202
rect 39058 29150 39060 29202
rect 39004 29148 39060 29150
rect 39452 28866 39508 28868
rect 39452 28814 39454 28866
rect 39454 28814 39506 28866
rect 39506 28814 39508 28866
rect 39452 28812 39508 28814
rect 39116 28588 39172 28644
rect 39004 28530 39060 28532
rect 39004 28478 39006 28530
rect 39006 28478 39058 28530
rect 39058 28478 39060 28530
rect 39004 28476 39060 28478
rect 39004 28028 39060 28084
rect 39004 26460 39060 26516
rect 39340 28530 39396 28532
rect 39340 28478 39342 28530
rect 39342 28478 39394 28530
rect 39394 28478 39396 28530
rect 39340 28476 39396 28478
rect 39452 28418 39508 28420
rect 39452 28366 39454 28418
rect 39454 28366 39506 28418
rect 39506 28366 39508 28418
rect 39452 28364 39508 28366
rect 39340 28028 39396 28084
rect 39564 27916 39620 27972
rect 40124 33122 40180 33124
rect 40124 33070 40126 33122
rect 40126 33070 40178 33122
rect 40178 33070 40180 33122
rect 40124 33068 40180 33070
rect 40012 32844 40068 32900
rect 40012 29708 40068 29764
rect 39900 29260 39956 29316
rect 40460 32732 40516 32788
rect 40348 32674 40404 32676
rect 40348 32622 40350 32674
rect 40350 32622 40402 32674
rect 40402 32622 40404 32674
rect 40348 32620 40404 32622
rect 40348 30044 40404 30100
rect 40348 29650 40404 29652
rect 40348 29598 40350 29650
rect 40350 29598 40402 29650
rect 40402 29598 40404 29650
rect 40348 29596 40404 29598
rect 41244 33628 41300 33684
rect 41132 33180 41188 33236
rect 40908 32732 40964 32788
rect 41356 33068 41412 33124
rect 41692 32956 41748 33012
rect 41244 32674 41300 32676
rect 41244 32622 41246 32674
rect 41246 32622 41298 32674
rect 41298 32622 41300 32674
rect 41244 32620 41300 32622
rect 40684 31554 40740 31556
rect 40684 31502 40686 31554
rect 40686 31502 40738 31554
rect 40738 31502 40740 31554
rect 40684 31500 40740 31502
rect 40572 29708 40628 29764
rect 40460 29260 40516 29316
rect 40460 28924 40516 28980
rect 40236 28082 40292 28084
rect 40236 28030 40238 28082
rect 40238 28030 40290 28082
rect 40290 28030 40292 28082
rect 40236 28028 40292 28030
rect 40124 27916 40180 27972
rect 40348 27858 40404 27860
rect 40348 27806 40350 27858
rect 40350 27806 40402 27858
rect 40402 27806 40404 27858
rect 40348 27804 40404 27806
rect 40236 27634 40292 27636
rect 40236 27582 40238 27634
rect 40238 27582 40290 27634
rect 40290 27582 40292 27634
rect 40236 27580 40292 27582
rect 39564 25116 39620 25172
rect 39788 27356 39844 27412
rect 39452 25004 39508 25060
rect 39900 27074 39956 27076
rect 39900 27022 39902 27074
rect 39902 27022 39954 27074
rect 39954 27022 39956 27074
rect 39900 27020 39956 27022
rect 38668 22764 38724 22820
rect 37884 22316 37940 22372
rect 38556 22316 38612 22372
rect 38332 22258 38388 22260
rect 38332 22206 38334 22258
rect 38334 22206 38386 22258
rect 38386 22206 38388 22258
rect 38332 22204 38388 22206
rect 37548 19906 37604 19908
rect 37548 19854 37550 19906
rect 37550 19854 37602 19906
rect 37602 19854 37604 19906
rect 37548 19852 37604 19854
rect 37884 19964 37940 20020
rect 37548 19516 37604 19572
rect 37436 18620 37492 18676
rect 37548 18732 37604 18788
rect 37660 18620 37716 18676
rect 38108 20130 38164 20132
rect 38108 20078 38110 20130
rect 38110 20078 38162 20130
rect 38162 20078 38164 20130
rect 38108 20076 38164 20078
rect 38220 20018 38276 20020
rect 38220 19966 38222 20018
rect 38222 19966 38274 20018
rect 38274 19966 38276 20018
rect 38220 19964 38276 19966
rect 37996 19740 38052 19796
rect 38332 19234 38388 19236
rect 38332 19182 38334 19234
rect 38334 19182 38386 19234
rect 38386 19182 38388 19234
rect 38332 19180 38388 19182
rect 37884 18620 37940 18676
rect 38220 19010 38276 19012
rect 38220 18958 38222 19010
rect 38222 18958 38274 19010
rect 38274 18958 38276 19010
rect 38220 18956 38276 18958
rect 38220 18732 38276 18788
rect 38332 18620 38388 18676
rect 39340 23154 39396 23156
rect 39340 23102 39342 23154
rect 39342 23102 39394 23154
rect 39394 23102 39396 23154
rect 39340 23100 39396 23102
rect 39900 25004 39956 25060
rect 39788 24722 39844 24724
rect 39788 24670 39790 24722
rect 39790 24670 39842 24722
rect 39842 24670 39844 24722
rect 39788 24668 39844 24670
rect 39788 23436 39844 23492
rect 39452 22540 39508 22596
rect 39340 21868 39396 21924
rect 39116 20914 39172 20916
rect 39116 20862 39118 20914
rect 39118 20862 39170 20914
rect 39170 20862 39172 20914
rect 39116 20860 39172 20862
rect 38556 19964 38612 20020
rect 38780 20018 38836 20020
rect 38780 19966 38782 20018
rect 38782 19966 38834 20018
rect 38834 19966 38836 20018
rect 38780 19964 38836 19966
rect 39788 20860 39844 20916
rect 39788 20300 39844 20356
rect 40012 24834 40068 24836
rect 40012 24782 40014 24834
rect 40014 24782 40066 24834
rect 40066 24782 40068 24834
rect 40012 24780 40068 24782
rect 40012 22482 40068 22484
rect 40012 22430 40014 22482
rect 40014 22430 40066 22482
rect 40066 22430 40068 22482
rect 40012 22428 40068 22430
rect 39900 20076 39956 20132
rect 39564 19292 39620 19348
rect 38668 18620 38724 18676
rect 39228 18620 39284 18676
rect 38108 18396 38164 18452
rect 39004 18450 39060 18452
rect 39004 18398 39006 18450
rect 39006 18398 39058 18450
rect 39058 18398 39060 18450
rect 39004 18396 39060 18398
rect 38668 18172 38724 18228
rect 38780 18284 38836 18340
rect 37884 17554 37940 17556
rect 37884 17502 37886 17554
rect 37886 17502 37938 17554
rect 37938 17502 37940 17554
rect 37884 17500 37940 17502
rect 38556 17948 38612 18004
rect 38332 17442 38388 17444
rect 38332 17390 38334 17442
rect 38334 17390 38386 17442
rect 38386 17390 38388 17442
rect 38332 17388 38388 17390
rect 38556 17388 38612 17444
rect 37548 15538 37604 15540
rect 37548 15486 37550 15538
rect 37550 15486 37602 15538
rect 37602 15486 37604 15538
rect 37548 15484 37604 15486
rect 37436 15314 37492 15316
rect 37436 15262 37438 15314
rect 37438 15262 37490 15314
rect 37490 15262 37492 15314
rect 37436 15260 37492 15262
rect 36876 14476 36932 14532
rect 36988 15148 37044 15204
rect 36876 14306 36932 14308
rect 36876 14254 36878 14306
rect 36878 14254 36930 14306
rect 36930 14254 36932 14306
rect 36876 14252 36932 14254
rect 36092 14140 36148 14196
rect 37996 15484 38052 15540
rect 37772 15314 37828 15316
rect 37772 15262 37774 15314
rect 37774 15262 37826 15314
rect 37826 15262 37828 15314
rect 37772 15260 37828 15262
rect 37100 14140 37156 14196
rect 37212 14530 37268 14532
rect 37212 14478 37214 14530
rect 37214 14478 37266 14530
rect 37266 14478 37268 14530
rect 37212 14476 37268 14478
rect 36204 13356 36260 13412
rect 35532 12236 35588 12292
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34972 10668 35028 10724
rect 33628 9884 33684 9940
rect 34188 10444 34244 10500
rect 33516 8988 33572 9044
rect 33180 6524 33236 6580
rect 33404 7980 33460 8036
rect 34972 10444 35028 10500
rect 34524 8428 34580 8484
rect 34412 8204 34468 8260
rect 34636 8034 34692 8036
rect 34636 7982 34638 8034
rect 34638 7982 34690 8034
rect 34690 7982 34692 8034
rect 34636 7980 34692 7982
rect 35644 10722 35700 10724
rect 35644 10670 35646 10722
rect 35646 10670 35698 10722
rect 35698 10670 35700 10722
rect 35644 10668 35700 10670
rect 35532 10556 35588 10612
rect 35420 10444 35476 10500
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35084 8482 35140 8484
rect 35084 8430 35086 8482
rect 35086 8430 35138 8482
rect 35138 8430 35140 8482
rect 35084 8428 35140 8430
rect 37548 13858 37604 13860
rect 37548 13806 37550 13858
rect 37550 13806 37602 13858
rect 37602 13806 37604 13858
rect 37548 13804 37604 13806
rect 36652 13356 36708 13412
rect 36204 11282 36260 11284
rect 36204 11230 36206 11282
rect 36206 11230 36258 11282
rect 36258 11230 36260 11282
rect 36204 11228 36260 11230
rect 36316 11340 36372 11396
rect 36764 10498 36820 10500
rect 36764 10446 36766 10498
rect 36766 10446 36818 10498
rect 36818 10446 36820 10498
rect 36764 10444 36820 10446
rect 36540 8988 36596 9044
rect 37100 13356 37156 13412
rect 37324 11394 37380 11396
rect 37324 11342 37326 11394
rect 37326 11342 37378 11394
rect 37378 11342 37380 11394
rect 37324 11340 37380 11342
rect 37548 10610 37604 10612
rect 37548 10558 37550 10610
rect 37550 10558 37602 10610
rect 37602 10558 37604 10610
rect 37548 10556 37604 10558
rect 37436 9714 37492 9716
rect 37436 9662 37438 9714
rect 37438 9662 37490 9714
rect 37490 9662 37492 9714
rect 37436 9660 37492 9662
rect 38556 15372 38612 15428
rect 38332 14642 38388 14644
rect 38332 14590 38334 14642
rect 38334 14590 38386 14642
rect 38386 14590 38388 14642
rect 38332 14588 38388 14590
rect 38220 14364 38276 14420
rect 38220 13970 38276 13972
rect 38220 13918 38222 13970
rect 38222 13918 38274 13970
rect 38274 13918 38276 13970
rect 38220 13916 38276 13918
rect 38108 13858 38164 13860
rect 38108 13806 38110 13858
rect 38110 13806 38162 13858
rect 38162 13806 38164 13858
rect 38108 13804 38164 13806
rect 38444 13580 38500 13636
rect 38220 11340 38276 11396
rect 37996 9826 38052 9828
rect 37996 9774 37998 9826
rect 37998 9774 38050 9826
rect 38050 9774 38052 9826
rect 37996 9772 38052 9774
rect 38892 17836 38948 17892
rect 38780 17612 38836 17668
rect 38780 17106 38836 17108
rect 38780 17054 38782 17106
rect 38782 17054 38834 17106
rect 38834 17054 38836 17106
rect 38780 17052 38836 17054
rect 38780 15260 38836 15316
rect 38780 13746 38836 13748
rect 38780 13694 38782 13746
rect 38782 13694 38834 13746
rect 38834 13694 38836 13746
rect 38780 13692 38836 13694
rect 38668 13356 38724 13412
rect 38780 11900 38836 11956
rect 39452 18450 39508 18452
rect 39452 18398 39454 18450
rect 39454 18398 39506 18450
rect 39506 18398 39508 18450
rect 39452 18396 39508 18398
rect 39676 19234 39732 19236
rect 39676 19182 39678 19234
rect 39678 19182 39730 19234
rect 39730 19182 39732 19234
rect 39676 19180 39732 19182
rect 39900 19180 39956 19236
rect 39228 17724 39284 17780
rect 39004 17666 39060 17668
rect 39004 17614 39006 17666
rect 39006 17614 39058 17666
rect 39058 17614 39060 17666
rect 39004 17612 39060 17614
rect 39676 17778 39732 17780
rect 39676 17726 39678 17778
rect 39678 17726 39730 17778
rect 39730 17726 39732 17778
rect 39676 17724 39732 17726
rect 40684 29372 40740 29428
rect 40908 29708 40964 29764
rect 41356 31890 41412 31892
rect 41356 31838 41358 31890
rect 41358 31838 41410 31890
rect 41410 31838 41412 31890
rect 41356 31836 41412 31838
rect 41244 30716 41300 30772
rect 41132 30210 41188 30212
rect 41132 30158 41134 30210
rect 41134 30158 41186 30210
rect 41186 30158 41188 30210
rect 41132 30156 41188 30158
rect 41356 30044 41412 30100
rect 41692 32786 41748 32788
rect 41692 32734 41694 32786
rect 41694 32734 41746 32786
rect 41746 32734 41748 32786
rect 41692 32732 41748 32734
rect 42700 46620 42756 46676
rect 42588 44716 42644 44772
rect 43260 45836 43316 45892
rect 42588 44492 42644 44548
rect 43484 50652 43540 50708
rect 43820 51490 43876 51492
rect 43820 51438 43822 51490
rect 43822 51438 43874 51490
rect 43874 51438 43876 51490
rect 43820 51436 43876 51438
rect 44044 51324 44100 51380
rect 43820 51212 43876 51268
rect 43708 49532 43764 49588
rect 43820 48300 43876 48356
rect 43820 46674 43876 46676
rect 43820 46622 43822 46674
rect 43822 46622 43874 46674
rect 43874 46622 43876 46674
rect 43820 46620 43876 46622
rect 43708 46002 43764 46004
rect 43708 45950 43710 46002
rect 43710 45950 43762 46002
rect 43762 45950 43764 46002
rect 43708 45948 43764 45950
rect 42812 43708 42868 43764
rect 43036 43538 43092 43540
rect 43036 43486 43038 43538
rect 43038 43486 43090 43538
rect 43090 43486 43092 43538
rect 43036 43484 43092 43486
rect 42476 42530 42532 42532
rect 42476 42478 42478 42530
rect 42478 42478 42530 42530
rect 42530 42478 42532 42530
rect 42476 42476 42532 42478
rect 42700 41020 42756 41076
rect 42476 39564 42532 39620
rect 43036 39564 43092 39620
rect 44268 53842 44324 53844
rect 44268 53790 44270 53842
rect 44270 53790 44322 53842
rect 44322 53790 44324 53842
rect 44268 53788 44324 53790
rect 44268 50482 44324 50484
rect 44268 50430 44270 50482
rect 44270 50430 44322 50482
rect 44322 50430 44324 50482
rect 44268 50428 44324 50430
rect 44492 48354 44548 48356
rect 44492 48302 44494 48354
rect 44494 48302 44546 48354
rect 44546 48302 44548 48354
rect 44492 48300 44548 48302
rect 44156 46620 44212 46676
rect 44044 45890 44100 45892
rect 44044 45838 44046 45890
rect 44046 45838 44098 45890
rect 44098 45838 44100 45890
rect 44044 45836 44100 45838
rect 44940 53788 44996 53844
rect 45052 56924 45108 56980
rect 46060 57148 46116 57204
rect 45500 57036 45556 57092
rect 45276 55020 45332 55076
rect 45164 53900 45220 53956
rect 43596 40796 43652 40852
rect 43708 40402 43764 40404
rect 43708 40350 43710 40402
rect 43710 40350 43762 40402
rect 43762 40350 43764 40402
rect 43708 40348 43764 40350
rect 43596 39900 43652 39956
rect 43932 40348 43988 40404
rect 44156 39900 44212 39956
rect 44156 39564 44212 39620
rect 43708 38946 43764 38948
rect 43708 38894 43710 38946
rect 43710 38894 43762 38946
rect 43762 38894 43764 38946
rect 43708 38892 43764 38894
rect 42364 38556 42420 38612
rect 42364 35810 42420 35812
rect 42364 35758 42366 35810
rect 42366 35758 42418 35810
rect 42418 35758 42420 35810
rect 42364 35756 42420 35758
rect 42028 33628 42084 33684
rect 41916 31836 41972 31892
rect 42476 34914 42532 34916
rect 42476 34862 42478 34914
rect 42478 34862 42530 34914
rect 42530 34862 42532 34914
rect 42476 34860 42532 34862
rect 43036 37212 43092 37268
rect 43484 37212 43540 37268
rect 43596 36540 43652 36596
rect 43148 35420 43204 35476
rect 42924 33628 42980 33684
rect 44044 38892 44100 38948
rect 42700 33346 42756 33348
rect 42700 33294 42702 33346
rect 42702 33294 42754 33346
rect 42754 33294 42756 33346
rect 42700 33292 42756 33294
rect 42476 33122 42532 33124
rect 42476 33070 42478 33122
rect 42478 33070 42530 33122
rect 42530 33070 42532 33122
rect 42476 33068 42532 33070
rect 42028 31388 42084 31444
rect 41468 29426 41524 29428
rect 41468 29374 41470 29426
rect 41470 29374 41522 29426
rect 41522 29374 41524 29426
rect 41468 29372 41524 29374
rect 41244 28924 41300 28980
rect 41020 27356 41076 27412
rect 41244 27298 41300 27300
rect 41244 27246 41246 27298
rect 41246 27246 41298 27298
rect 41298 27246 41300 27298
rect 41244 27244 41300 27246
rect 40348 24722 40404 24724
rect 40348 24670 40350 24722
rect 40350 24670 40402 24722
rect 40402 24670 40404 24722
rect 40348 24668 40404 24670
rect 40236 23436 40292 23492
rect 40572 22482 40628 22484
rect 40572 22430 40574 22482
rect 40574 22430 40626 22482
rect 40626 22430 40628 22482
rect 40572 22428 40628 22430
rect 40236 20018 40292 20020
rect 40236 19966 40238 20018
rect 40238 19966 40290 20018
rect 40290 19966 40292 20018
rect 40236 19964 40292 19966
rect 40236 19292 40292 19348
rect 40348 18562 40404 18564
rect 40348 18510 40350 18562
rect 40350 18510 40402 18562
rect 40402 18510 40404 18562
rect 40348 18508 40404 18510
rect 40124 18284 40180 18340
rect 40348 18284 40404 18340
rect 40124 17778 40180 17780
rect 40124 17726 40126 17778
rect 40126 17726 40178 17778
rect 40178 17726 40180 17778
rect 40124 17724 40180 17726
rect 39116 14530 39172 14532
rect 39116 14478 39118 14530
rect 39118 14478 39170 14530
rect 39170 14478 39172 14530
rect 39116 14476 39172 14478
rect 39452 13692 39508 13748
rect 39004 13522 39060 13524
rect 39004 13470 39006 13522
rect 39006 13470 39058 13522
rect 39058 13470 39060 13522
rect 39004 13468 39060 13470
rect 40460 14642 40516 14644
rect 40460 14590 40462 14642
rect 40462 14590 40514 14642
rect 40514 14590 40516 14642
rect 40460 14588 40516 14590
rect 39900 13522 39956 13524
rect 39900 13470 39902 13522
rect 39902 13470 39954 13522
rect 39954 13470 39956 13522
rect 39900 13468 39956 13470
rect 40124 14476 40180 14532
rect 39340 12908 39396 12964
rect 38668 9826 38724 9828
rect 38668 9774 38670 9826
rect 38670 9774 38722 9826
rect 38722 9774 38724 9826
rect 38668 9772 38724 9774
rect 37772 9660 37828 9716
rect 38108 9714 38164 9716
rect 38108 9662 38110 9714
rect 38110 9662 38162 9714
rect 38162 9662 38164 9714
rect 38108 9660 38164 9662
rect 38332 9714 38388 9716
rect 38332 9662 38334 9714
rect 38334 9662 38386 9714
rect 38386 9662 38388 9714
rect 38332 9660 38388 9662
rect 37660 9212 37716 9268
rect 37212 9042 37268 9044
rect 37212 8990 37214 9042
rect 37214 8990 37266 9042
rect 37266 8990 37268 9042
rect 37212 8988 37268 8990
rect 38668 9266 38724 9268
rect 38668 9214 38670 9266
rect 38670 9214 38722 9266
rect 38722 9214 38724 9266
rect 38668 9212 38724 9214
rect 38444 9042 38500 9044
rect 38444 8990 38446 9042
rect 38446 8990 38498 9042
rect 38498 8990 38500 9042
rect 38444 8988 38500 8990
rect 35084 8258 35140 8260
rect 35084 8206 35086 8258
rect 35086 8206 35138 8258
rect 35138 8206 35140 8258
rect 35084 8204 35140 8206
rect 34972 7420 35028 7476
rect 35532 7420 35588 7476
rect 34412 6690 34468 6692
rect 34412 6638 34414 6690
rect 34414 6638 34466 6690
rect 34466 6638 34468 6690
rect 34412 6636 34468 6638
rect 33852 6524 33908 6580
rect 34636 6578 34692 6580
rect 34636 6526 34638 6578
rect 34638 6526 34690 6578
rect 34690 6526 34692 6578
rect 34636 6524 34692 6526
rect 33180 6130 33236 6132
rect 33180 6078 33182 6130
rect 33182 6078 33234 6130
rect 33234 6078 33236 6130
rect 33180 6076 33236 6078
rect 33852 6076 33908 6132
rect 33628 5852 33684 5908
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35420 6466 35476 6468
rect 35420 6414 35422 6466
rect 35422 6414 35474 6466
rect 35474 6414 35476 6466
rect 35420 6412 35476 6414
rect 36092 6748 36148 6804
rect 35532 5852 35588 5908
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5740 35700 5796
rect 36428 6076 36484 6132
rect 36764 6748 36820 6804
rect 36092 5906 36148 5908
rect 36092 5854 36094 5906
rect 36094 5854 36146 5906
rect 36146 5854 36148 5906
rect 36092 5852 36148 5854
rect 31500 4284 31556 4340
rect 37772 6748 37828 6804
rect 37324 6076 37380 6132
rect 37548 5964 37604 6020
rect 37436 5794 37492 5796
rect 37436 5742 37438 5794
rect 37438 5742 37490 5794
rect 37490 5742 37492 5794
rect 37436 5740 37492 5742
rect 38780 6748 38836 6804
rect 37884 6076 37940 6132
rect 37996 5740 38052 5796
rect 38892 6130 38948 6132
rect 38892 6078 38894 6130
rect 38894 6078 38946 6130
rect 38946 6078 38948 6130
rect 38892 6076 38948 6078
rect 38108 5010 38164 5012
rect 38108 4958 38110 5010
rect 38110 4958 38162 5010
rect 38162 4958 38164 5010
rect 38108 4956 38164 4958
rect 39340 9714 39396 9716
rect 39340 9662 39342 9714
rect 39342 9662 39394 9714
rect 39394 9662 39396 9714
rect 39340 9660 39396 9662
rect 39788 12962 39844 12964
rect 39788 12910 39790 12962
rect 39790 12910 39842 12962
rect 39842 12910 39844 12962
rect 39788 12908 39844 12910
rect 39900 12850 39956 12852
rect 39900 12798 39902 12850
rect 39902 12798 39954 12850
rect 39954 12798 39956 12850
rect 39900 12796 39956 12798
rect 40124 9548 40180 9604
rect 39004 5010 39060 5012
rect 39004 4958 39006 5010
rect 39006 4958 39058 5010
rect 39058 4958 39060 5010
rect 39004 4956 39060 4958
rect 39564 6130 39620 6132
rect 39564 6078 39566 6130
rect 39566 6078 39618 6130
rect 39618 6078 39620 6130
rect 39564 6076 39620 6078
rect 39452 4844 39508 4900
rect 40460 4844 40516 4900
rect 40236 4732 40292 4788
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 24892 3612 24948 3668
rect 41020 24668 41076 24724
rect 40908 23436 40964 23492
rect 41132 24780 41188 24836
rect 43036 32956 43092 33012
rect 42588 31836 42644 31892
rect 42476 31500 42532 31556
rect 42252 30770 42308 30772
rect 42252 30718 42254 30770
rect 42254 30718 42306 30770
rect 42306 30718 42308 30770
rect 42252 30716 42308 30718
rect 42364 30210 42420 30212
rect 42364 30158 42366 30210
rect 42366 30158 42418 30210
rect 42418 30158 42420 30210
rect 42364 30156 42420 30158
rect 42588 30156 42644 30212
rect 42700 29426 42756 29428
rect 42700 29374 42702 29426
rect 42702 29374 42754 29426
rect 42754 29374 42756 29426
rect 42700 29372 42756 29374
rect 42140 25282 42196 25284
rect 42140 25230 42142 25282
rect 42142 25230 42194 25282
rect 42194 25230 42196 25282
rect 42140 25228 42196 25230
rect 41692 24780 41748 24836
rect 41916 24780 41972 24836
rect 41580 24668 41636 24724
rect 41020 20300 41076 20356
rect 41020 19346 41076 19348
rect 41020 19294 41022 19346
rect 41022 19294 41074 19346
rect 41074 19294 41076 19346
rect 41020 19292 41076 19294
rect 40908 19234 40964 19236
rect 40908 19182 40910 19234
rect 40910 19182 40962 19234
rect 40962 19182 40964 19234
rect 40908 19180 40964 19182
rect 40908 14642 40964 14644
rect 40908 14590 40910 14642
rect 40910 14590 40962 14642
rect 40962 14590 40964 14642
rect 40908 14588 40964 14590
rect 41132 14530 41188 14532
rect 41132 14478 41134 14530
rect 41134 14478 41186 14530
rect 41186 14478 41188 14530
rect 41132 14476 41188 14478
rect 41580 23436 41636 23492
rect 41468 22428 41524 22484
rect 42476 25228 42532 25284
rect 42588 24780 42644 24836
rect 42700 24556 42756 24612
rect 42700 23548 42756 23604
rect 42252 22482 42308 22484
rect 42252 22430 42254 22482
rect 42254 22430 42306 22482
rect 42306 22430 42308 22482
rect 42252 22428 42308 22430
rect 41580 19292 41636 19348
rect 41692 18508 41748 18564
rect 41580 17612 41636 17668
rect 41804 18284 41860 18340
rect 42700 21756 42756 21812
rect 43596 33346 43652 33348
rect 43596 33294 43598 33346
rect 43598 33294 43650 33346
rect 43650 33294 43652 33346
rect 43596 33292 43652 33294
rect 43484 30156 43540 30212
rect 43708 31836 43764 31892
rect 43484 29596 43540 29652
rect 43372 28812 43428 28868
rect 43484 28754 43540 28756
rect 43484 28702 43486 28754
rect 43486 28702 43538 28754
rect 43538 28702 43540 28754
rect 43484 28700 43540 28702
rect 43596 29372 43652 29428
rect 44380 42252 44436 42308
rect 46172 55244 46228 55300
rect 46060 54796 46116 54852
rect 45836 53564 45892 53620
rect 45500 48972 45556 49028
rect 45612 50204 45668 50260
rect 45164 47852 45220 47908
rect 45388 48130 45444 48132
rect 45388 48078 45390 48130
rect 45390 48078 45442 48130
rect 45442 48078 45444 48130
rect 45388 48076 45444 48078
rect 46284 54796 46340 54852
rect 46284 51324 46340 51380
rect 46844 57762 46900 57764
rect 46844 57710 46846 57762
rect 46846 57710 46898 57762
rect 46898 57710 46900 57762
rect 46844 57708 46900 57710
rect 46732 55970 46788 55972
rect 46732 55918 46734 55970
rect 46734 55918 46786 55970
rect 46786 55918 46788 55970
rect 46732 55916 46788 55918
rect 47068 55916 47124 55972
rect 46732 55356 46788 55412
rect 46732 54796 46788 54852
rect 46620 54124 46676 54180
rect 47068 55298 47124 55300
rect 47068 55246 47070 55298
rect 47070 55246 47122 55298
rect 47122 55246 47124 55298
rect 47068 55244 47124 55246
rect 47068 53676 47124 53732
rect 46956 53452 47012 53508
rect 46844 51324 46900 51380
rect 46284 49868 46340 49924
rect 46396 49756 46452 49812
rect 46732 48972 46788 49028
rect 45164 46002 45220 46004
rect 45164 45950 45166 46002
rect 45166 45950 45218 46002
rect 45218 45950 45220 46002
rect 45164 45948 45220 45950
rect 45052 44940 45108 44996
rect 45724 48076 45780 48132
rect 45724 44994 45780 44996
rect 45724 44942 45726 44994
rect 45726 44942 45778 44994
rect 45778 44942 45780 44994
rect 45724 44940 45780 44942
rect 45836 44882 45892 44884
rect 45836 44830 45838 44882
rect 45838 44830 45890 44882
rect 45890 44830 45892 44882
rect 45836 44828 45892 44830
rect 46620 47852 46676 47908
rect 46620 46898 46676 46900
rect 46620 46846 46622 46898
rect 46622 46846 46674 46898
rect 46674 46846 46676 46898
rect 46620 46844 46676 46846
rect 46956 49026 47012 49028
rect 46956 48974 46958 49026
rect 46958 48974 47010 49026
rect 47010 48974 47012 49026
rect 46956 48972 47012 48974
rect 47180 48466 47236 48468
rect 47180 48414 47182 48466
rect 47182 48414 47234 48466
rect 47234 48414 47236 48466
rect 47180 48412 47236 48414
rect 48188 77980 48244 78036
rect 48188 75570 48244 75572
rect 48188 75518 48190 75570
rect 48190 75518 48242 75570
rect 48242 75518 48244 75570
rect 48188 75516 48244 75518
rect 48188 73052 48244 73108
rect 48188 70588 48244 70644
rect 48188 68124 48244 68180
rect 48188 65660 48244 65716
rect 48188 63196 48244 63252
rect 48188 60732 48244 60788
rect 48076 58322 48132 58324
rect 48076 58270 48078 58322
rect 48078 58270 48130 58322
rect 48130 58270 48132 58322
rect 48076 58268 48132 58270
rect 48076 55804 48132 55860
rect 47404 53676 47460 53732
rect 48076 53618 48132 53620
rect 48076 53566 48078 53618
rect 48078 53566 48130 53618
rect 48130 53566 48132 53618
rect 48076 53564 48132 53566
rect 48076 50876 48132 50932
rect 47516 49810 47572 49812
rect 47516 49758 47518 49810
rect 47518 49758 47570 49810
rect 47570 49758 47572 49810
rect 47516 49756 47572 49758
rect 47292 48188 47348 48244
rect 46956 46844 47012 46900
rect 45948 44434 46004 44436
rect 45948 44382 45950 44434
rect 45950 44382 46002 44434
rect 46002 44382 46004 44434
rect 45948 44380 46004 44382
rect 46508 44828 46564 44884
rect 45276 43426 45332 43428
rect 45276 43374 45278 43426
rect 45278 43374 45330 43426
rect 45330 43374 45332 43426
rect 45276 43372 45332 43374
rect 46620 43708 46676 43764
rect 47068 44380 47124 44436
rect 46620 43538 46676 43540
rect 46620 43486 46622 43538
rect 46622 43486 46674 43538
rect 46674 43486 46676 43538
rect 46620 43484 46676 43486
rect 46508 43372 46564 43428
rect 45836 42140 45892 42196
rect 44940 41916 44996 41972
rect 45724 41746 45780 41748
rect 45724 41694 45726 41746
rect 45726 41694 45778 41746
rect 45778 41694 45780 41746
rect 45724 41692 45780 41694
rect 45388 41020 45444 41076
rect 45164 40796 45220 40852
rect 44492 40514 44548 40516
rect 44492 40462 44494 40514
rect 44494 40462 44546 40514
rect 44546 40462 44548 40514
rect 44492 40460 44548 40462
rect 45388 40460 45444 40516
rect 44380 39788 44436 39844
rect 44492 39564 44548 39620
rect 47180 43538 47236 43540
rect 47180 43486 47182 43538
rect 47182 43486 47234 43538
rect 47234 43486 47236 43538
rect 47180 43484 47236 43486
rect 46172 41692 46228 41748
rect 46396 42028 46452 42084
rect 46172 41074 46228 41076
rect 46172 41022 46174 41074
rect 46174 41022 46226 41074
rect 46226 41022 46228 41074
rect 46172 41020 46228 41022
rect 44044 32844 44100 32900
rect 43932 29596 43988 29652
rect 43932 29426 43988 29428
rect 43932 29374 43934 29426
rect 43934 29374 43986 29426
rect 43986 29374 43988 29426
rect 43932 29372 43988 29374
rect 43708 28588 43764 28644
rect 42924 24722 42980 24724
rect 42924 24670 42926 24722
rect 42926 24670 42978 24722
rect 42978 24670 42980 24722
rect 42924 24668 42980 24670
rect 43148 24780 43204 24836
rect 43596 24668 43652 24724
rect 43036 24556 43092 24612
rect 42140 19292 42196 19348
rect 42028 17666 42084 17668
rect 42028 17614 42030 17666
rect 42030 17614 42082 17666
rect 42082 17614 42084 17666
rect 42028 17612 42084 17614
rect 43708 24556 43764 24612
rect 43820 24444 43876 24500
rect 43260 21756 43316 21812
rect 43036 16210 43092 16212
rect 43036 16158 43038 16210
rect 43038 16158 43090 16210
rect 43090 16158 43092 16210
rect 43036 16156 43092 16158
rect 43484 18284 43540 18340
rect 41692 12850 41748 12852
rect 41692 12798 41694 12850
rect 41694 12798 41746 12850
rect 41746 12798 41748 12850
rect 41692 12796 41748 12798
rect 41468 12066 41524 12068
rect 41468 12014 41470 12066
rect 41470 12014 41522 12066
rect 41522 12014 41524 12066
rect 41468 12012 41524 12014
rect 41692 11954 41748 11956
rect 41692 11902 41694 11954
rect 41694 11902 41746 11954
rect 41746 11902 41748 11954
rect 41692 11900 41748 11902
rect 42252 12796 42308 12852
rect 42364 12066 42420 12068
rect 42364 12014 42366 12066
rect 42366 12014 42418 12066
rect 42418 12014 42420 12066
rect 42364 12012 42420 12014
rect 42588 11954 42644 11956
rect 42588 11902 42590 11954
rect 42590 11902 42642 11954
rect 42642 11902 42644 11954
rect 42588 11900 42644 11902
rect 40908 9602 40964 9604
rect 40908 9550 40910 9602
rect 40910 9550 40962 9602
rect 40962 9550 40964 9602
rect 40908 9548 40964 9550
rect 43708 15820 43764 15876
rect 43596 14588 43652 14644
rect 43484 14476 43540 14532
rect 43260 13074 43316 13076
rect 43260 13022 43262 13074
rect 43262 13022 43314 13074
rect 43314 13022 43316 13074
rect 43260 13020 43316 13022
rect 44268 37378 44324 37380
rect 44268 37326 44270 37378
rect 44270 37326 44322 37378
rect 44322 37326 44324 37378
rect 44268 37324 44324 37326
rect 45836 39340 45892 39396
rect 44828 37324 44884 37380
rect 45612 36482 45668 36484
rect 45612 36430 45614 36482
rect 45614 36430 45666 36482
rect 45666 36430 45668 36482
rect 45612 36428 45668 36430
rect 45612 35532 45668 35588
rect 46060 37548 46116 37604
rect 46060 37212 46116 37268
rect 45948 36988 46004 37044
rect 46508 41916 46564 41972
rect 46172 36482 46228 36484
rect 46172 36430 46174 36482
rect 46174 36430 46226 36482
rect 46226 36430 46228 36482
rect 46172 36428 46228 36430
rect 45052 34242 45108 34244
rect 45052 34190 45054 34242
rect 45054 34190 45106 34242
rect 45106 34190 45108 34242
rect 45052 34188 45108 34190
rect 45724 34242 45780 34244
rect 45724 34190 45726 34242
rect 45726 34190 45778 34242
rect 45778 34190 45780 34242
rect 45724 34188 45780 34190
rect 44380 30380 44436 30436
rect 44604 29596 44660 29652
rect 46172 35532 46228 35588
rect 46284 34524 46340 34580
rect 47404 43596 47460 43652
rect 46620 36428 46676 36484
rect 46844 37548 46900 37604
rect 46844 37266 46900 37268
rect 46844 37214 46846 37266
rect 46846 37214 46898 37266
rect 46898 37214 46900 37266
rect 46844 37212 46900 37214
rect 46620 34412 46676 34468
rect 46508 34076 46564 34132
rect 46172 33346 46228 33348
rect 46172 33294 46174 33346
rect 46174 33294 46226 33346
rect 46226 33294 46228 33346
rect 46172 33292 46228 33294
rect 46620 33852 46676 33908
rect 46508 33292 46564 33348
rect 47068 34300 47124 34356
rect 45724 30156 45780 30212
rect 45164 28812 45220 28868
rect 45276 28754 45332 28756
rect 45276 28702 45278 28754
rect 45278 28702 45330 28754
rect 45330 28702 45332 28754
rect 45276 28700 45332 28702
rect 45388 28530 45444 28532
rect 45388 28478 45390 28530
rect 45390 28478 45442 28530
rect 45442 28478 45444 28530
rect 45388 28476 45444 28478
rect 45164 26908 45220 26964
rect 44156 26178 44212 26180
rect 44156 26126 44158 26178
rect 44158 26126 44210 26178
rect 44210 26126 44212 26178
rect 44156 26124 44212 26126
rect 44828 26178 44884 26180
rect 44828 26126 44830 26178
rect 44830 26126 44882 26178
rect 44882 26126 44884 26178
rect 44828 26124 44884 26126
rect 45164 26124 45220 26180
rect 44044 26012 44100 26068
rect 44044 24722 44100 24724
rect 44044 24670 44046 24722
rect 44046 24670 44098 24722
rect 44098 24670 44100 24722
rect 44044 24668 44100 24670
rect 44828 24668 44884 24724
rect 45388 25618 45444 25620
rect 45388 25566 45390 25618
rect 45390 25566 45442 25618
rect 45442 25566 45444 25618
rect 45388 25564 45444 25566
rect 45388 24722 45444 24724
rect 45388 24670 45390 24722
rect 45390 24670 45442 24722
rect 45442 24670 45444 24722
rect 45388 24668 45444 24670
rect 45052 24444 45108 24500
rect 44940 23996 44996 24052
rect 44828 20690 44884 20692
rect 44828 20638 44830 20690
rect 44830 20638 44882 20690
rect 44882 20638 44884 20690
rect 44828 20636 44884 20638
rect 44492 19404 44548 19460
rect 45724 26962 45780 26964
rect 45724 26910 45726 26962
rect 45726 26910 45778 26962
rect 45778 26910 45780 26962
rect 45724 26908 45780 26910
rect 46060 32674 46116 32676
rect 46060 32622 46062 32674
rect 46062 32622 46114 32674
rect 46114 32622 46116 32674
rect 46060 32620 46116 32622
rect 46732 32620 46788 32676
rect 47068 33740 47124 33796
rect 47292 33906 47348 33908
rect 47292 33854 47294 33906
rect 47294 33854 47346 33906
rect 47346 33854 47348 33906
rect 47292 33852 47348 33854
rect 47740 49922 47796 49924
rect 47740 49870 47742 49922
rect 47742 49870 47794 49922
rect 47794 49870 47796 49922
rect 47740 49868 47796 49870
rect 47964 49756 48020 49812
rect 47740 48802 47796 48804
rect 47740 48750 47742 48802
rect 47742 48750 47794 48802
rect 47794 48750 47796 48802
rect 47740 48748 47796 48750
rect 47740 48354 47796 48356
rect 47740 48302 47742 48354
rect 47742 48302 47794 48354
rect 47794 48302 47796 48354
rect 47740 48300 47796 48302
rect 47740 43708 47796 43764
rect 48076 45948 48132 46004
rect 48076 41074 48132 41076
rect 48076 41022 48078 41074
rect 48078 41022 48130 41074
rect 48130 41022 48132 41074
rect 48076 41020 48132 41022
rect 48188 38668 48244 38724
rect 47852 36988 47908 37044
rect 48188 36092 48244 36148
rect 47740 34412 47796 34468
rect 47628 33740 47684 33796
rect 48188 33628 48244 33684
rect 48300 33740 48356 33796
rect 46284 31836 46340 31892
rect 45948 28812 46004 28868
rect 47516 31836 47572 31892
rect 47180 29596 47236 29652
rect 48188 31164 48244 31220
rect 46620 28754 46676 28756
rect 46620 28702 46622 28754
rect 46622 28702 46674 28754
rect 46674 28702 46676 28754
rect 46620 28700 46676 28702
rect 48188 28530 48244 28532
rect 48188 28478 48190 28530
rect 48190 28478 48242 28530
rect 48242 28478 48244 28530
rect 48188 28476 48244 28478
rect 46620 26460 46676 26516
rect 47404 26460 47460 26516
rect 46732 26236 46788 26292
rect 46284 25564 46340 25620
rect 46396 25506 46452 25508
rect 46396 25454 46398 25506
rect 46398 25454 46450 25506
rect 46450 25454 46452 25506
rect 46396 25452 46452 25454
rect 46620 25452 46676 25508
rect 46508 25340 46564 25396
rect 45388 22988 45444 23044
rect 45276 22092 45332 22148
rect 45500 23324 45556 23380
rect 45836 23378 45892 23380
rect 45836 23326 45838 23378
rect 45838 23326 45890 23378
rect 45890 23326 45892 23378
rect 45836 23324 45892 23326
rect 45388 21868 45444 21924
rect 45948 22204 46004 22260
rect 44604 19180 44660 19236
rect 44044 14530 44100 14532
rect 44044 14478 44046 14530
rect 44046 14478 44098 14530
rect 44098 14478 44100 14530
rect 44044 14476 44100 14478
rect 44268 14530 44324 14532
rect 44268 14478 44270 14530
rect 44270 14478 44322 14530
rect 44322 14478 44324 14530
rect 44268 14476 44324 14478
rect 43932 13804 43988 13860
rect 43484 10668 43540 10724
rect 43260 10610 43316 10612
rect 43260 10558 43262 10610
rect 43262 10558 43314 10610
rect 43314 10558 43316 10610
rect 43260 10556 43316 10558
rect 44380 10722 44436 10724
rect 44380 10670 44382 10722
rect 44382 10670 44434 10722
rect 44434 10670 44436 10722
rect 44380 10668 44436 10670
rect 44044 10610 44100 10612
rect 44044 10558 44046 10610
rect 44046 10558 44098 10610
rect 44098 10558 44100 10610
rect 44044 10556 44100 10558
rect 42140 9826 42196 9828
rect 42140 9774 42142 9826
rect 42142 9774 42194 9826
rect 42194 9774 42196 9826
rect 42140 9772 42196 9774
rect 41132 8146 41188 8148
rect 41132 8094 41134 8146
rect 41134 8094 41186 8146
rect 41186 8094 41188 8146
rect 41132 8092 41188 8094
rect 40908 5964 40964 6020
rect 41916 7474 41972 7476
rect 41916 7422 41918 7474
rect 41918 7422 41970 7474
rect 41970 7422 41972 7474
rect 41916 7420 41972 7422
rect 41468 7196 41524 7252
rect 42812 10108 42868 10164
rect 42924 9772 42980 9828
rect 43372 9042 43428 9044
rect 43372 8990 43374 9042
rect 43374 8990 43426 9042
rect 43426 8990 43428 9042
rect 43372 8988 43428 8990
rect 44044 10108 44100 10164
rect 45388 19234 45444 19236
rect 45388 19182 45390 19234
rect 45390 19182 45442 19234
rect 45442 19182 45444 19234
rect 45388 19180 45444 19182
rect 42476 7420 42532 7476
rect 42812 7196 42868 7252
rect 41580 6018 41636 6020
rect 41580 5966 41582 6018
rect 41582 5966 41634 6018
rect 41634 5966 41636 6018
rect 41580 5964 41636 5966
rect 42364 5964 42420 6020
rect 44044 9042 44100 9044
rect 44044 8990 44046 9042
rect 44046 8990 44098 9042
rect 44098 8990 44100 9042
rect 44044 8988 44100 8990
rect 41132 4956 41188 5012
rect 44828 16156 44884 16212
rect 45052 15708 45108 15764
rect 45724 15874 45780 15876
rect 45724 15822 45726 15874
rect 45726 15822 45778 15874
rect 45778 15822 45780 15874
rect 45724 15820 45780 15822
rect 45500 15708 45556 15764
rect 44828 14642 44884 14644
rect 44828 14590 44830 14642
rect 44830 14590 44882 14642
rect 44882 14590 44884 14642
rect 44828 14588 44884 14590
rect 45388 14530 45444 14532
rect 45388 14478 45390 14530
rect 45390 14478 45442 14530
rect 45442 14478 45444 14530
rect 45388 14476 45444 14478
rect 45052 13020 45108 13076
rect 44604 4732 44660 4788
rect 45276 4060 45332 4116
rect 40684 3612 40740 3668
rect 44044 3666 44100 3668
rect 44044 3614 44046 3666
rect 44046 3614 44098 3666
rect 44098 3614 44100 3666
rect 44044 3612 44100 3614
rect 26908 3554 26964 3556
rect 26908 3502 26910 3554
rect 26910 3502 26962 3554
rect 26962 3502 26964 3554
rect 26908 3500 26964 3502
rect 21532 3388 21588 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 46172 23324 46228 23380
rect 46172 22370 46228 22372
rect 46172 22318 46174 22370
rect 46174 22318 46226 22370
rect 46226 22318 46228 22370
rect 46172 22316 46228 22318
rect 46396 21868 46452 21924
rect 48188 26236 48244 26292
rect 46732 24108 46788 24164
rect 48076 23826 48132 23828
rect 48076 23774 48078 23826
rect 48078 23774 48130 23826
rect 48130 23774 48132 23826
rect 48076 23772 48132 23774
rect 47068 22316 47124 22372
rect 46844 22258 46900 22260
rect 46844 22206 46846 22258
rect 46846 22206 46898 22258
rect 46898 22206 46900 22258
rect 46844 22204 46900 22206
rect 46956 22146 47012 22148
rect 46956 22094 46958 22146
rect 46958 22094 47010 22146
rect 47010 22094 47012 22146
rect 46956 22092 47012 22094
rect 48076 21308 48132 21364
rect 46732 20802 46788 20804
rect 46732 20750 46734 20802
rect 46734 20750 46786 20802
rect 46786 20750 46788 20802
rect 46732 20748 46788 20750
rect 47180 19906 47236 19908
rect 47180 19854 47182 19906
rect 47182 19854 47234 19906
rect 47234 19854 47236 19906
rect 47180 19852 47236 19854
rect 47628 19852 47684 19908
rect 48076 19122 48132 19124
rect 48076 19070 48078 19122
rect 48078 19070 48130 19122
rect 48130 19070 48132 19122
rect 48076 19068 48132 19070
rect 47068 18844 47124 18900
rect 47068 16210 47124 16212
rect 47068 16158 47070 16210
rect 47070 16158 47122 16210
rect 47122 16158 47124 16210
rect 47068 16156 47124 16158
rect 47740 16380 47796 16436
rect 47628 16156 47684 16212
rect 46732 14700 46788 14756
rect 48076 13916 48132 13972
rect 46620 13804 46676 13860
rect 46732 12178 46788 12180
rect 46732 12126 46734 12178
rect 46734 12126 46786 12178
rect 46786 12126 46788 12178
rect 46732 12124 46788 12126
rect 47740 11452 47796 11508
rect 46732 9938 46788 9940
rect 46732 9886 46734 9938
rect 46734 9886 46786 9938
rect 46786 9886 46788 9938
rect 46732 9884 46788 9886
rect 48076 8988 48132 9044
rect 48076 6578 48132 6580
rect 48076 6526 48078 6578
rect 48078 6526 48130 6578
rect 48130 6526 48132 6578
rect 48076 6524 48132 6526
rect 46620 4450 46676 4452
rect 46620 4398 46622 4450
rect 46622 4398 46674 4450
rect 46674 4398 46676 4450
rect 46620 4396 46676 4398
rect 46060 3500 46116 3556
rect 31164 3330 31220 3332
rect 31164 3278 31166 3330
rect 31166 3278 31218 3330
rect 31218 3278 31220 3330
rect 31164 3276 31220 3278
rect 48076 4060 48132 4116
rect 47740 1596 47796 1652
<< metal3 >>
rect 0 78036 800 78064
rect 49200 78036 50000 78064
rect 0 77980 2604 78036
rect 2660 77980 2670 78036
rect 48178 77980 48188 78036
rect 48244 77980 50000 78036
rect 0 77952 800 77980
rect 49200 77952 50000 77980
rect 29362 77196 29372 77252
rect 29428 77196 30380 77252
rect 30436 77196 30446 77252
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 13234 76636 13244 76692
rect 13300 76636 13916 76692
rect 13972 76636 13982 76692
rect 27570 76636 27580 76692
rect 27636 76636 29260 76692
rect 29316 76636 29326 76692
rect 31154 76636 31164 76692
rect 31220 76636 32620 76692
rect 32676 76636 32686 76692
rect 36866 76636 36876 76692
rect 36932 76636 37548 76692
rect 37604 76636 37614 76692
rect 42354 76636 42364 76692
rect 42420 76636 42924 76692
rect 42980 76636 42990 76692
rect 24322 76524 24332 76580
rect 24388 76524 33236 76580
rect 35074 76524 35084 76580
rect 35140 76524 36092 76580
rect 36148 76524 36158 76580
rect 40114 76524 40124 76580
rect 40180 76524 40796 76580
rect 40852 76524 41468 76580
rect 41524 76524 41534 76580
rect 1922 76412 1932 76468
rect 1988 76412 3724 76468
rect 3780 76412 3790 76468
rect 13570 76412 13580 76468
rect 13636 76412 15148 76468
rect 15204 76412 15214 76468
rect 27234 76412 27244 76468
rect 27300 76412 29148 76468
rect 29204 76412 29214 76468
rect 31154 76412 31164 76468
rect 31220 76412 32396 76468
rect 32452 76412 32462 76468
rect 33180 76356 33236 76524
rect 33394 76412 33404 76468
rect 33460 76412 34748 76468
rect 34804 76412 34814 76468
rect 43652 76356 43708 76468
rect 43764 76412 43774 76468
rect 20066 76300 20076 76356
rect 20132 76300 22092 76356
rect 22148 76300 22158 76356
rect 33180 76300 43708 76356
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 24770 75852 24780 75908
rect 24836 75852 38332 75908
rect 38388 75852 38398 75908
rect 2594 75740 2604 75796
rect 2660 75740 3612 75796
rect 3668 75740 3678 75796
rect 19058 75740 19068 75796
rect 19124 75740 20076 75796
rect 20132 75740 40012 75796
rect 40068 75740 40078 75796
rect 3154 75628 3164 75684
rect 3220 75628 5180 75684
rect 5236 75628 5246 75684
rect 14690 75628 14700 75684
rect 14756 75628 15932 75684
rect 15988 75628 15998 75684
rect 20626 75628 20636 75684
rect 20692 75628 22428 75684
rect 22484 75628 22494 75684
rect 29250 75628 29260 75684
rect 29316 75628 29596 75684
rect 29652 75628 31500 75684
rect 31556 75628 31948 75684
rect 32004 75628 32014 75684
rect 0 75572 800 75600
rect 49200 75572 50000 75600
rect 0 75516 1708 75572
rect 1764 75516 1774 75572
rect 48178 75516 48188 75572
rect 48244 75516 50000 75572
rect 0 75488 800 75516
rect 49200 75488 50000 75516
rect 19068 75404 20524 75460
rect 20580 75404 20590 75460
rect 19068 75236 19124 75404
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 19058 75180 19068 75236
rect 19124 75180 19134 75236
rect 5394 74956 5404 75012
rect 5460 74956 6636 75012
rect 6692 74956 9100 75012
rect 9156 74956 44380 75012
rect 44436 74956 44446 75012
rect 4162 74844 4172 74900
rect 4228 74844 4844 74900
rect 4900 74844 5740 74900
rect 5796 74844 5806 74900
rect 23538 74844 23548 74900
rect 23604 74844 23996 74900
rect 24052 74844 24668 74900
rect 24724 74844 26012 74900
rect 26068 74844 29596 74900
rect 29652 74844 29662 74900
rect 9090 74732 9100 74788
rect 9156 74732 9660 74788
rect 9716 74732 10668 74788
rect 10724 74732 10734 74788
rect 18162 74732 18172 74788
rect 18228 74732 19404 74788
rect 19460 74732 19470 74788
rect 22754 74732 22764 74788
rect 22820 74732 27244 74788
rect 27300 74732 27310 74788
rect 28578 74732 28588 74788
rect 28644 74732 31276 74788
rect 31332 74732 31342 74788
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 22754 74396 22764 74452
rect 22820 74396 24332 74452
rect 24388 74396 24398 74452
rect 15586 74284 15596 74340
rect 15652 74284 26348 74340
rect 26404 74284 26414 74340
rect 18162 74172 18172 74228
rect 18228 74172 19180 74228
rect 19236 74172 19246 74228
rect 20514 74172 20524 74228
rect 20580 74172 22316 74228
rect 22372 74172 23212 74228
rect 23268 74172 23278 74228
rect 23874 74172 23884 74228
rect 23940 74172 25228 74228
rect 25284 74172 25294 74228
rect 8372 74060 9100 74116
rect 9156 74060 9166 74116
rect 3938 73948 3948 74004
rect 4004 73948 4732 74004
rect 4788 73948 4798 74004
rect 5730 73948 5740 74004
rect 5796 73948 7588 74004
rect 7532 73892 7588 73948
rect 8372 73892 8428 74060
rect 10882 73948 10892 74004
rect 10948 73948 12460 74004
rect 12516 73948 14028 74004
rect 14084 73948 16380 74004
rect 16436 73948 16828 74004
rect 16884 73948 17388 74004
rect 17444 73948 19068 74004
rect 19124 73948 19134 74004
rect 19730 73948 19740 74004
rect 19796 73948 20748 74004
rect 20804 73948 20814 74004
rect 40338 73948 40348 74004
rect 40404 73948 45500 74004
rect 45556 73948 45566 74004
rect 7532 73836 8428 73892
rect 7532 73780 7588 73836
rect 7522 73724 7532 73780
rect 7588 73724 7598 73780
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 20626 73612 20636 73668
rect 20692 73612 33964 73668
rect 34020 73612 34030 73668
rect 26674 73500 26684 73556
rect 26740 73500 27692 73556
rect 27748 73500 27758 73556
rect 8306 73388 8316 73444
rect 8372 73388 9548 73444
rect 9604 73388 9614 73444
rect 11778 73388 11788 73444
rect 11844 73388 25452 73444
rect 25508 73388 25518 73444
rect 17938 73276 17948 73332
rect 18004 73276 18620 73332
rect 18676 73276 18686 73332
rect 18946 73276 18956 73332
rect 19012 73276 24780 73332
rect 24836 73276 24846 73332
rect 4834 73164 4844 73220
rect 4900 73164 5628 73220
rect 5684 73164 5694 73220
rect 16594 73164 16604 73220
rect 16660 73164 17164 73220
rect 17220 73164 17612 73220
rect 17668 73164 17678 73220
rect 26226 73164 26236 73220
rect 26292 73164 36540 73220
rect 36596 73164 36606 73220
rect 0 73108 800 73136
rect 49200 73108 50000 73136
rect 0 73052 1708 73108
rect 1764 73052 1774 73108
rect 24882 73052 24892 73108
rect 24948 73052 26684 73108
rect 26740 73052 26750 73108
rect 48178 73052 48188 73108
rect 48244 73052 50000 73108
rect 0 73024 800 73052
rect 49200 73024 50000 73052
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 18834 72828 18844 72884
rect 18900 72828 20748 72884
rect 20804 72828 20814 72884
rect 18162 72604 18172 72660
rect 18228 72604 18956 72660
rect 19012 72604 19180 72660
rect 19236 72604 19246 72660
rect 24546 72604 24556 72660
rect 24612 72604 25676 72660
rect 25732 72604 34300 72660
rect 34356 72604 34366 72660
rect 1250 72380 1260 72436
rect 1316 72380 5852 72436
rect 5908 72380 6524 72436
rect 6580 72380 6590 72436
rect 12786 72380 12796 72436
rect 12852 72380 21644 72436
rect 21700 72380 22204 72436
rect 22260 72380 22270 72436
rect 12898 72268 12908 72324
rect 12964 72268 17948 72324
rect 18004 72268 18014 72324
rect 23874 72268 23884 72324
rect 23940 72268 25340 72324
rect 25396 72268 26236 72324
rect 26292 72268 26302 72324
rect 32732 72268 33852 72324
rect 33908 72268 33918 72324
rect 36988 72268 42028 72324
rect 42084 72268 42094 72324
rect 32732 72212 32788 72268
rect 32722 72156 32732 72212
rect 32788 72156 32798 72212
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 28018 72044 28028 72100
rect 28084 72044 28364 72100
rect 28420 72044 28430 72100
rect 31154 71932 31164 71988
rect 31220 71932 31948 71988
rect 32004 71932 32014 71988
rect 28130 71820 28140 71876
rect 28196 71820 28476 71876
rect 28532 71820 28542 71876
rect 29810 71820 29820 71876
rect 29876 71820 30492 71876
rect 30548 71820 30558 71876
rect 36988 71764 37044 72268
rect 22418 71708 22428 71764
rect 22484 71708 22764 71764
rect 22820 71708 24332 71764
rect 24388 71708 37044 71764
rect 34962 71596 34972 71652
rect 35028 71596 37324 71652
rect 37380 71596 37996 71652
rect 38052 71596 38062 71652
rect 2146 71484 2156 71540
rect 2212 71484 4956 71540
rect 5012 71484 5022 71540
rect 3378 71372 3388 71428
rect 3444 71372 4284 71428
rect 4340 71372 4350 71428
rect 16594 71372 16604 71428
rect 16660 71372 17724 71428
rect 17780 71372 21980 71428
rect 22036 71372 22046 71428
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 11106 71260 11116 71316
rect 11172 71260 16716 71316
rect 16772 71260 16782 71316
rect 17042 71260 17052 71316
rect 17108 71260 22652 71316
rect 22708 71260 22718 71316
rect 8418 71148 8428 71204
rect 8484 71148 9212 71204
rect 9268 71148 23156 71204
rect 23100 71092 23156 71148
rect 31892 71148 35868 71204
rect 35924 71148 35934 71204
rect 4274 71036 4284 71092
rect 4340 71036 6300 71092
rect 6356 71036 6366 71092
rect 23090 71036 23100 71092
rect 23156 71036 23166 71092
rect 31892 70980 31948 71148
rect 34066 71036 34076 71092
rect 34132 71036 34860 71092
rect 34916 71036 35532 71092
rect 35588 71036 35598 71092
rect 25890 70924 25900 70980
rect 25956 70924 26908 70980
rect 26964 70924 26974 70980
rect 29922 70924 29932 70980
rect 29988 70924 30492 70980
rect 30548 70924 31948 70980
rect 11778 70812 11788 70868
rect 11844 70812 20524 70868
rect 20580 70812 20590 70868
rect 30930 70812 30940 70868
rect 30996 70812 35644 70868
rect 35700 70812 36988 70868
rect 37044 70812 37054 70868
rect 8194 70700 8204 70756
rect 8260 70700 18508 70756
rect 18564 70700 18574 70756
rect 21410 70700 21420 70756
rect 21476 70700 40348 70756
rect 40404 70700 40414 70756
rect 0 70644 800 70672
rect 8204 70644 8260 70700
rect 49200 70644 50000 70672
rect 0 70588 1708 70644
rect 1764 70588 1774 70644
rect 6748 70588 7084 70644
rect 7140 70588 8260 70644
rect 9874 70588 9884 70644
rect 9940 70588 11452 70644
rect 11508 70588 11518 70644
rect 15362 70588 15372 70644
rect 15428 70588 17164 70644
rect 17220 70588 17836 70644
rect 17892 70588 17902 70644
rect 18386 70588 18396 70644
rect 18452 70588 19404 70644
rect 19460 70588 19470 70644
rect 29372 70588 29596 70644
rect 29652 70588 30268 70644
rect 30324 70588 30334 70644
rect 33842 70588 33852 70644
rect 33908 70588 34076 70644
rect 34132 70588 35980 70644
rect 36036 70588 36046 70644
rect 48178 70588 48188 70644
rect 48244 70588 50000 70644
rect 0 70560 800 70588
rect 6748 70532 6804 70588
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 6178 70476 6188 70532
rect 6244 70476 6804 70532
rect 28242 70476 28252 70532
rect 28308 70476 29148 70532
rect 29204 70476 29214 70532
rect 29372 70420 29428 70588
rect 49200 70560 50000 70588
rect 37762 70476 37772 70532
rect 37828 70476 38892 70532
rect 38948 70476 38958 70532
rect 6514 70364 6524 70420
rect 6580 70364 7644 70420
rect 7700 70364 8428 70420
rect 8484 70364 8494 70420
rect 9986 70364 9996 70420
rect 10052 70364 10444 70420
rect 10500 70364 12460 70420
rect 12516 70364 13692 70420
rect 13748 70364 13758 70420
rect 18274 70364 18284 70420
rect 18340 70364 18732 70420
rect 18788 70364 21420 70420
rect 21476 70364 21486 70420
rect 29026 70364 29036 70420
rect 29092 70364 29428 70420
rect 8194 70252 8204 70308
rect 8260 70252 11788 70308
rect 11844 70252 11854 70308
rect 19282 70252 19292 70308
rect 19348 70252 20188 70308
rect 20244 70252 20254 70308
rect 27346 70252 27356 70308
rect 27412 70252 27804 70308
rect 27860 70252 41804 70308
rect 41860 70252 41870 70308
rect 10210 70140 10220 70196
rect 10276 70140 14140 70196
rect 14196 70140 14206 70196
rect 16258 70140 16268 70196
rect 16324 70140 25004 70196
rect 25060 70140 25070 70196
rect 37762 70140 37772 70196
rect 37828 70140 39004 70196
rect 39060 70140 39564 70196
rect 39620 70140 41692 70196
rect 41748 70140 41758 70196
rect 16818 70028 16828 70084
rect 16884 70028 17612 70084
rect 17668 70028 17678 70084
rect 25442 70028 25452 70084
rect 25508 70028 26908 70084
rect 36418 70028 36428 70084
rect 36484 70028 37660 70084
rect 37716 70028 37726 70084
rect 8418 69916 8428 69972
rect 8484 69916 23436 69972
rect 23492 69916 23502 69972
rect 26852 69860 26908 70028
rect 37986 69916 37996 69972
rect 38052 69916 38780 69972
rect 38836 69916 38846 69972
rect 26852 69804 27132 69860
rect 27188 69804 28028 69860
rect 28084 69804 29820 69860
rect 29876 69804 29886 69860
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 20626 69580 20636 69636
rect 20692 69580 21308 69636
rect 21364 69580 21374 69636
rect 25890 69580 25900 69636
rect 25956 69580 38444 69636
rect 38500 69580 38510 69636
rect 20636 69524 20692 69580
rect 12002 69468 12012 69524
rect 12068 69468 12796 69524
rect 12852 69468 20692 69524
rect 35634 69468 35644 69524
rect 35700 69468 39004 69524
rect 39060 69468 39070 69524
rect 6626 69244 6636 69300
rect 6692 69244 6972 69300
rect 7028 69244 8764 69300
rect 8820 69244 8830 69300
rect 36306 69244 36316 69300
rect 36372 69244 37324 69300
rect 37380 69244 37390 69300
rect 7046 69132 7084 69188
rect 7140 69132 7150 69188
rect 24210 69132 24220 69188
rect 24276 69132 24668 69188
rect 24724 69132 25676 69188
rect 25732 69132 25742 69188
rect 34962 69132 34972 69188
rect 35028 69132 35196 69188
rect 35252 69132 37772 69188
rect 37828 69132 37838 69188
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 6402 68908 6412 68964
rect 6468 68908 8540 68964
rect 8596 68908 8606 68964
rect 8754 68908 8764 68964
rect 8820 68908 9996 68964
rect 10052 68908 10062 68964
rect 33394 68684 33404 68740
rect 33460 68684 34300 68740
rect 34356 68684 34366 68740
rect 5842 68572 5852 68628
rect 5908 68572 6636 68628
rect 6692 68572 6702 68628
rect 8082 68572 8092 68628
rect 8148 68572 9548 68628
rect 9604 68572 9614 68628
rect 33058 68572 33068 68628
rect 33124 68572 34188 68628
rect 34244 68572 34254 68628
rect 38658 68572 38668 68628
rect 38724 68572 39228 68628
rect 39284 68572 39564 68628
rect 39620 68572 39630 68628
rect 32386 68460 32396 68516
rect 32452 68460 35196 68516
rect 35252 68460 35756 68516
rect 35812 68460 37436 68516
rect 37492 68460 37502 68516
rect 38770 68348 38780 68404
rect 38836 68348 40572 68404
rect 40628 68348 40638 68404
rect 0 68180 800 68208
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 49200 68180 50000 68208
rect 0 68124 1820 68180
rect 1876 68124 1886 68180
rect 48178 68124 48188 68180
rect 48244 68124 50000 68180
rect 0 68096 800 68124
rect 49200 68096 50000 68124
rect 7606 67900 7644 67956
rect 7700 67900 7710 67956
rect 29810 67788 29820 67844
rect 29876 67788 30940 67844
rect 30996 67788 31006 67844
rect 7522 67676 7532 67732
rect 7588 67676 8204 67732
rect 8260 67676 8270 67732
rect 32946 67676 32956 67732
rect 33012 67676 33404 67732
rect 33460 67676 34076 67732
rect 34132 67676 34142 67732
rect 40898 67676 40908 67732
rect 40964 67676 42252 67732
rect 42308 67676 43596 67732
rect 43652 67676 43662 67732
rect 6514 67564 6524 67620
rect 6580 67564 7756 67620
rect 7812 67564 7980 67620
rect 8036 67564 8046 67620
rect 14466 67564 14476 67620
rect 14532 67564 15260 67620
rect 15316 67564 15326 67620
rect 17378 67564 17388 67620
rect 17444 67564 19292 67620
rect 19348 67564 19358 67620
rect 31378 67564 31388 67620
rect 31444 67564 31724 67620
rect 31780 67564 32396 67620
rect 32452 67564 32462 67620
rect 23650 67452 23660 67508
rect 23716 67452 24444 67508
rect 24500 67452 24510 67508
rect 31042 67452 31052 67508
rect 31108 67452 35644 67508
rect 35700 67452 35710 67508
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 10658 67340 10668 67396
rect 10724 67340 11676 67396
rect 11732 67340 11742 67396
rect 6626 67228 6636 67284
rect 6692 67228 7756 67284
rect 7812 67228 7822 67284
rect 18162 67228 18172 67284
rect 18228 67228 19068 67284
rect 19124 67228 19134 67284
rect 17938 67116 17948 67172
rect 18004 67116 18620 67172
rect 18676 67116 21308 67172
rect 21364 67116 21374 67172
rect 23314 67116 23324 67172
rect 23380 67116 23996 67172
rect 24052 67116 24062 67172
rect 29250 67116 29260 67172
rect 29316 67116 29596 67172
rect 29652 67116 29662 67172
rect 14802 67004 14812 67060
rect 14868 67004 14878 67060
rect 26562 67004 26572 67060
rect 26628 67004 27356 67060
rect 27412 67004 27422 67060
rect 28354 67004 28364 67060
rect 28420 67004 29484 67060
rect 29540 67004 29550 67060
rect 35298 67004 35308 67060
rect 35364 67004 36316 67060
rect 36372 67004 36382 67060
rect 38994 67004 39004 67060
rect 39060 67004 39564 67060
rect 39620 67004 39630 67060
rect 42578 67004 42588 67060
rect 42644 67004 43372 67060
rect 43428 67004 44604 67060
rect 44660 67004 44670 67060
rect 14812 66948 14868 67004
rect 14812 66892 15932 66948
rect 15988 66892 17276 66948
rect 17332 66892 17500 66948
rect 17556 66892 17566 66948
rect 25442 66892 25452 66948
rect 25508 66892 26684 66948
rect 26740 66892 27692 66948
rect 27748 66892 27916 66948
rect 27972 66892 27982 66948
rect 27346 66780 27356 66836
rect 27412 66780 28588 66836
rect 28644 66780 29596 66836
rect 29652 66780 30604 66836
rect 30660 66780 30670 66836
rect 43250 66780 43260 66836
rect 43316 66780 44268 66836
rect 44324 66780 44334 66836
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 30604 66332 31836 66388
rect 31892 66332 31902 66388
rect 32162 66332 32172 66388
rect 32228 66332 34300 66388
rect 34356 66332 34366 66388
rect 37538 66332 37548 66388
rect 37604 66332 39116 66388
rect 39172 66332 39182 66388
rect 41346 66332 41356 66388
rect 41412 66332 42252 66388
rect 42308 66332 42318 66388
rect 30604 66276 30660 66332
rect 1586 66220 1596 66276
rect 1652 66220 2268 66276
rect 2324 66220 2334 66276
rect 6738 66220 6748 66276
rect 6804 66220 9436 66276
rect 9492 66220 10108 66276
rect 10164 66220 10174 66276
rect 15026 66220 15036 66276
rect 15092 66220 17388 66276
rect 17444 66220 17454 66276
rect 29474 66220 29484 66276
rect 29540 66220 29820 66276
rect 29876 66220 30604 66276
rect 30660 66220 30670 66276
rect 31266 66220 31276 66276
rect 31332 66220 32060 66276
rect 32116 66220 32844 66276
rect 32900 66220 32910 66276
rect 33394 66220 33404 66276
rect 33460 66220 34412 66276
rect 34468 66220 37436 66276
rect 37492 66220 37502 66276
rect 38322 66220 38332 66276
rect 38388 66220 39228 66276
rect 39284 66220 39294 66276
rect 12198 66108 12236 66164
rect 12292 66108 12302 66164
rect 21746 66108 21756 66164
rect 21812 66108 22428 66164
rect 22484 66108 22494 66164
rect 37538 66108 37548 66164
rect 37604 66108 38444 66164
rect 38500 66108 38510 66164
rect 5058 65996 5068 66052
rect 5124 65996 5628 66052
rect 5684 65996 5694 66052
rect 13906 65996 13916 66052
rect 13972 65996 15596 66052
rect 15652 65996 15662 66052
rect 29138 65996 29148 66052
rect 29204 65996 29932 66052
rect 29988 65996 31052 66052
rect 31108 65996 31118 66052
rect 40114 65996 40124 66052
rect 40180 65996 41020 66052
rect 41076 65996 41086 66052
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 5394 65772 5404 65828
rect 5460 65772 7308 65828
rect 7364 65772 7374 65828
rect 13010 65772 13020 65828
rect 13076 65772 14252 65828
rect 14308 65772 14924 65828
rect 14980 65772 14990 65828
rect 41906 65772 41916 65828
rect 41972 65772 42364 65828
rect 42420 65772 42430 65828
rect 0 65716 800 65744
rect 49200 65716 50000 65744
rect 0 65660 1820 65716
rect 1876 65660 1886 65716
rect 15026 65660 15036 65716
rect 15092 65660 17612 65716
rect 17668 65660 17678 65716
rect 32386 65660 32396 65716
rect 32452 65660 33740 65716
rect 33796 65660 33806 65716
rect 48178 65660 48188 65716
rect 48244 65660 50000 65716
rect 0 65632 800 65660
rect 49200 65632 50000 65660
rect 2146 65548 2156 65604
rect 2212 65548 4172 65604
rect 4228 65548 4238 65604
rect 7186 65548 7196 65604
rect 7252 65548 7644 65604
rect 7700 65548 7710 65604
rect 14130 65548 14140 65604
rect 14196 65548 15260 65604
rect 15316 65548 15326 65604
rect 31826 65548 31836 65604
rect 31892 65548 34524 65604
rect 34580 65548 34590 65604
rect 4386 65436 4396 65492
rect 4452 65436 8316 65492
rect 8372 65436 8382 65492
rect 11778 65436 11788 65492
rect 11844 65436 12572 65492
rect 12628 65436 12638 65492
rect 13570 65436 13580 65492
rect 13636 65436 14252 65492
rect 14308 65436 14318 65492
rect 14690 65436 14700 65492
rect 14756 65436 15596 65492
rect 15652 65436 15662 65492
rect 15820 65436 16492 65492
rect 16548 65436 16558 65492
rect 20850 65436 20860 65492
rect 20916 65436 22092 65492
rect 22148 65436 22158 65492
rect 32274 65436 32284 65492
rect 32340 65436 33628 65492
rect 33684 65436 33694 65492
rect 36866 65436 36876 65492
rect 36932 65436 37660 65492
rect 37716 65436 37726 65492
rect 15820 65380 15876 65436
rect 7746 65324 7756 65380
rect 7812 65324 8652 65380
rect 8708 65324 8718 65380
rect 10882 65324 10892 65380
rect 10948 65324 13468 65380
rect 13524 65324 15820 65380
rect 15876 65324 15886 65380
rect 16370 65324 16380 65380
rect 16436 65324 16446 65380
rect 20738 65324 20748 65380
rect 20804 65324 22988 65380
rect 23044 65324 23054 65380
rect 32498 65324 32508 65380
rect 32564 65324 33180 65380
rect 33236 65324 33246 65380
rect 37538 65324 37548 65380
rect 37604 65324 40572 65380
rect 40628 65324 41020 65380
rect 41076 65324 41356 65380
rect 41412 65324 41422 65380
rect 16380 65268 16436 65324
rect 6178 65212 6188 65268
rect 6244 65212 7644 65268
rect 7700 65212 7710 65268
rect 12338 65212 12348 65268
rect 12404 65212 12796 65268
rect 12852 65212 12862 65268
rect 14802 65212 14812 65268
rect 14868 65212 16436 65268
rect 18162 65212 18172 65268
rect 18228 65212 18844 65268
rect 18900 65212 18910 65268
rect 40002 65212 40012 65268
rect 40068 65212 40348 65268
rect 40404 65212 40908 65268
rect 40964 65212 40974 65268
rect 15586 65100 15596 65156
rect 15652 65100 17612 65156
rect 17668 65100 20188 65156
rect 20244 65100 21308 65156
rect 21364 65100 21374 65156
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 10882 64988 10892 65044
rect 10948 64988 10958 65044
rect 10892 64820 10948 64988
rect 11554 64876 11564 64932
rect 11620 64876 12012 64932
rect 12068 64876 12078 64932
rect 10770 64764 10780 64820
rect 10836 64764 10948 64820
rect 16706 64764 16716 64820
rect 16772 64764 25340 64820
rect 25396 64764 25406 64820
rect 27794 64764 27804 64820
rect 27860 64764 31948 64820
rect 34402 64764 34412 64820
rect 34468 64764 35420 64820
rect 35476 64764 35486 64820
rect 37874 64764 37884 64820
rect 37940 64764 38668 64820
rect 38724 64764 38734 64820
rect 31892 64708 31948 64764
rect 6738 64652 6748 64708
rect 6804 64652 7196 64708
rect 7252 64652 7262 64708
rect 9538 64652 9548 64708
rect 9604 64652 10108 64708
rect 10164 64652 10668 64708
rect 10724 64652 10734 64708
rect 15138 64652 15148 64708
rect 15204 64652 16044 64708
rect 16100 64652 16110 64708
rect 20972 64652 22092 64708
rect 22148 64652 22158 64708
rect 31892 64652 41076 64708
rect 20972 64596 21028 64652
rect 41020 64596 41076 64652
rect 8754 64540 8764 64596
rect 8820 64540 10220 64596
rect 10276 64540 10286 64596
rect 11554 64540 11564 64596
rect 11620 64540 12572 64596
rect 12628 64540 12638 64596
rect 13906 64540 13916 64596
rect 13972 64540 14588 64596
rect 14644 64540 16268 64596
rect 16324 64540 16334 64596
rect 17266 64540 17276 64596
rect 17332 64540 18396 64596
rect 18452 64540 19740 64596
rect 19796 64540 20972 64596
rect 21028 64540 21038 64596
rect 21858 64540 21868 64596
rect 21924 64540 24556 64596
rect 24612 64540 24622 64596
rect 41010 64540 41020 64596
rect 41076 64540 41086 64596
rect 6514 64428 6524 64484
rect 6580 64428 7196 64484
rect 7252 64428 7262 64484
rect 15446 64428 15484 64484
rect 15540 64428 15550 64484
rect 17042 64428 17052 64484
rect 17108 64428 17612 64484
rect 17668 64428 17678 64484
rect 19506 64428 19516 64484
rect 19572 64428 20636 64484
rect 20692 64428 23660 64484
rect 23716 64428 23726 64484
rect 10322 64316 10332 64372
rect 10388 64316 11228 64372
rect 11284 64316 13020 64372
rect 13076 64316 13086 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 10546 64204 10556 64260
rect 10612 64204 11116 64260
rect 11172 64204 11182 64260
rect 11442 64204 11452 64260
rect 11508 64204 15148 64260
rect 15092 64148 15148 64204
rect 8978 64092 8988 64148
rect 9044 64092 9884 64148
rect 9940 64092 9950 64148
rect 12198 64092 12236 64148
rect 12292 64092 12302 64148
rect 15092 64092 26236 64148
rect 26292 64092 26302 64148
rect 39778 64092 39788 64148
rect 39844 64092 40684 64148
rect 40740 64092 40750 64148
rect 9884 63924 9940 64092
rect 10770 63980 10780 64036
rect 10836 63980 11788 64036
rect 11844 63980 13244 64036
rect 13300 63980 14252 64036
rect 14308 63980 14318 64036
rect 16034 63980 16044 64036
rect 16100 63980 16940 64036
rect 16996 63980 18396 64036
rect 18452 63980 18462 64036
rect 35746 63980 35756 64036
rect 35812 63980 36652 64036
rect 36708 63980 36718 64036
rect 9884 63868 13468 63924
rect 13524 63868 13916 63924
rect 13972 63868 13982 63924
rect 38770 63868 38780 63924
rect 38836 63868 39900 63924
rect 39956 63868 39966 63924
rect 10780 63812 10836 63868
rect 10770 63756 10780 63812
rect 10836 63756 10846 63812
rect 25778 63756 25788 63812
rect 25844 63756 26684 63812
rect 26740 63756 26750 63812
rect 29250 63756 29260 63812
rect 29316 63756 29932 63812
rect 29988 63756 30380 63812
rect 30436 63756 30446 63812
rect 34626 63756 34636 63812
rect 34692 63756 35196 63812
rect 35252 63756 36428 63812
rect 36484 63756 36494 63812
rect 37874 63756 37884 63812
rect 37940 63756 39004 63812
rect 39060 63756 39070 63812
rect 43474 63756 43484 63812
rect 43540 63756 45836 63812
rect 45892 63756 46060 63812
rect 46116 63756 46126 63812
rect 11890 63644 11900 63700
rect 11956 63644 15596 63700
rect 15652 63644 15662 63700
rect 18162 63644 18172 63700
rect 18228 63644 19068 63700
rect 19124 63644 19134 63700
rect 26562 63644 26572 63700
rect 26628 63644 27692 63700
rect 27748 63644 27758 63700
rect 30482 63644 30492 63700
rect 30548 63644 31164 63700
rect 31220 63644 31230 63700
rect 38210 63644 38220 63700
rect 38276 63644 39676 63700
rect 39732 63644 39742 63700
rect 41010 63644 41020 63700
rect 41076 63644 44268 63700
rect 44324 63644 44334 63700
rect 14914 63532 14924 63588
rect 14980 63532 18284 63588
rect 18340 63532 18350 63588
rect 25330 63532 25340 63588
rect 25396 63532 32284 63588
rect 32340 63532 32350 63588
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 17826 63308 17836 63364
rect 17892 63308 18172 63364
rect 18228 63308 19180 63364
rect 19236 63308 19964 63364
rect 20020 63308 20030 63364
rect 25442 63308 25452 63364
rect 25508 63308 27020 63364
rect 27076 63308 27086 63364
rect 30930 63308 30940 63364
rect 30996 63308 31948 63364
rect 32004 63308 32014 63364
rect 0 63252 800 63280
rect 49200 63252 50000 63280
rect 0 63196 1820 63252
rect 1876 63196 1886 63252
rect 6626 63196 6636 63252
rect 6692 63196 6972 63252
rect 7028 63196 7756 63252
rect 7812 63196 7822 63252
rect 13122 63196 13132 63252
rect 13188 63196 16828 63252
rect 16884 63196 16894 63252
rect 20290 63196 20300 63252
rect 20356 63196 21644 63252
rect 21700 63196 21710 63252
rect 45938 63196 45948 63252
rect 46004 63196 46844 63252
rect 46900 63196 46910 63252
rect 48178 63196 48188 63252
rect 48244 63196 50000 63252
rect 0 63168 800 63196
rect 49200 63168 50000 63196
rect 7158 63084 7196 63140
rect 7252 63084 7262 63140
rect 7606 63084 7644 63140
rect 7700 63084 7710 63140
rect 17266 63084 17276 63140
rect 17332 63084 18844 63140
rect 18900 63084 18910 63140
rect 26562 63084 26572 63140
rect 26628 63084 27356 63140
rect 27412 63084 28028 63140
rect 28084 63084 28094 63140
rect 34290 63084 34300 63140
rect 34356 63084 35420 63140
rect 35476 63084 35486 63140
rect 44930 63084 44940 63140
rect 44996 63084 45612 63140
rect 45668 63084 46620 63140
rect 46676 63084 46686 63140
rect 25330 62972 25340 63028
rect 25396 62972 26348 63028
rect 26404 62972 28924 63028
rect 28980 62972 29484 63028
rect 29540 62972 29550 63028
rect 33394 62972 33404 63028
rect 33460 62972 34188 63028
rect 34244 62972 35196 63028
rect 35252 62972 35262 63028
rect 6290 62860 6300 62916
rect 6356 62860 7196 62916
rect 7252 62860 7262 62916
rect 16370 62860 16380 62916
rect 16436 62860 16828 62916
rect 16884 62860 17500 62916
rect 17556 62860 17566 62916
rect 19394 62860 19404 62916
rect 19460 62860 19740 62916
rect 19796 62860 19806 62916
rect 21522 62860 21532 62916
rect 21588 62860 25676 62916
rect 25732 62860 25742 62916
rect 29362 62860 29372 62916
rect 29428 62860 30044 62916
rect 30100 62860 30110 62916
rect 42802 62860 42812 62916
rect 42868 62860 44268 62916
rect 44324 62860 44334 62916
rect 17826 62748 17836 62804
rect 17892 62748 18172 62804
rect 18228 62748 18238 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 2258 62636 2268 62692
rect 2324 62636 4620 62692
rect 4676 62636 4686 62692
rect 15250 62636 15260 62692
rect 15316 62636 16660 62692
rect 16604 62580 16660 62636
rect 21532 62580 21588 62860
rect 10434 62524 10444 62580
rect 10500 62524 11116 62580
rect 11172 62524 11452 62580
rect 11508 62524 14028 62580
rect 14084 62524 14094 62580
rect 14690 62524 14700 62580
rect 14756 62524 15932 62580
rect 15988 62524 15998 62580
rect 16594 62524 16604 62580
rect 16660 62524 21588 62580
rect 44034 62524 44044 62580
rect 44100 62524 44604 62580
rect 44660 62524 44670 62580
rect 1474 62412 1484 62468
rect 1540 62412 5740 62468
rect 5796 62412 5806 62468
rect 28018 62412 28028 62468
rect 28084 62412 43260 62468
rect 43316 62412 43326 62468
rect 6402 62300 6412 62356
rect 6468 62300 7196 62356
rect 7252 62300 7756 62356
rect 7812 62300 8204 62356
rect 8260 62300 8270 62356
rect 8642 62300 8652 62356
rect 8708 62300 14924 62356
rect 14980 62300 14990 62356
rect 15586 62300 15596 62356
rect 15652 62300 16044 62356
rect 16100 62300 16110 62356
rect 16706 62300 16716 62356
rect 16772 62300 17948 62356
rect 18004 62300 18014 62356
rect 30482 62300 30492 62356
rect 30548 62300 31388 62356
rect 31444 62300 31724 62356
rect 31780 62300 33180 62356
rect 33236 62300 33246 62356
rect 41682 62300 41692 62356
rect 41748 62300 42924 62356
rect 42980 62300 44044 62356
rect 44100 62300 44110 62356
rect 8204 62244 8260 62300
rect 8204 62188 8988 62244
rect 9044 62188 9054 62244
rect 10098 62188 10108 62244
rect 10164 62188 12908 62244
rect 12964 62188 12974 62244
rect 15362 62188 15372 62244
rect 15428 62188 18508 62244
rect 18564 62188 18574 62244
rect 18834 62188 18844 62244
rect 18900 62188 20300 62244
rect 20356 62188 20366 62244
rect 22866 62188 22876 62244
rect 22932 62188 23884 62244
rect 23940 62188 24668 62244
rect 24724 62188 24734 62244
rect 31154 62188 31164 62244
rect 31220 62188 32060 62244
rect 32116 62188 32126 62244
rect 12562 62076 12572 62132
rect 12628 62076 14924 62132
rect 14980 62076 14990 62132
rect 26674 62076 26684 62132
rect 26740 62076 27244 62132
rect 27300 62076 27310 62132
rect 29362 62076 29372 62132
rect 29428 62076 31724 62132
rect 31780 62076 31790 62132
rect 26450 61964 26460 62020
rect 26516 61964 26796 62020
rect 26852 61964 26862 62020
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 18498 61852 18508 61908
rect 18564 61852 19404 61908
rect 19460 61852 19470 61908
rect 7298 61740 7308 61796
rect 7364 61740 7868 61796
rect 7924 61740 8428 61796
rect 8484 61740 8494 61796
rect 20962 61628 20972 61684
rect 21028 61628 25340 61684
rect 25396 61628 27132 61684
rect 27188 61628 27198 61684
rect 29922 61628 29932 61684
rect 29988 61628 31612 61684
rect 31668 61628 31678 61684
rect 41906 61628 41916 61684
rect 41972 61628 42476 61684
rect 42532 61628 43036 61684
rect 43092 61628 43102 61684
rect 5170 61516 5180 61572
rect 5236 61516 5852 61572
rect 5908 61516 5918 61572
rect 6290 61516 6300 61572
rect 6356 61516 6366 61572
rect 11218 61516 11228 61572
rect 11284 61516 11788 61572
rect 11844 61516 11854 61572
rect 12674 61516 12684 61572
rect 12740 61516 14364 61572
rect 14420 61516 14430 61572
rect 15474 61516 15484 61572
rect 15540 61516 16492 61572
rect 16548 61516 16558 61572
rect 18918 61516 18956 61572
rect 19012 61516 19022 61572
rect 24434 61516 24444 61572
rect 24500 61516 24892 61572
rect 24948 61516 24958 61572
rect 41010 61516 41020 61572
rect 41076 61516 42140 61572
rect 42196 61516 43148 61572
rect 43204 61516 43214 61572
rect 6300 61460 6356 61516
rect 2930 61404 2940 61460
rect 2996 61404 4060 61460
rect 4116 61404 4126 61460
rect 5506 61404 5516 61460
rect 5572 61404 6356 61460
rect 13010 61404 13020 61460
rect 13076 61404 13692 61460
rect 13748 61404 13758 61460
rect 19506 61404 19516 61460
rect 19572 61404 21644 61460
rect 21700 61404 21710 61460
rect 31490 61404 31500 61460
rect 31556 61404 32620 61460
rect 32676 61404 32686 61460
rect 37762 61404 37772 61460
rect 37828 61404 39452 61460
rect 39508 61404 39518 61460
rect 43922 61404 43932 61460
rect 43988 61404 44940 61460
rect 44996 61404 45006 61460
rect 5730 61292 5740 61348
rect 5796 61292 6860 61348
rect 6916 61292 7196 61348
rect 7252 61292 7262 61348
rect 12002 61292 12012 61348
rect 12068 61292 13580 61348
rect 13636 61292 13646 61348
rect 13794 61292 13804 61348
rect 13860 61292 18844 61348
rect 18900 61292 19292 61348
rect 19348 61292 19358 61348
rect 20514 61292 20524 61348
rect 20580 61292 22652 61348
rect 22708 61292 22718 61348
rect 5842 61180 5852 61236
rect 5908 61180 6972 61236
rect 7028 61180 7038 61236
rect 11554 61180 11564 61236
rect 11620 61180 13468 61236
rect 13524 61180 13534 61236
rect 17154 61180 17164 61236
rect 17220 61180 17612 61236
rect 17668 61180 18620 61236
rect 18676 61180 19180 61236
rect 19236 61180 19516 61236
rect 19572 61180 19582 61236
rect 37090 61180 37100 61236
rect 37156 61180 37166 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 12786 61068 12796 61124
rect 12852 61068 14140 61124
rect 14196 61068 15372 61124
rect 15428 61068 15438 61124
rect 15586 61068 15596 61124
rect 15652 61068 15932 61124
rect 15988 61068 17892 61124
rect 19030 61068 19068 61124
rect 19124 61068 19134 61124
rect 17836 60900 17892 61068
rect 18050 60956 18060 61012
rect 18116 60956 20524 61012
rect 20580 60956 20590 61012
rect 31378 60956 31388 61012
rect 31444 60956 33180 61012
rect 33236 60956 36876 61012
rect 36932 60956 36942 61012
rect 14018 60844 14028 60900
rect 14084 60844 15932 60900
rect 15988 60844 15998 60900
rect 17836 60844 22372 60900
rect 22530 60844 22540 60900
rect 22596 60844 25228 60900
rect 25284 60844 25294 60900
rect 0 60788 800 60816
rect 22316 60788 22372 60844
rect 0 60732 1708 60788
rect 1764 60732 1774 60788
rect 5506 60732 5516 60788
rect 5572 60732 6636 60788
rect 6692 60732 9660 60788
rect 9716 60732 9726 60788
rect 15250 60732 15260 60788
rect 15316 60732 15596 60788
rect 15652 60732 15662 60788
rect 16482 60732 16492 60788
rect 16548 60732 18508 60788
rect 18564 60732 21756 60788
rect 21812 60732 21822 60788
rect 22316 60732 24108 60788
rect 24164 60732 24892 60788
rect 24948 60732 25564 60788
rect 25620 60732 25630 60788
rect 0 60704 800 60732
rect 31724 60676 31780 60956
rect 31938 60844 31948 60900
rect 32004 60844 33628 60900
rect 33684 60844 33694 60900
rect 34850 60844 34860 60900
rect 34916 60844 36764 60900
rect 36820 60844 36830 60900
rect 37100 60788 37156 61180
rect 41010 60956 41020 61012
rect 41076 60956 41916 61012
rect 41972 60956 41982 61012
rect 49200 60788 50000 60816
rect 32610 60732 32620 60788
rect 32676 60732 34748 60788
rect 34804 60732 34814 60788
rect 34962 60732 34972 60788
rect 35028 60732 35756 60788
rect 35812 60732 35822 60788
rect 36306 60732 36316 60788
rect 36372 60732 37212 60788
rect 37268 60732 37278 60788
rect 40002 60732 40012 60788
rect 40068 60732 41132 60788
rect 41188 60732 41468 60788
rect 41524 60732 41534 60788
rect 48178 60732 48188 60788
rect 48244 60732 50000 60788
rect 49200 60704 50000 60732
rect 14802 60620 14812 60676
rect 14868 60620 17612 60676
rect 17668 60620 17836 60676
rect 17892 60620 17902 60676
rect 19170 60620 19180 60676
rect 19236 60620 19964 60676
rect 20020 60620 20030 60676
rect 20402 60620 20412 60676
rect 20468 60620 21308 60676
rect 21364 60620 21374 60676
rect 23314 60620 23324 60676
rect 23380 60620 24444 60676
rect 24500 60620 24510 60676
rect 27794 60620 27804 60676
rect 27860 60620 28924 60676
rect 28980 60620 29260 60676
rect 29316 60620 29326 60676
rect 31724 60620 31836 60676
rect 31892 60620 31902 60676
rect 32162 60620 32172 60676
rect 32228 60620 33852 60676
rect 33908 60620 33918 60676
rect 12114 60508 12124 60564
rect 12180 60508 16940 60564
rect 16996 60508 17006 60564
rect 18274 60508 18284 60564
rect 18340 60508 18732 60564
rect 18788 60508 18798 60564
rect 31602 60508 31612 60564
rect 31668 60508 32508 60564
rect 32564 60508 32956 60564
rect 33012 60508 33022 60564
rect 33366 60508 33404 60564
rect 33460 60508 33470 60564
rect 34972 60508 35308 60564
rect 35364 60508 35374 60564
rect 36306 60508 36316 60564
rect 36372 60508 37324 60564
rect 37380 60508 37390 60564
rect 40338 60508 40348 60564
rect 40404 60508 42028 60564
rect 42084 60508 42094 60564
rect 1586 60396 1596 60452
rect 1652 60396 3388 60452
rect 3444 60396 3454 60452
rect 7074 60396 7084 60452
rect 7140 60396 8092 60452
rect 8148 60396 10108 60452
rect 10164 60396 10668 60452
rect 10724 60396 11228 60452
rect 11284 60396 11294 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 33170 60284 33180 60340
rect 33236 60284 33740 60340
rect 33796 60284 33806 60340
rect 33740 60228 33796 60284
rect 34972 60228 35028 60508
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 38658 60284 38668 60340
rect 38724 60284 39788 60340
rect 39844 60284 40684 60340
rect 40740 60284 40750 60340
rect 33740 60172 35196 60228
rect 35252 60172 35262 60228
rect 19254 60060 19292 60116
rect 19348 60060 19358 60116
rect 22082 60060 22092 60116
rect 22148 60060 22764 60116
rect 22820 60060 22830 60116
rect 39106 60060 39116 60116
rect 39172 60060 39564 60116
rect 39620 60060 40460 60116
rect 40516 60060 40526 60116
rect 12674 59948 12684 60004
rect 12740 59948 15820 60004
rect 15876 59948 15886 60004
rect 18946 59948 18956 60004
rect 19012 59948 19852 60004
rect 19908 59948 19918 60004
rect 20290 59948 20300 60004
rect 20356 59948 21644 60004
rect 21700 59948 21710 60004
rect 24882 59948 24892 60004
rect 24948 59948 26460 60004
rect 26516 59948 26526 60004
rect 34850 59948 34860 60004
rect 34916 59948 37884 60004
rect 37940 59948 37950 60004
rect 34860 59892 34916 59948
rect 20514 59836 20524 59892
rect 20580 59836 22316 59892
rect 22372 59836 22382 59892
rect 22754 59836 22764 59892
rect 22820 59836 23324 59892
rect 23380 59836 23390 59892
rect 31714 59836 31724 59892
rect 31780 59836 32172 59892
rect 32228 59836 34916 59892
rect 37090 59836 37100 59892
rect 37156 59836 37660 59892
rect 37716 59836 37726 59892
rect 17378 59724 17388 59780
rect 17444 59724 18060 59780
rect 18116 59724 18126 59780
rect 31266 59724 31276 59780
rect 31332 59724 31612 59780
rect 31668 59724 31678 59780
rect 32386 59724 32396 59780
rect 32452 59724 33180 59780
rect 33236 59724 34076 59780
rect 34132 59724 34142 59780
rect 13346 59612 13356 59668
rect 13412 59612 17500 59668
rect 17556 59612 17566 59668
rect 31350 59612 31388 59668
rect 31444 59612 31454 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 25554 59500 25564 59556
rect 25620 59500 34972 59556
rect 35028 59500 35980 59556
rect 36036 59500 36046 59556
rect 7410 59388 7420 59444
rect 7476 59388 8652 59444
rect 8708 59388 8718 59444
rect 21858 59388 21868 59444
rect 21924 59388 41916 59444
rect 41972 59388 41982 59444
rect 16482 59276 16492 59332
rect 16548 59276 18060 59332
rect 18116 59276 18126 59332
rect 31266 59276 31276 59332
rect 31332 59276 32620 59332
rect 32676 59276 32686 59332
rect 43250 59276 43260 59332
rect 43316 59276 45836 59332
rect 45892 59276 45902 59332
rect 7970 59164 7980 59220
rect 8036 59164 9548 59220
rect 9604 59164 9614 59220
rect 18162 59164 18172 59220
rect 18228 59164 19628 59220
rect 19684 59164 19694 59220
rect 35634 59164 35644 59220
rect 35700 59164 36428 59220
rect 36484 59164 36876 59220
rect 36932 59164 36942 59220
rect 37202 59164 37212 59220
rect 37268 59164 38108 59220
rect 38164 59164 38174 59220
rect 6178 59052 6188 59108
rect 6244 59052 6412 59108
rect 6468 59052 6860 59108
rect 6916 59052 9996 59108
rect 10052 59052 10062 59108
rect 15474 59052 15484 59108
rect 15540 59052 17724 59108
rect 17780 59052 20636 59108
rect 20692 59052 20702 59108
rect 26114 59052 26124 59108
rect 26180 59052 27804 59108
rect 27860 59052 27870 59108
rect 31042 59052 31052 59108
rect 31108 59052 31724 59108
rect 31780 59052 31790 59108
rect 32162 59052 32172 59108
rect 32228 59052 32956 59108
rect 33012 59052 33516 59108
rect 33572 59052 33964 59108
rect 34020 59052 34030 59108
rect 34178 59052 34188 59108
rect 34244 59052 35980 59108
rect 36036 59052 36764 59108
rect 36820 59052 36830 59108
rect 38546 59052 38556 59108
rect 38612 59052 39004 59108
rect 39060 59052 39900 59108
rect 39956 59052 39966 59108
rect 6514 58940 6524 58996
rect 6580 58940 7868 58996
rect 7924 58940 7934 58996
rect 10658 58940 10668 58996
rect 10724 58940 11564 58996
rect 11620 58940 23548 58996
rect 23604 58940 24220 58996
rect 24276 58940 24286 58996
rect 36306 58940 36316 58996
rect 36372 58940 36988 58996
rect 37044 58940 38668 58996
rect 38724 58940 38734 58996
rect 4946 58828 4956 58884
rect 5012 58828 8484 58884
rect 8642 58828 8652 58884
rect 8708 58828 23100 58884
rect 23156 58828 23996 58884
rect 24052 58828 24062 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 8428 58772 8484 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 8428 58716 10668 58772
rect 10724 58716 10734 58772
rect 18386 58716 18396 58772
rect 18452 58716 18956 58772
rect 19012 58716 19022 58772
rect 9436 58660 9492 58716
rect 8754 58604 8764 58660
rect 8820 58604 9212 58660
rect 9268 58604 9278 58660
rect 9426 58604 9436 58660
rect 9492 58604 9502 58660
rect 26338 58604 26348 58660
rect 26404 58604 26908 58660
rect 26964 58604 26974 58660
rect 5954 58492 5964 58548
rect 6020 58492 6300 58548
rect 6356 58492 6748 58548
rect 6804 58492 6814 58548
rect 16370 58492 16380 58548
rect 16436 58492 16716 58548
rect 16772 58492 16782 58548
rect 25554 58492 25564 58548
rect 25620 58492 25900 58548
rect 25956 58492 28140 58548
rect 28196 58492 28206 58548
rect 5170 58380 5180 58436
rect 5236 58380 6636 58436
rect 6692 58380 7420 58436
rect 7476 58380 7486 58436
rect 12226 58380 12236 58436
rect 12292 58380 18060 58436
rect 18116 58380 18620 58436
rect 18676 58380 18686 58436
rect 25666 58380 25676 58436
rect 25732 58380 27020 58436
rect 27076 58380 27086 58436
rect 0 58324 800 58352
rect 49200 58324 50000 58352
rect 0 58268 1708 58324
rect 1764 58268 2492 58324
rect 2548 58268 2558 58324
rect 8306 58268 8316 58324
rect 8372 58268 11564 58324
rect 11620 58268 23100 58324
rect 23156 58268 23166 58324
rect 24434 58268 24444 58324
rect 24500 58268 25788 58324
rect 25844 58268 25854 58324
rect 40114 58268 40124 58324
rect 40180 58268 41132 58324
rect 41188 58268 41198 58324
rect 48066 58268 48076 58324
rect 48132 58268 50000 58324
rect 0 58240 800 58268
rect 49200 58240 50000 58268
rect 4610 58156 4620 58212
rect 4676 58156 5740 58212
rect 5796 58156 5806 58212
rect 9986 58156 9996 58212
rect 10052 58156 10556 58212
rect 10612 58156 10622 58212
rect 12338 58156 12348 58212
rect 12404 58156 13804 58212
rect 13860 58156 13870 58212
rect 20514 58156 20524 58212
rect 20580 58156 23884 58212
rect 23940 58156 23950 58212
rect 24994 58156 25004 58212
rect 25060 58156 26348 58212
rect 26404 58156 26414 58212
rect 28578 58156 28588 58212
rect 28644 58156 29148 58212
rect 29204 58156 29596 58212
rect 29652 58156 29662 58212
rect 36978 58156 36988 58212
rect 37044 58156 37996 58212
rect 38052 58156 38062 58212
rect 39218 58156 39228 58212
rect 39284 58156 39564 58212
rect 39620 58156 40012 58212
rect 40068 58156 40572 58212
rect 40628 58156 40638 58212
rect 43362 58156 43372 58212
rect 43428 58156 44044 58212
rect 44100 58156 44110 58212
rect 7410 58044 7420 58100
rect 7476 58044 7868 58100
rect 7924 58044 7934 58100
rect 9538 58044 9548 58100
rect 9604 58044 11004 58100
rect 11060 58044 11070 58100
rect 25218 58044 25228 58100
rect 25284 58044 25564 58100
rect 25620 58044 25630 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 8418 57932 8428 57988
rect 8484 57932 10108 57988
rect 10164 57932 10668 57988
rect 10724 57932 10734 57988
rect 15222 57932 15260 57988
rect 15316 57932 15326 57988
rect 16930 57932 16940 57988
rect 16996 57932 17948 57988
rect 18004 57932 18014 57988
rect 7186 57820 7196 57876
rect 7252 57820 7644 57876
rect 7700 57820 7710 57876
rect 8082 57820 8092 57876
rect 8148 57820 9940 57876
rect 10658 57820 10668 57876
rect 10724 57820 22652 57876
rect 22708 57820 23884 57876
rect 23940 57820 23950 57876
rect 24434 57820 24444 57876
rect 24500 57820 26908 57876
rect 44482 57820 44492 57876
rect 44548 57820 45612 57876
rect 45668 57820 45678 57876
rect 9884 57764 9940 57820
rect 26852 57764 26908 57820
rect 5954 57708 5964 57764
rect 6020 57708 6524 57764
rect 6580 57708 8764 57764
rect 8820 57708 8830 57764
rect 9874 57708 9884 57764
rect 9940 57708 9950 57764
rect 11442 57708 11452 57764
rect 11508 57708 11676 57764
rect 11732 57708 11742 57764
rect 13794 57708 13804 57764
rect 13860 57708 17500 57764
rect 17556 57708 17566 57764
rect 26852 57708 46844 57764
rect 46900 57708 46910 57764
rect 10742 57596 10780 57652
rect 10836 57596 10846 57652
rect 12562 57596 12572 57652
rect 12628 57596 14700 57652
rect 14756 57596 14766 57652
rect 15250 57596 15260 57652
rect 15316 57596 15484 57652
rect 15540 57596 15550 57652
rect 15698 57596 15708 57652
rect 15764 57596 15802 57652
rect 16818 57596 16828 57652
rect 16884 57596 17612 57652
rect 17668 57596 17678 57652
rect 17826 57596 17836 57652
rect 17892 57596 17902 57652
rect 19954 57596 19964 57652
rect 20020 57596 22204 57652
rect 22260 57596 22270 57652
rect 28354 57596 28364 57652
rect 28420 57596 28700 57652
rect 28756 57596 28766 57652
rect 33506 57596 33516 57652
rect 33572 57596 34076 57652
rect 34132 57596 39228 57652
rect 39284 57596 39676 57652
rect 39732 57596 39742 57652
rect 44566 57596 44604 57652
rect 44660 57596 44670 57652
rect 17836 57540 17892 57596
rect 7074 57484 7084 57540
rect 7140 57484 8764 57540
rect 8820 57484 8830 57540
rect 10098 57484 10108 57540
rect 10164 57484 10444 57540
rect 10500 57484 15148 57540
rect 15204 57484 15820 57540
rect 15876 57484 15886 57540
rect 16828 57484 17892 57540
rect 28914 57484 28924 57540
rect 28980 57484 38668 57540
rect 44258 57484 44268 57540
rect 44324 57484 45500 57540
rect 45556 57484 45566 57540
rect 16828 57428 16884 57484
rect 38612 57428 38668 57484
rect 6066 57372 6076 57428
rect 6132 57372 8540 57428
rect 8596 57372 8606 57428
rect 16818 57372 16828 57428
rect 16884 57372 16894 57428
rect 18722 57372 18732 57428
rect 18788 57372 18956 57428
rect 19012 57372 19404 57428
rect 19460 57372 19470 57428
rect 26898 57372 26908 57428
rect 26964 57372 28140 57428
rect 28196 57372 37324 57428
rect 37380 57372 38332 57428
rect 38388 57372 38398 57428
rect 38612 57372 44604 57428
rect 44660 57372 44670 57428
rect 30482 57260 30492 57316
rect 30548 57260 31052 57316
rect 31108 57260 31118 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 8950 57148 8988 57204
rect 9044 57148 9054 57204
rect 15250 57148 15260 57204
rect 15316 57148 16716 57204
rect 16772 57148 16782 57204
rect 20178 57148 20188 57204
rect 20244 57148 21420 57204
rect 21476 57148 21486 57204
rect 30258 57148 30268 57204
rect 30324 57148 30716 57204
rect 30772 57148 30782 57204
rect 45154 57148 45164 57204
rect 45220 57148 46060 57204
rect 46116 57148 46126 57204
rect 2034 57036 2044 57092
rect 2100 57036 2828 57092
rect 2884 57036 2894 57092
rect 14578 57036 14588 57092
rect 14644 57036 15708 57092
rect 15764 57036 15774 57092
rect 15922 57036 15932 57092
rect 15988 57036 16026 57092
rect 19842 57036 19852 57092
rect 19908 57036 21756 57092
rect 21812 57036 22428 57092
rect 22484 57036 22494 57092
rect 24210 57036 24220 57092
rect 24276 57036 27916 57092
rect 27972 57036 30156 57092
rect 30212 57036 31276 57092
rect 31332 57036 31342 57092
rect 41906 57036 41916 57092
rect 41972 57036 45500 57092
rect 45556 57036 45566 57092
rect 1362 56924 1372 56980
rect 1428 56924 5740 56980
rect 5796 56924 5806 56980
rect 12124 56924 18508 56980
rect 18564 56924 18574 56980
rect 23090 56924 23100 56980
rect 23156 56924 24108 56980
rect 24164 56924 25228 56980
rect 25284 56924 25294 56980
rect 44594 56924 44604 56980
rect 44660 56924 45052 56980
rect 45108 56924 45118 56980
rect 7074 56812 7084 56868
rect 7140 56812 7644 56868
rect 7700 56812 7710 56868
rect 8082 56812 8092 56868
rect 8148 56812 8988 56868
rect 9044 56812 9054 56868
rect 9874 56812 9884 56868
rect 9940 56812 10332 56868
rect 10388 56812 10398 56868
rect 12124 56756 12180 56924
rect 25666 56812 25676 56868
rect 25732 56812 26460 56868
rect 26516 56812 28252 56868
rect 28308 56812 29260 56868
rect 29316 56812 29326 56868
rect 40758 56812 40796 56868
rect 40852 56812 40862 56868
rect 43138 56812 43148 56868
rect 43204 56812 43708 56868
rect 43764 56812 43774 56868
rect 12114 56700 12124 56756
rect 12180 56700 12190 56756
rect 12338 56700 12348 56756
rect 12404 56700 13356 56756
rect 13412 56700 13422 56756
rect 15698 56700 15708 56756
rect 15764 56700 16492 56756
rect 16548 56700 16558 56756
rect 43026 56700 43036 56756
rect 43092 56700 43652 56756
rect 43596 56644 43652 56700
rect 11106 56588 11116 56644
rect 11172 56588 11564 56644
rect 11620 56588 12684 56644
rect 12740 56588 12750 56644
rect 26114 56588 26124 56644
rect 26180 56588 26460 56644
rect 26516 56588 26526 56644
rect 27570 56588 27580 56644
rect 27636 56588 29708 56644
rect 29764 56588 31612 56644
rect 31668 56588 31678 56644
rect 35746 56588 35756 56644
rect 35812 56588 37100 56644
rect 37156 56588 37166 56644
rect 43586 56588 43596 56644
rect 43652 56588 43662 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 14914 56364 14924 56420
rect 14980 56364 16940 56420
rect 16996 56364 18956 56420
rect 19012 56364 19022 56420
rect 23202 56364 23212 56420
rect 23268 56364 23324 56420
rect 23380 56364 25340 56420
rect 25396 56364 25406 56420
rect 26114 56364 26124 56420
rect 26180 56364 29036 56420
rect 29092 56364 29102 56420
rect 24434 56252 24444 56308
rect 24500 56252 24510 56308
rect 28438 56252 28476 56308
rect 28532 56252 28542 56308
rect 35634 56252 35644 56308
rect 35700 56252 37100 56308
rect 37156 56252 37166 56308
rect 5730 56140 5740 56196
rect 5796 56140 11564 56196
rect 11620 56140 12124 56196
rect 12180 56140 12190 56196
rect 13458 56140 13468 56196
rect 13524 56140 13916 56196
rect 13972 56140 13982 56196
rect 17154 56140 17164 56196
rect 17220 56140 17500 56196
rect 17556 56140 17566 56196
rect 18162 56140 18172 56196
rect 18228 56140 20636 56196
rect 20692 56140 20702 56196
rect 24444 56084 24500 56252
rect 30706 56140 30716 56196
rect 30772 56140 31500 56196
rect 31556 56140 31566 56196
rect 36642 56140 36652 56196
rect 36708 56140 37212 56196
rect 37268 56140 37278 56196
rect 38882 56140 38892 56196
rect 38948 56140 39788 56196
rect 39844 56140 40124 56196
rect 40180 56140 41020 56196
rect 41076 56140 42028 56196
rect 42084 56140 42094 56196
rect 13766 56028 13804 56084
rect 13860 56028 13870 56084
rect 24444 56028 31612 56084
rect 31668 56028 31678 56084
rect 13346 55916 13356 55972
rect 13412 55916 13916 55972
rect 13972 55916 13982 55972
rect 22418 55916 22428 55972
rect 22484 55916 26124 55972
rect 26180 55916 26190 55972
rect 30594 55916 30604 55972
rect 30660 55916 32844 55972
rect 32900 55916 32910 55972
rect 40898 55916 40908 55972
rect 40964 55916 41020 55972
rect 41076 55916 41580 55972
rect 41636 55916 41646 55972
rect 44566 55916 44604 55972
rect 44660 55916 44670 55972
rect 46722 55916 46732 55972
rect 46788 55916 47068 55972
rect 47124 55916 47134 55972
rect 0 55860 800 55888
rect 49200 55860 50000 55888
rect 0 55804 1708 55860
rect 1764 55804 2492 55860
rect 2548 55804 2558 55860
rect 7858 55804 7868 55860
rect 7924 55804 8204 55860
rect 8260 55804 9660 55860
rect 9716 55804 9726 55860
rect 18386 55804 18396 55860
rect 18452 55804 18732 55860
rect 18788 55804 18798 55860
rect 19058 55804 19068 55860
rect 19124 55804 20188 55860
rect 20244 55804 20254 55860
rect 48066 55804 48076 55860
rect 48132 55804 50000 55860
rect 0 55776 800 55804
rect 49200 55776 50000 55804
rect 29698 55692 29708 55748
rect 29764 55692 30604 55748
rect 30660 55692 30670 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 9650 55580 9660 55636
rect 9716 55580 11004 55636
rect 11060 55580 11070 55636
rect 17154 55580 17164 55636
rect 17220 55580 17948 55636
rect 18004 55580 18014 55636
rect 19170 55580 19180 55636
rect 19236 55580 26908 55636
rect 26852 55524 26908 55580
rect 12114 55468 12124 55524
rect 12180 55468 13580 55524
rect 13636 55468 13646 55524
rect 26852 55468 42140 55524
rect 42196 55468 42206 55524
rect 20402 55356 20412 55412
rect 20468 55356 21532 55412
rect 21588 55356 24892 55412
rect 24948 55356 24958 55412
rect 25666 55356 25676 55412
rect 25732 55356 27580 55412
rect 27636 55356 28028 55412
rect 28084 55356 32172 55412
rect 32228 55356 32238 55412
rect 35522 55356 35532 55412
rect 35588 55356 46732 55412
rect 46788 55356 46798 55412
rect 16930 55244 16940 55300
rect 16996 55244 18396 55300
rect 18452 55244 18462 55300
rect 22278 55244 22316 55300
rect 22372 55244 22382 55300
rect 22978 55244 22988 55300
rect 23044 55244 24668 55300
rect 24724 55244 24734 55300
rect 25414 55244 25452 55300
rect 25508 55244 25518 55300
rect 32498 55244 32508 55300
rect 32564 55244 33516 55300
rect 33572 55244 34412 55300
rect 34468 55244 34636 55300
rect 34692 55244 34702 55300
rect 46162 55244 46172 55300
rect 46228 55244 47068 55300
rect 47124 55244 47134 55300
rect 10770 55132 10780 55188
rect 10836 55132 11900 55188
rect 11956 55132 11966 55188
rect 15922 55132 15932 55188
rect 15988 55132 17052 55188
rect 17108 55132 17118 55188
rect 20290 55132 20300 55188
rect 20356 55132 21420 55188
rect 21476 55132 22876 55188
rect 22932 55132 22942 55188
rect 25554 55132 25564 55188
rect 25620 55132 26124 55188
rect 26180 55132 26190 55188
rect 27234 55132 27244 55188
rect 27300 55132 27916 55188
rect 27972 55132 28476 55188
rect 28532 55132 28542 55188
rect 33282 55132 33292 55188
rect 33348 55132 34188 55188
rect 34244 55132 34254 55188
rect 43474 55132 43484 55188
rect 43540 55132 43932 55188
rect 43988 55132 43998 55188
rect 20066 55020 20076 55076
rect 20132 55020 21980 55076
rect 22036 55020 22046 55076
rect 22754 55020 22764 55076
rect 22820 55020 25340 55076
rect 25396 55020 25406 55076
rect 34066 55020 34076 55076
rect 34132 55020 35756 55076
rect 35812 55020 36204 55076
rect 36260 55020 36270 55076
rect 40674 55020 40684 55076
rect 40740 55020 43148 55076
rect 43204 55020 43214 55076
rect 44034 55020 44044 55076
rect 44100 55020 45276 55076
rect 45332 55020 45342 55076
rect 12898 54908 12908 54964
rect 12964 54908 13580 54964
rect 13636 54908 13646 54964
rect 33394 54908 33404 54964
rect 33460 54908 33516 54964
rect 33572 54908 33964 54964
rect 34020 54908 34030 54964
rect 13580 54740 13636 54908
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 14438 54796 14476 54852
rect 14532 54796 14542 54852
rect 33730 54796 33740 54852
rect 33796 54796 34188 54852
rect 34244 54796 34254 54852
rect 46050 54796 46060 54852
rect 46116 54796 46284 54852
rect 46340 54796 46732 54852
rect 46788 54796 46798 54852
rect 6066 54684 6076 54740
rect 6132 54684 8540 54740
rect 8596 54684 8606 54740
rect 13580 54684 17948 54740
rect 18004 54684 18014 54740
rect 22418 54684 22428 54740
rect 22484 54684 38668 54740
rect 41654 54684 41692 54740
rect 41748 54684 41758 54740
rect 38612 54628 38668 54684
rect 4834 54572 4844 54628
rect 4900 54572 6188 54628
rect 6244 54572 6254 54628
rect 13570 54572 13580 54628
rect 13636 54572 13804 54628
rect 13860 54572 13870 54628
rect 14242 54572 14252 54628
rect 14308 54572 15036 54628
rect 15092 54572 15102 54628
rect 15474 54572 15484 54628
rect 15540 54572 16156 54628
rect 16212 54572 16222 54628
rect 17266 54572 17276 54628
rect 17332 54572 17612 54628
rect 17668 54572 21196 54628
rect 21252 54572 21262 54628
rect 26114 54572 26124 54628
rect 26180 54572 27132 54628
rect 27188 54572 27198 54628
rect 38612 54572 42028 54628
rect 42084 54572 42094 54628
rect 43026 54572 43036 54628
rect 43092 54572 43596 54628
rect 43652 54572 43662 54628
rect 5170 54460 5180 54516
rect 5236 54460 5852 54516
rect 5908 54460 6524 54516
rect 6580 54460 8092 54516
rect 8148 54460 8158 54516
rect 25778 54460 25788 54516
rect 25844 54460 25854 54516
rect 26226 54460 26236 54516
rect 26292 54460 26572 54516
rect 26628 54460 26638 54516
rect 26786 54460 26796 54516
rect 26852 54460 26908 54516
rect 26964 54460 26974 54516
rect 27570 54460 27580 54516
rect 27636 54460 28140 54516
rect 28196 54460 28206 54516
rect 25788 54404 25844 54460
rect 1922 54348 1932 54404
rect 1988 54348 2492 54404
rect 2548 54348 3388 54404
rect 3444 54348 3454 54404
rect 8418 54348 8428 54404
rect 8484 54348 10220 54404
rect 10276 54348 10286 54404
rect 25788 54348 29260 54404
rect 29316 54348 29326 54404
rect 32050 54348 32060 54404
rect 32116 54348 40796 54404
rect 40852 54348 41020 54404
rect 41076 54348 41086 54404
rect 41682 54348 41692 54404
rect 41748 54348 43148 54404
rect 43204 54348 43820 54404
rect 43876 54348 43886 54404
rect 20178 54236 20188 54292
rect 20244 54236 20972 54292
rect 21028 54236 21038 54292
rect 26002 54236 26012 54292
rect 26068 54236 27580 54292
rect 27636 54236 27646 54292
rect 39190 54236 39228 54292
rect 39284 54236 39294 54292
rect 14130 54124 14140 54180
rect 14196 54124 14924 54180
rect 14980 54124 14990 54180
rect 24434 54124 24444 54180
rect 24500 54124 27244 54180
rect 27300 54124 27468 54180
rect 27524 54124 27534 54180
rect 38770 54124 38780 54180
rect 38836 54124 40012 54180
rect 40068 54124 40078 54180
rect 41206 54124 41244 54180
rect 41300 54124 41310 54180
rect 42130 54124 42140 54180
rect 42196 54124 46620 54180
rect 46676 54124 46686 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 11442 54012 11452 54068
rect 11508 54012 11900 54068
rect 11956 54012 11966 54068
rect 24770 54012 24780 54068
rect 24836 54012 26796 54068
rect 26852 54012 26862 54068
rect 28102 54012 28140 54068
rect 28196 54012 28206 54068
rect 37426 54012 37436 54068
rect 37492 54012 37884 54068
rect 37940 54012 38332 54068
rect 38388 54012 42924 54068
rect 42980 54012 43484 54068
rect 43540 54012 43550 54068
rect 6038 53900 6076 53956
rect 6132 53900 6142 53956
rect 19170 53900 19180 53956
rect 19236 53900 45164 53956
rect 45220 53900 45230 53956
rect 13122 53788 13132 53844
rect 13188 53788 22316 53844
rect 22372 53788 22382 53844
rect 27906 53788 27916 53844
rect 27972 53788 29148 53844
rect 29204 53788 29214 53844
rect 32946 53788 32956 53844
rect 33012 53788 33516 53844
rect 33572 53788 40684 53844
rect 40740 53788 41916 53844
rect 41972 53788 41982 53844
rect 44258 53788 44268 53844
rect 44324 53788 44940 53844
rect 44996 53788 45006 53844
rect 1810 53676 1820 53732
rect 1876 53676 3388 53732
rect 13234 53676 13244 53732
rect 13300 53676 14812 53732
rect 14868 53676 14878 53732
rect 20514 53676 20524 53732
rect 20580 53676 21532 53732
rect 21588 53676 21598 53732
rect 23986 53676 23996 53732
rect 24052 53676 25676 53732
rect 25732 53676 25742 53732
rect 27122 53676 27132 53732
rect 27188 53676 29932 53732
rect 29988 53676 29998 53732
rect 47058 53676 47068 53732
rect 47124 53676 47404 53732
rect 47460 53676 47470 53732
rect 3332 53508 3388 53676
rect 21532 53620 21588 53676
rect 5954 53564 5964 53620
rect 6020 53564 6636 53620
rect 6692 53564 6702 53620
rect 9762 53564 9772 53620
rect 9828 53564 10556 53620
rect 10612 53564 10622 53620
rect 10994 53564 11004 53620
rect 11060 53564 11564 53620
rect 11620 53564 14028 53620
rect 14084 53564 14700 53620
rect 14756 53564 14766 53620
rect 15810 53564 15820 53620
rect 15876 53564 16268 53620
rect 16324 53564 16334 53620
rect 21532 53564 22988 53620
rect 23044 53564 25452 53620
rect 25508 53564 26796 53620
rect 26852 53564 26862 53620
rect 27570 53564 27580 53620
rect 27636 53564 28252 53620
rect 28308 53564 28318 53620
rect 31602 53564 31612 53620
rect 31668 53564 38668 53620
rect 41122 53564 41132 53620
rect 41188 53564 41468 53620
rect 41524 53564 41534 53620
rect 42130 53564 42140 53620
rect 42196 53564 45836 53620
rect 45892 53564 45902 53620
rect 48066 53564 48076 53620
rect 48132 53564 48142 53620
rect 38612 53508 38668 53564
rect 3332 53452 5068 53508
rect 5124 53452 5516 53508
rect 5572 53452 5582 53508
rect 16370 53452 16380 53508
rect 16436 53452 17724 53508
rect 17780 53452 18620 53508
rect 18676 53452 18686 53508
rect 25330 53452 25340 53508
rect 25396 53452 25406 53508
rect 26226 53452 26236 53508
rect 26292 53452 28140 53508
rect 28196 53452 28206 53508
rect 31826 53452 31836 53508
rect 31892 53452 33404 53508
rect 33460 53452 33470 53508
rect 38612 53452 46956 53508
rect 47012 53452 47022 53508
rect 0 53312 800 53424
rect 25340 53396 25396 53452
rect 48076 53396 48132 53564
rect 49200 53396 50000 53424
rect 20738 53340 20748 53396
rect 20804 53340 20814 53396
rect 25340 53340 35532 53396
rect 35588 53340 35598 53396
rect 41122 53340 41132 53396
rect 41188 53340 41916 53396
rect 41972 53340 42364 53396
rect 42420 53340 42430 53396
rect 48076 53340 50000 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 4162 53116 4172 53172
rect 4228 53116 7532 53172
rect 7588 53116 8876 53172
rect 8932 53116 8942 53172
rect 13570 53116 13580 53172
rect 13636 53116 20524 53172
rect 20580 53116 20590 53172
rect 3332 53004 10780 53060
rect 10836 53004 11228 53060
rect 11284 53004 11294 53060
rect 13794 53004 13804 53060
rect 13860 53004 13870 53060
rect 3332 52948 3388 53004
rect 13804 52948 13860 53004
rect 20748 52948 20804 53340
rect 49200 53312 50000 53340
rect 27458 53228 27468 53284
rect 27524 53228 27916 53284
rect 27972 53228 27982 53284
rect 31378 53228 31388 53284
rect 31444 53228 41020 53284
rect 41076 53228 42028 53284
rect 42084 53228 42094 53284
rect 23202 53004 23212 53060
rect 23268 53004 24556 53060
rect 24612 53004 24622 53060
rect 33394 53004 33404 53060
rect 33460 53004 33740 53060
rect 33796 53004 33806 53060
rect 40226 53004 40236 53060
rect 40292 53004 41244 53060
rect 41300 53004 41310 53060
rect 1698 52892 1708 52948
rect 1764 52892 3388 52948
rect 9874 52892 9884 52948
rect 9940 52892 10332 52948
rect 10388 52892 10398 52948
rect 10630 52892 10668 52948
rect 10724 52892 10734 52948
rect 13804 52892 14140 52948
rect 14196 52892 14206 52948
rect 14466 52892 14476 52948
rect 14532 52892 15260 52948
rect 15316 52892 15326 52948
rect 15698 52892 15708 52948
rect 15764 52892 16604 52948
rect 16660 52892 16670 52948
rect 18498 52892 18508 52948
rect 18564 52892 19852 52948
rect 19908 52892 19918 52948
rect 20738 52892 20748 52948
rect 20804 52892 20814 52948
rect 21970 52892 21980 52948
rect 22036 52892 22652 52948
rect 22708 52892 22718 52948
rect 35634 52892 35644 52948
rect 35700 52892 36316 52948
rect 36372 52892 37436 52948
rect 37492 52892 37502 52948
rect 40870 52892 40908 52948
rect 40964 52892 40974 52948
rect 2258 52780 2268 52836
rect 2324 52780 9548 52836
rect 9604 52780 9614 52836
rect 12898 52780 12908 52836
rect 12964 52780 19180 52836
rect 19236 52780 19246 52836
rect 21858 52780 21868 52836
rect 21924 52780 25900 52836
rect 25956 52780 25966 52836
rect 29474 52780 29484 52836
rect 29540 52780 30156 52836
rect 30212 52780 30716 52836
rect 30772 52780 30782 52836
rect 31378 52780 31388 52836
rect 31444 52780 32172 52836
rect 32228 52780 39116 52836
rect 39172 52780 41244 52836
rect 41300 52780 41310 52836
rect 6290 52668 6300 52724
rect 6356 52668 6748 52724
rect 6804 52668 8428 52724
rect 8484 52668 10556 52724
rect 10612 52668 10622 52724
rect 15222 52668 15260 52724
rect 15316 52668 15326 52724
rect 22866 52668 22876 52724
rect 22932 52668 23548 52724
rect 23604 52668 24444 52724
rect 24500 52668 24510 52724
rect 26226 52668 26236 52724
rect 26292 52668 28700 52724
rect 28756 52668 28766 52724
rect 33618 52668 33628 52724
rect 33684 52668 34300 52724
rect 34356 52668 39564 52724
rect 39620 52668 41804 52724
rect 41860 52668 41870 52724
rect 8866 52556 8876 52612
rect 8932 52556 16604 52612
rect 16660 52556 20300 52612
rect 20356 52556 20366 52612
rect 23202 52556 23212 52612
rect 23268 52556 24108 52612
rect 24164 52556 24174 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 5842 52444 5852 52500
rect 5908 52444 6244 52500
rect 8082 52444 8092 52500
rect 8148 52444 8764 52500
rect 8820 52444 10780 52500
rect 10836 52444 18396 52500
rect 18452 52444 18462 52500
rect 22530 52444 22540 52500
rect 22596 52444 22988 52500
rect 23044 52444 23054 52500
rect 6188 52388 6244 52444
rect 4722 52332 4732 52388
rect 4788 52332 5964 52388
rect 6020 52332 6030 52388
rect 6178 52332 6188 52388
rect 6244 52332 23436 52388
rect 23492 52332 23502 52388
rect 30258 52332 30268 52388
rect 30324 52332 41132 52388
rect 41188 52332 41198 52388
rect 41654 52332 41692 52388
rect 41748 52332 41758 52388
rect 4834 52220 4844 52276
rect 4900 52220 4910 52276
rect 16118 52220 16156 52276
rect 16212 52220 16222 52276
rect 28466 52220 28476 52276
rect 28532 52220 32284 52276
rect 32340 52220 33404 52276
rect 33460 52220 33470 52276
rect 37202 52220 37212 52276
rect 37268 52220 37996 52276
rect 38052 52220 38062 52276
rect 41010 52220 41020 52276
rect 41076 52220 41244 52276
rect 41300 52220 41916 52276
rect 41972 52220 41982 52276
rect 4844 52164 4900 52220
rect 4162 52108 4172 52164
rect 4228 52108 5628 52164
rect 5684 52108 5694 52164
rect 12562 52108 12572 52164
rect 12628 52108 13356 52164
rect 13412 52108 13422 52164
rect 13570 52108 13580 52164
rect 13636 52108 13916 52164
rect 13972 52108 13982 52164
rect 19058 52108 19068 52164
rect 19124 52108 19852 52164
rect 19908 52108 19918 52164
rect 21420 52108 22316 52164
rect 22372 52108 22382 52164
rect 24658 52108 24668 52164
rect 24724 52108 26684 52164
rect 26740 52108 29260 52164
rect 29316 52108 29708 52164
rect 29764 52108 29774 52164
rect 31714 52108 31724 52164
rect 31780 52108 32172 52164
rect 32228 52108 32238 52164
rect 41020 52108 41804 52164
rect 41860 52108 41870 52164
rect 21420 52052 21476 52108
rect 3602 51996 3612 52052
rect 3668 51996 4956 52052
rect 5012 51996 6300 52052
rect 6356 51996 6366 52052
rect 6738 51996 6748 52052
rect 6804 51996 8316 52052
rect 8372 51996 8382 52052
rect 15362 51996 15372 52052
rect 15428 51996 15708 52052
rect 15764 51996 15774 52052
rect 18834 51996 18844 52052
rect 18900 51996 21420 52052
rect 21476 51996 21486 52052
rect 24434 51996 24444 52052
rect 24500 51996 25340 52052
rect 25396 51996 25406 52052
rect 31602 51996 31612 52052
rect 31668 51996 32620 52052
rect 32676 51996 32686 52052
rect 41020 51940 41076 52108
rect 3826 51884 3836 51940
rect 3892 51884 8652 51940
rect 8708 51884 8718 51940
rect 11778 51884 11788 51940
rect 11844 51884 12348 51940
rect 12404 51884 12414 51940
rect 19394 51884 19404 51940
rect 19460 51884 21196 51940
rect 21252 51884 22764 51940
rect 22820 51884 25004 51940
rect 25060 51884 25070 51940
rect 25778 51884 25788 51940
rect 25844 51884 26236 51940
rect 26292 51884 26302 51940
rect 32722 51884 32732 51940
rect 32788 51884 34972 51940
rect 35028 51884 35532 51940
rect 35588 51884 35598 51940
rect 41010 51884 41020 51940
rect 41076 51884 41086 51940
rect 18946 51772 18956 51828
rect 19012 51772 19516 51828
rect 19572 51772 19582 51828
rect 22306 51772 22316 51828
rect 22372 51772 22876 51828
rect 22932 51772 22942 51828
rect 26786 51772 26796 51828
rect 26852 51772 38668 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 8642 51660 8652 51716
rect 8708 51660 9660 51716
rect 9716 51660 9726 51716
rect 17826 51660 17836 51716
rect 17892 51660 18732 51716
rect 18788 51660 18798 51716
rect 27010 51660 27020 51716
rect 27076 51660 29036 51716
rect 29092 51660 29372 51716
rect 29428 51660 29438 51716
rect 8530 51548 8540 51604
rect 8596 51548 9772 51604
rect 9828 51548 9838 51604
rect 22530 51548 22540 51604
rect 22596 51548 23884 51604
rect 23940 51548 23950 51604
rect 24210 51548 24220 51604
rect 24276 51548 25452 51604
rect 25508 51548 25518 51604
rect 27356 51548 29820 51604
rect 29876 51548 29886 51604
rect 2706 51436 2716 51492
rect 2772 51436 4172 51492
rect 4228 51436 4238 51492
rect 20514 51436 20524 51492
rect 20580 51436 27132 51492
rect 27188 51436 27198 51492
rect 4834 51324 4844 51380
rect 4900 51324 5628 51380
rect 5684 51324 6524 51380
rect 6580 51324 6590 51380
rect 7634 51324 7644 51380
rect 7700 51324 8764 51380
rect 8820 51324 8830 51380
rect 22754 51324 22764 51380
rect 22820 51324 23324 51380
rect 23380 51324 23390 51380
rect 24882 51324 24892 51380
rect 24948 51324 26908 51380
rect 26852 51268 26908 51324
rect 27356 51268 27412 51548
rect 28802 51436 28812 51492
rect 28868 51436 38164 51492
rect 32498 51324 32508 51380
rect 32564 51324 32844 51380
rect 32900 51324 32910 51380
rect 34402 51324 34412 51380
rect 34468 51324 35420 51380
rect 35476 51324 35486 51380
rect 10322 51212 10332 51268
rect 10388 51212 10556 51268
rect 10612 51212 23436 51268
rect 23492 51212 23502 51268
rect 26852 51212 27412 51268
rect 28466 51212 28476 51268
rect 28532 51212 30268 51268
rect 30324 51212 30334 51268
rect 35746 51212 35756 51268
rect 35812 51212 36316 51268
rect 36372 51212 36382 51268
rect 38108 51156 38164 51436
rect 38612 51268 38668 51772
rect 40786 51660 40796 51716
rect 40852 51660 41132 51716
rect 41188 51660 41198 51716
rect 38882 51548 38892 51604
rect 38948 51548 40012 51604
rect 40068 51548 40078 51604
rect 42690 51436 42700 51492
rect 42756 51436 43820 51492
rect 43876 51436 43886 51492
rect 42018 51324 42028 51380
rect 42084 51324 42588 51380
rect 42644 51324 44044 51380
rect 44100 51324 44110 51380
rect 46274 51324 46284 51380
rect 46340 51324 46844 51380
rect 46900 51324 46910 51380
rect 38612 51212 43820 51268
rect 43876 51212 43886 51268
rect 28774 51100 28812 51156
rect 28868 51100 28878 51156
rect 31490 51100 31500 51156
rect 31556 51100 35588 51156
rect 38108 51100 38668 51156
rect 38724 51100 38734 51156
rect 40870 51100 40908 51156
rect 40964 51100 40974 51156
rect 35532 51044 35588 51100
rect 6178 50988 6188 51044
rect 6244 50988 7756 51044
rect 7812 50988 7822 51044
rect 12674 50988 12684 51044
rect 12740 50988 13916 51044
rect 13972 50988 13982 51044
rect 18722 50988 18732 51044
rect 18788 50988 18956 51044
rect 19012 50988 19022 51044
rect 35532 50988 42028 51044
rect 42084 50988 42094 51044
rect 0 50848 800 50960
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 49200 50932 50000 50960
rect 18610 50876 18620 50932
rect 18676 50876 20076 50932
rect 20132 50876 26796 50932
rect 26852 50876 26862 50932
rect 34514 50876 34524 50932
rect 34580 50876 34590 50932
rect 35532 50876 35756 50932
rect 35812 50876 35822 50932
rect 48066 50876 48076 50932
rect 48132 50876 50000 50932
rect 34524 50820 34580 50876
rect 35532 50820 35588 50876
rect 49200 50848 50000 50876
rect 26226 50764 26236 50820
rect 26292 50764 28252 50820
rect 28308 50764 28318 50820
rect 28476 50764 30324 50820
rect 34524 50764 35588 50820
rect 35644 50764 40348 50820
rect 40404 50764 41580 50820
rect 41636 50764 41646 50820
rect 28476 50708 28532 50764
rect 3714 50652 3724 50708
rect 3780 50652 5628 50708
rect 5684 50652 6860 50708
rect 6916 50652 6926 50708
rect 15362 50652 15372 50708
rect 15428 50652 17052 50708
rect 17108 50652 17118 50708
rect 21186 50652 21196 50708
rect 21252 50652 21262 50708
rect 26674 50652 26684 50708
rect 26740 50652 28140 50708
rect 28196 50652 28532 50708
rect 29596 50652 29820 50708
rect 29876 50652 29886 50708
rect 2482 50540 2492 50596
rect 2548 50540 3164 50596
rect 3220 50540 3230 50596
rect 4498 50540 4508 50596
rect 4564 50540 6076 50596
rect 6132 50540 6142 50596
rect 8306 50540 8316 50596
rect 8372 50540 9772 50596
rect 9828 50540 9838 50596
rect 18498 50540 18508 50596
rect 18564 50540 19068 50596
rect 19124 50540 19404 50596
rect 19460 50540 19470 50596
rect 21196 50484 21252 50652
rect 21410 50540 21420 50596
rect 21476 50540 22204 50596
rect 22260 50540 22270 50596
rect 27458 50540 27468 50596
rect 27524 50540 28364 50596
rect 28420 50540 28430 50596
rect 2818 50428 2828 50484
rect 2884 50428 3836 50484
rect 3892 50428 3902 50484
rect 4050 50428 4060 50484
rect 4116 50428 7644 50484
rect 7700 50428 7710 50484
rect 8418 50428 8428 50484
rect 8484 50428 8876 50484
rect 8932 50428 10220 50484
rect 10276 50428 10286 50484
rect 21196 50428 21364 50484
rect 25890 50428 25900 50484
rect 25956 50428 27020 50484
rect 27076 50428 27086 50484
rect 28018 50428 28028 50484
rect 28084 50428 29036 50484
rect 29092 50428 29102 50484
rect 21308 50372 21364 50428
rect 29596 50372 29652 50652
rect 30268 50596 30324 50764
rect 33282 50652 33292 50708
rect 33348 50652 33964 50708
rect 34020 50652 34524 50708
rect 34580 50652 34590 50708
rect 35644 50596 35700 50764
rect 36306 50652 36316 50708
rect 36372 50652 39452 50708
rect 39508 50652 39518 50708
rect 43026 50652 43036 50708
rect 43092 50652 43484 50708
rect 43540 50652 43550 50708
rect 30258 50540 30268 50596
rect 30324 50540 35700 50596
rect 37650 50540 37660 50596
rect 37716 50540 38332 50596
rect 38388 50540 38398 50596
rect 38098 50428 38108 50484
rect 38164 50428 38892 50484
rect 38948 50428 38958 50484
rect 44258 50428 44268 50484
rect 44324 50428 44334 50484
rect 10322 50316 10332 50372
rect 10388 50316 10668 50372
rect 10724 50316 10734 50372
rect 12226 50316 12236 50372
rect 12292 50316 12684 50372
rect 12740 50316 20636 50372
rect 20692 50316 20702 50372
rect 20962 50316 20972 50372
rect 21028 50316 21364 50372
rect 28578 50316 28588 50372
rect 28644 50316 28924 50372
rect 28980 50316 28990 50372
rect 29250 50316 29260 50372
rect 29316 50316 29652 50372
rect 31042 50316 31052 50372
rect 31108 50316 31724 50372
rect 31780 50316 31790 50372
rect 33170 50316 33180 50372
rect 33236 50316 33246 50372
rect 33394 50316 33404 50372
rect 33460 50316 34188 50372
rect 34244 50316 34254 50372
rect 33180 50260 33236 50316
rect 1922 50204 1932 50260
rect 1988 50204 2380 50260
rect 2436 50204 3276 50260
rect 3332 50204 8764 50260
rect 8820 50204 8830 50260
rect 10434 50204 10444 50260
rect 10500 50204 10780 50260
rect 10836 50204 10846 50260
rect 11330 50204 11340 50260
rect 11396 50204 11406 50260
rect 25778 50204 25788 50260
rect 25844 50204 28252 50260
rect 28308 50204 28318 50260
rect 30370 50204 30380 50260
rect 30436 50204 33236 50260
rect 44268 50260 44324 50428
rect 44268 50204 45612 50260
rect 45668 50204 45678 50260
rect 11340 50148 11396 50204
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 2034 50092 2044 50148
rect 2100 50092 2492 50148
rect 2548 50092 2558 50148
rect 11340 50092 11564 50148
rect 11620 50092 11630 50148
rect 15922 50092 15932 50148
rect 15988 50092 16380 50148
rect 16436 50092 16446 50148
rect 11414 49980 11452 50036
rect 11508 49980 11518 50036
rect 11732 49980 17612 50036
rect 17668 49980 17678 50036
rect 17910 49980 17948 50036
rect 18004 49980 18014 50036
rect 18834 49980 18844 50036
rect 18900 49980 20412 50036
rect 20468 49980 21644 50036
rect 21700 49980 21710 50036
rect 23492 49980 25340 50036
rect 25396 49980 25452 50036
rect 25508 49980 25518 50036
rect 40898 49980 40908 50036
rect 40964 49980 41580 50036
rect 41636 49980 41646 50036
rect 11732 49924 11788 49980
rect 10994 49868 11004 49924
rect 11060 49868 11788 49924
rect 12338 49868 12348 49924
rect 12404 49868 13468 49924
rect 13524 49868 13534 49924
rect 21410 49868 21420 49924
rect 21476 49868 21868 49924
rect 21924 49868 22316 49924
rect 22372 49868 22382 49924
rect 2370 49756 2380 49812
rect 2436 49756 4060 49812
rect 4116 49756 4126 49812
rect 11106 49756 11116 49812
rect 11172 49756 12124 49812
rect 12180 49756 12190 49812
rect 13794 49756 13804 49812
rect 13860 49756 15596 49812
rect 15652 49756 19740 49812
rect 19796 49756 19806 49812
rect 23426 49756 23436 49812
rect 23492 49756 23548 49980
rect 26114 49868 26124 49924
rect 26180 49868 26572 49924
rect 26628 49868 28028 49924
rect 28084 49868 28094 49924
rect 33394 49868 33404 49924
rect 33460 49868 34300 49924
rect 34356 49868 34366 49924
rect 39554 49868 39564 49924
rect 39620 49868 41020 49924
rect 41076 49868 41086 49924
rect 46274 49868 46284 49924
rect 46340 49868 47740 49924
rect 47796 49868 47806 49924
rect 27122 49756 27132 49812
rect 27188 49756 28364 49812
rect 28420 49756 28430 49812
rect 32722 49756 32732 49812
rect 32788 49756 33068 49812
rect 33124 49756 33740 49812
rect 33796 49756 33806 49812
rect 46386 49756 46396 49812
rect 46452 49756 47516 49812
rect 47572 49756 47964 49812
rect 48020 49756 48030 49812
rect 1922 49644 1932 49700
rect 1988 49644 2940 49700
rect 2996 49644 5908 49700
rect 10546 49644 10556 49700
rect 10612 49644 10780 49700
rect 10836 49644 10846 49700
rect 15250 49644 15260 49700
rect 15316 49644 16156 49700
rect 16212 49644 16222 49700
rect 23986 49644 23996 49700
rect 24052 49644 24668 49700
rect 24724 49644 24734 49700
rect 25330 49644 25340 49700
rect 25396 49644 28588 49700
rect 28644 49644 28654 49700
rect 31490 49644 31500 49700
rect 31556 49644 33180 49700
rect 33236 49644 33246 49700
rect 5852 49588 5908 49644
rect 5842 49532 5852 49588
rect 5908 49532 5918 49588
rect 11106 49532 11116 49588
rect 11172 49532 12236 49588
rect 12292 49532 12302 49588
rect 15026 49532 15036 49588
rect 15092 49532 16268 49588
rect 16324 49532 16334 49588
rect 19058 49532 19068 49588
rect 19124 49532 20636 49588
rect 20692 49532 21756 49588
rect 21812 49532 21822 49588
rect 34850 49532 34860 49588
rect 34916 49532 35868 49588
rect 35924 49532 35934 49588
rect 41010 49532 41020 49588
rect 41076 49532 42812 49588
rect 42868 49532 43708 49588
rect 43764 49532 43774 49588
rect 5506 49420 5516 49476
rect 5572 49420 6636 49476
rect 6692 49420 23324 49476
rect 23380 49420 23660 49476
rect 23716 49420 23726 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 15586 49308 15596 49364
rect 15652 49308 15932 49364
rect 15988 49308 15998 49364
rect 17714 49308 17724 49364
rect 17780 49308 18620 49364
rect 18676 49308 18686 49364
rect 19618 49308 19628 49364
rect 19684 49308 20300 49364
rect 20356 49308 21196 49364
rect 21252 49308 21262 49364
rect 26002 49308 26012 49364
rect 26068 49308 27132 49364
rect 27188 49308 27198 49364
rect 18386 49196 18396 49252
rect 18452 49196 43260 49252
rect 43316 49196 43326 49252
rect 16034 49084 16044 49140
rect 16100 49084 22484 49140
rect 24658 49084 24668 49140
rect 24724 49084 26460 49140
rect 26516 49084 26740 49140
rect 27346 49084 27356 49140
rect 27412 49084 31388 49140
rect 31444 49084 31454 49140
rect 32050 49084 32060 49140
rect 32116 49084 39676 49140
rect 39732 49084 39742 49140
rect 22428 49028 22484 49084
rect 26684 49028 26740 49084
rect 8194 48972 8204 49028
rect 8260 48972 8988 49028
rect 9044 48972 9054 49028
rect 9202 48972 9212 49028
rect 9268 48972 15708 49028
rect 15764 48972 18620 49028
rect 18676 48972 18686 49028
rect 19394 48972 19404 49028
rect 19460 48972 20188 49028
rect 20244 48972 20254 49028
rect 20738 48972 20748 49028
rect 20804 48972 22204 49028
rect 22260 48972 22270 49028
rect 22428 48972 26012 49028
rect 26068 48972 26078 49028
rect 26674 48972 26684 49028
rect 26740 48972 26750 49028
rect 27010 48972 27020 49028
rect 27076 48972 27804 49028
rect 27860 48972 29148 49028
rect 29204 48972 29214 49028
rect 30156 48972 32620 49028
rect 32676 48972 32686 49028
rect 38612 48972 38668 49084
rect 38724 48972 38734 49028
rect 39554 48972 39564 49028
rect 39620 48972 40012 49028
rect 40068 48972 41132 49028
rect 41188 48972 41198 49028
rect 45490 48972 45500 49028
rect 45556 48972 46732 49028
rect 46788 48972 46956 49028
rect 47012 48972 47022 49028
rect 13794 48860 13804 48916
rect 13860 48860 14140 48916
rect 14196 48860 14206 48916
rect 16258 48860 16268 48916
rect 16324 48860 19516 48916
rect 19572 48860 19582 48916
rect 24322 48860 24332 48916
rect 24388 48860 29932 48916
rect 29988 48860 29998 48916
rect 30156 48804 30212 48972
rect 30594 48860 30604 48916
rect 30660 48860 31724 48916
rect 31780 48860 32396 48916
rect 32452 48860 32462 48916
rect 32946 48860 32956 48916
rect 33012 48860 33628 48916
rect 33684 48860 34972 48916
rect 35028 48860 35532 48916
rect 35588 48860 35598 48916
rect 40114 48860 40124 48916
rect 40180 48860 41580 48916
rect 41636 48860 41646 48916
rect 1586 48748 1596 48804
rect 1652 48748 11228 48804
rect 11284 48748 14252 48804
rect 14308 48748 14318 48804
rect 15250 48748 15260 48804
rect 15316 48748 15820 48804
rect 15876 48748 16156 48804
rect 16212 48748 16222 48804
rect 20178 48748 20188 48804
rect 20244 48748 21308 48804
rect 21364 48748 21374 48804
rect 27794 48748 27804 48804
rect 27860 48748 28028 48804
rect 28084 48748 30212 48804
rect 30706 48748 30716 48804
rect 30772 48748 32732 48804
rect 32788 48748 32798 48804
rect 33282 48748 33292 48804
rect 33348 48748 33404 48804
rect 33460 48748 34300 48804
rect 34356 48748 34366 48804
rect 34850 48748 34860 48804
rect 34916 48748 35308 48804
rect 35364 48748 36876 48804
rect 36932 48748 36942 48804
rect 39106 48748 39116 48804
rect 39172 48748 39228 48804
rect 39284 48748 39294 48804
rect 40002 48748 40012 48804
rect 40068 48748 40684 48804
rect 40740 48748 40750 48804
rect 47730 48748 47740 48804
rect 47796 48748 47806 48804
rect 33292 48692 33348 48748
rect 13794 48636 13804 48692
rect 13860 48636 14476 48692
rect 14532 48636 14542 48692
rect 31826 48636 31836 48692
rect 31892 48636 33348 48692
rect 35718 48636 35756 48692
rect 35812 48636 35822 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 30034 48524 30044 48580
rect 30100 48524 38668 48580
rect 41122 48524 41132 48580
rect 41188 48524 41580 48580
rect 41636 48524 41646 48580
rect 0 48384 800 48496
rect 38612 48468 38668 48524
rect 47740 48468 47796 48748
rect 49200 48468 50000 48496
rect 1698 48412 1708 48468
rect 1764 48412 3388 48468
rect 4386 48412 4396 48468
rect 4452 48412 4844 48468
rect 4900 48412 6076 48468
rect 6132 48412 6636 48468
rect 6692 48412 6702 48468
rect 7074 48412 7084 48468
rect 7140 48412 8540 48468
rect 8596 48412 8988 48468
rect 9044 48412 9548 48468
rect 9604 48412 9614 48468
rect 9874 48412 9884 48468
rect 9940 48412 13020 48468
rect 13076 48412 13086 48468
rect 38612 48412 39340 48468
rect 39396 48412 39406 48468
rect 43250 48412 43260 48468
rect 43316 48412 47180 48468
rect 47236 48412 47246 48468
rect 47740 48412 50000 48468
rect 3332 48356 3388 48412
rect 9884 48356 9940 48412
rect 47180 48356 47236 48412
rect 49200 48384 50000 48412
rect 3332 48300 3612 48356
rect 3668 48300 9940 48356
rect 12562 48300 12572 48356
rect 12628 48300 13580 48356
rect 13636 48300 17948 48356
rect 18004 48300 18014 48356
rect 20972 48300 33852 48356
rect 33908 48300 33918 48356
rect 36418 48300 36428 48356
rect 36484 48300 37212 48356
rect 37268 48300 37278 48356
rect 37874 48300 37884 48356
rect 37940 48300 38668 48356
rect 38724 48300 38734 48356
rect 39554 48300 39564 48356
rect 39620 48300 40460 48356
rect 40516 48300 41356 48356
rect 41412 48300 41422 48356
rect 43810 48300 43820 48356
rect 43876 48300 44492 48356
rect 44548 48300 44558 48356
rect 47180 48300 47740 48356
rect 47796 48300 47806 48356
rect 20972 48244 21028 48300
rect 2482 48188 2492 48244
rect 2548 48188 3500 48244
rect 3556 48188 4284 48244
rect 4340 48188 4350 48244
rect 7186 48188 7196 48244
rect 7252 48188 8204 48244
rect 8260 48188 8270 48244
rect 8950 48188 8988 48244
rect 9044 48188 9054 48244
rect 9212 48188 21028 48244
rect 23650 48188 23660 48244
rect 23716 48188 47292 48244
rect 47348 48188 47358 48244
rect 9212 48132 9268 48188
rect 1138 48076 1148 48132
rect 1204 48076 9268 48132
rect 13570 48076 13580 48132
rect 13636 48076 18620 48132
rect 18676 48076 23548 48132
rect 23604 48076 23614 48132
rect 24546 48076 24556 48132
rect 24612 48076 25788 48132
rect 25844 48076 25854 48132
rect 34402 48076 34412 48132
rect 34468 48076 34972 48132
rect 35028 48076 35038 48132
rect 35858 48076 35868 48132
rect 35924 48076 37100 48132
rect 37156 48076 37166 48132
rect 37986 48076 37996 48132
rect 38052 48076 38556 48132
rect 38612 48076 38622 48132
rect 40114 48076 40124 48132
rect 40180 48076 41020 48132
rect 41076 48076 41086 48132
rect 45378 48076 45388 48132
rect 45444 48076 45724 48132
rect 45780 48076 45790 48132
rect 10742 47964 10780 48020
rect 10836 47964 10846 48020
rect 18050 47964 18060 48020
rect 18116 47964 19516 48020
rect 19572 47964 20300 48020
rect 20356 47964 20366 48020
rect 34290 47964 34300 48020
rect 34356 47964 35196 48020
rect 35252 47964 35262 48020
rect 45154 47852 45164 47908
rect 45220 47852 46620 47908
rect 46676 47852 46686 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 13010 47740 13020 47796
rect 13076 47740 13356 47796
rect 13412 47740 13422 47796
rect 20962 47740 20972 47796
rect 21028 47740 33068 47796
rect 33124 47740 33134 47796
rect 3602 47628 3612 47684
rect 3668 47628 4732 47684
rect 4788 47628 4798 47684
rect 40226 47628 40236 47684
rect 40292 47628 41804 47684
rect 41860 47628 42812 47684
rect 42868 47628 42878 47684
rect 3378 47516 3388 47572
rect 3444 47516 3836 47572
rect 3892 47516 15148 47572
rect 17714 47516 17724 47572
rect 17780 47516 19740 47572
rect 19796 47516 22652 47572
rect 22708 47516 22718 47572
rect 23874 47516 23884 47572
rect 23940 47516 24556 47572
rect 24612 47516 24622 47572
rect 25106 47516 25116 47572
rect 25172 47516 25676 47572
rect 25732 47516 25742 47572
rect 26226 47516 26236 47572
rect 26292 47516 26572 47572
rect 26628 47516 31724 47572
rect 31780 47516 31790 47572
rect 32946 47516 32956 47572
rect 33012 47516 33628 47572
rect 33684 47516 34748 47572
rect 34804 47516 34814 47572
rect 38994 47516 39004 47572
rect 39060 47516 39900 47572
rect 39956 47516 39966 47572
rect 2482 47404 2492 47460
rect 2548 47404 2828 47460
rect 2884 47404 2894 47460
rect 4162 47404 4172 47460
rect 4228 47404 4844 47460
rect 4900 47404 4910 47460
rect 8194 47404 8204 47460
rect 8260 47404 10556 47460
rect 10612 47404 10622 47460
rect 2828 47124 2884 47404
rect 15092 47348 15148 47516
rect 23426 47404 23436 47460
rect 23492 47404 25228 47460
rect 25284 47404 25294 47460
rect 33842 47404 33852 47460
rect 33908 47404 34972 47460
rect 35028 47404 35038 47460
rect 39004 47404 39788 47460
rect 39844 47404 39854 47460
rect 39004 47348 39060 47404
rect 4386 47292 4396 47348
rect 4452 47292 4956 47348
rect 5012 47292 5022 47348
rect 15092 47292 24276 47348
rect 24220 47236 24276 47292
rect 25900 47292 27580 47348
rect 27636 47292 27646 47348
rect 30258 47292 30268 47348
rect 30324 47292 30716 47348
rect 30772 47292 32284 47348
rect 32340 47292 32956 47348
rect 33012 47292 33022 47348
rect 38882 47292 38892 47348
rect 38948 47292 39060 47348
rect 39330 47292 39340 47348
rect 39396 47292 40292 47348
rect 40450 47292 40460 47348
rect 40516 47292 40908 47348
rect 40964 47292 40974 47348
rect 25900 47236 25956 47292
rect 3332 47180 7476 47236
rect 7606 47180 7644 47236
rect 7700 47180 7710 47236
rect 9202 47180 9212 47236
rect 9268 47180 10892 47236
rect 10948 47180 10958 47236
rect 20290 47180 20300 47236
rect 20356 47180 20748 47236
rect 20804 47180 20814 47236
rect 22194 47180 22204 47236
rect 22260 47180 22988 47236
rect 23044 47180 23054 47236
rect 23314 47180 23324 47236
rect 23380 47180 23996 47236
rect 24052 47180 24062 47236
rect 24220 47180 25956 47236
rect 26114 47180 26124 47236
rect 26180 47180 26190 47236
rect 26786 47180 26796 47236
rect 26852 47180 26908 47292
rect 40236 47236 40292 47292
rect 38098 47180 38108 47236
rect 38164 47180 38444 47236
rect 38500 47180 39676 47236
rect 39732 47180 39742 47236
rect 40226 47180 40236 47236
rect 40292 47180 40572 47236
rect 40628 47180 40638 47236
rect 40786 47180 40796 47236
rect 40852 47180 42252 47236
rect 42308 47180 42812 47236
rect 42868 47180 42878 47236
rect 3332 47124 3388 47180
rect 7420 47124 7476 47180
rect 26124 47124 26180 47180
rect 2828 47068 3388 47124
rect 4834 47068 4844 47124
rect 4900 47068 5404 47124
rect 5460 47068 5470 47124
rect 7420 47068 13356 47124
rect 13412 47068 13422 47124
rect 22642 47068 22652 47124
rect 22708 47068 22876 47124
rect 22932 47068 22942 47124
rect 26124 47068 28252 47124
rect 28308 47068 28588 47124
rect 28644 47068 28654 47124
rect 33842 47068 33852 47124
rect 33908 47068 38780 47124
rect 38836 47068 39564 47124
rect 39620 47068 39630 47124
rect 41010 47068 41020 47124
rect 41076 47068 41804 47124
rect 41860 47068 41870 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 8754 46956 8764 47012
rect 8820 46956 15708 47012
rect 15764 46956 15774 47012
rect 20412 46956 24892 47012
rect 24948 46956 24958 47012
rect 20412 46900 20468 46956
rect 1474 46844 1484 46900
rect 1540 46844 6748 46900
rect 6804 46844 7532 46900
rect 7588 46844 8316 46900
rect 8372 46844 8382 46900
rect 9874 46844 9884 46900
rect 9940 46844 10668 46900
rect 10724 46844 11564 46900
rect 11620 46844 13468 46900
rect 13524 46844 13692 46900
rect 13748 46844 13758 46900
rect 15474 46844 15484 46900
rect 15540 46844 15932 46900
rect 15988 46844 15998 46900
rect 17490 46844 17500 46900
rect 17556 46844 19068 46900
rect 19124 46844 20468 46900
rect 26562 46844 26572 46900
rect 26628 46844 26684 46900
rect 26740 46844 26750 46900
rect 46610 46844 46620 46900
rect 46676 46844 46956 46900
rect 47012 46844 47022 46900
rect 5394 46732 5404 46788
rect 5460 46732 5740 46788
rect 5796 46732 5806 46788
rect 8978 46732 8988 46788
rect 9044 46732 11228 46788
rect 11284 46732 11294 46788
rect 22978 46732 22988 46788
rect 23044 46732 23772 46788
rect 23828 46732 24220 46788
rect 24276 46732 24286 46788
rect 29138 46732 29148 46788
rect 29204 46732 29596 46788
rect 29652 46732 29662 46788
rect 33170 46732 33180 46788
rect 33236 46732 33628 46788
rect 33684 46732 33694 46788
rect 3826 46620 3836 46676
rect 3892 46620 4172 46676
rect 4228 46620 4238 46676
rect 20738 46620 20748 46676
rect 20804 46620 21196 46676
rect 21252 46620 21262 46676
rect 23090 46620 23100 46676
rect 23156 46620 23166 46676
rect 24546 46620 24556 46676
rect 24612 46620 25116 46676
rect 25172 46620 25182 46676
rect 34514 46620 34524 46676
rect 34580 46620 34748 46676
rect 34804 46620 34814 46676
rect 42690 46620 42700 46676
rect 42756 46620 43820 46676
rect 43876 46620 44156 46676
rect 44212 46620 44222 46676
rect 23100 46564 23156 46620
rect 11666 46508 11676 46564
rect 11732 46508 22652 46564
rect 22708 46508 23156 46564
rect 25330 46508 25340 46564
rect 25396 46508 27468 46564
rect 27524 46508 27534 46564
rect 29586 46508 29596 46564
rect 29652 46508 31500 46564
rect 31556 46508 31566 46564
rect 15810 46396 15820 46452
rect 15876 46396 17500 46452
rect 17556 46396 17566 46452
rect 20626 46396 20636 46452
rect 20692 46396 21420 46452
rect 21476 46396 21486 46452
rect 25554 46396 25564 46452
rect 25620 46396 26236 46452
rect 26292 46396 26302 46452
rect 26646 46396 26684 46452
rect 26740 46396 26750 46452
rect 34598 46396 34636 46452
rect 34692 46396 34702 46452
rect 5842 46284 5852 46340
rect 5908 46284 10556 46340
rect 10612 46284 11116 46340
rect 11172 46284 11182 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 15698 46172 15708 46228
rect 15764 46172 22764 46228
rect 22820 46172 22830 46228
rect 37510 46172 37548 46228
rect 37604 46172 37614 46228
rect 12562 46060 12572 46116
rect 12628 46060 24332 46116
rect 24388 46060 24892 46116
rect 24948 46060 24958 46116
rect 0 45920 800 46032
rect 49200 46004 50000 46032
rect 15922 45948 15932 46004
rect 15988 45948 17164 46004
rect 17220 45948 17230 46004
rect 20402 45948 20412 46004
rect 20468 45948 21532 46004
rect 21588 45948 21598 46004
rect 22642 45948 22652 46004
rect 22708 45948 22764 46004
rect 22820 45948 22830 46004
rect 26236 45948 26796 46004
rect 26852 45948 26908 46004
rect 26964 45948 26974 46004
rect 39218 45948 39228 46004
rect 39284 45948 39900 46004
rect 39956 45948 40572 46004
rect 40628 45948 41020 46004
rect 41076 45948 41086 46004
rect 43698 45948 43708 46004
rect 43764 45948 45164 46004
rect 45220 45948 45230 46004
rect 48066 45948 48076 46004
rect 48132 45948 50000 46004
rect 5730 45836 5740 45892
rect 5796 45836 7980 45892
rect 8036 45836 8046 45892
rect 9986 45836 9996 45892
rect 10052 45836 14140 45892
rect 14196 45836 14812 45892
rect 14868 45836 15036 45892
rect 15092 45836 15102 45892
rect 16604 45836 23548 45892
rect 23604 45836 23884 45892
rect 23940 45836 23950 45892
rect 24434 45836 24444 45892
rect 24500 45836 25676 45892
rect 25732 45836 25742 45892
rect 16604 45780 16660 45836
rect 26236 45780 26292 45948
rect 49200 45920 50000 45948
rect 40786 45836 40796 45892
rect 40852 45836 42252 45892
rect 42308 45836 42318 45892
rect 43250 45836 43260 45892
rect 43316 45836 44044 45892
rect 44100 45836 44110 45892
rect 9314 45724 9324 45780
rect 9380 45724 9548 45780
rect 9604 45724 10220 45780
rect 10276 45724 10286 45780
rect 11218 45724 11228 45780
rect 11284 45724 11900 45780
rect 11956 45724 13692 45780
rect 13748 45724 13758 45780
rect 14466 45724 14476 45780
rect 14532 45724 16604 45780
rect 16660 45724 16670 45780
rect 20738 45724 20748 45780
rect 20804 45724 21308 45780
rect 21364 45724 21868 45780
rect 21924 45724 21934 45780
rect 22866 45724 22876 45780
rect 22932 45724 23436 45780
rect 23492 45724 23502 45780
rect 26226 45724 26236 45780
rect 26292 45724 26302 45780
rect 30818 45724 30828 45780
rect 30884 45724 32060 45780
rect 32116 45724 32126 45780
rect 12226 45612 12236 45668
rect 12292 45612 15596 45668
rect 15652 45612 15662 45668
rect 18946 45612 18956 45668
rect 19012 45612 19628 45668
rect 19684 45612 20188 45668
rect 20244 45612 21532 45668
rect 21588 45612 21598 45668
rect 29222 45612 29260 45668
rect 29316 45612 29326 45668
rect 32722 45612 32732 45668
rect 32788 45612 33404 45668
rect 33460 45612 33470 45668
rect 36866 45612 36876 45668
rect 36932 45612 41916 45668
rect 41972 45612 41982 45668
rect 10994 45500 11004 45556
rect 11060 45500 12348 45556
rect 12404 45500 12414 45556
rect 29026 45500 29036 45556
rect 29092 45500 29708 45556
rect 29764 45500 29774 45556
rect 31154 45500 31164 45556
rect 31220 45500 32284 45556
rect 32340 45500 32350 45556
rect 37762 45500 37772 45556
rect 37828 45500 40460 45556
rect 40516 45500 41244 45556
rect 41300 45500 41310 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 15250 45388 15260 45444
rect 15316 45388 15708 45444
rect 15764 45388 15774 45444
rect 24630 45388 24668 45444
rect 24724 45388 24734 45444
rect 28690 45388 28700 45444
rect 28756 45388 29484 45444
rect 29540 45388 29550 45444
rect 30258 45388 30268 45444
rect 30324 45388 33628 45444
rect 33684 45388 33694 45444
rect 36754 45388 36764 45444
rect 36820 45388 36830 45444
rect 38658 45388 38668 45444
rect 38724 45388 38762 45444
rect 36764 45332 36820 45388
rect 1922 45276 1932 45332
rect 1988 45276 2380 45332
rect 2436 45276 2828 45332
rect 2884 45276 3668 45332
rect 3826 45276 3836 45332
rect 3892 45276 6860 45332
rect 6916 45276 6926 45332
rect 7074 45276 7084 45332
rect 7140 45276 8540 45332
rect 8596 45276 8606 45332
rect 8866 45276 8876 45332
rect 8932 45276 8942 45332
rect 13346 45276 13356 45332
rect 13412 45276 14588 45332
rect 14644 45276 14654 45332
rect 15138 45276 15148 45332
rect 15204 45276 16716 45332
rect 16772 45276 16782 45332
rect 17826 45276 17836 45332
rect 17892 45276 18396 45332
rect 18452 45276 18462 45332
rect 19366 45276 19404 45332
rect 19460 45276 19470 45332
rect 20300 45276 22484 45332
rect 23314 45276 23324 45332
rect 23380 45276 25452 45332
rect 25508 45276 25518 45332
rect 27916 45276 28140 45332
rect 28196 45276 30492 45332
rect 30548 45276 30558 45332
rect 30930 45276 30940 45332
rect 30996 45276 31388 45332
rect 31444 45276 31454 45332
rect 35298 45276 35308 45332
rect 35364 45276 37324 45332
rect 37380 45276 37390 45332
rect 38612 45276 40348 45332
rect 40404 45276 40414 45332
rect 3612 45220 3668 45276
rect 8876 45220 8932 45276
rect 2258 45164 2268 45220
rect 2324 45164 3164 45220
rect 3220 45164 3388 45220
rect 3444 45164 3454 45220
rect 3612 45164 5180 45220
rect 5236 45164 5246 45220
rect 8306 45164 8316 45220
rect 8372 45164 8932 45220
rect 16716 45220 16772 45276
rect 20300 45220 20356 45276
rect 22428 45220 22484 45276
rect 16716 45164 20356 45220
rect 20514 45164 20524 45220
rect 20580 45164 22204 45220
rect 22260 45164 22270 45220
rect 22428 45164 24444 45220
rect 24500 45164 25228 45220
rect 25284 45164 25294 45220
rect 25890 45164 25900 45220
rect 25956 45164 27132 45220
rect 27188 45164 27198 45220
rect 27916 45108 27972 45276
rect 30034 45164 30044 45220
rect 30100 45164 30828 45220
rect 30884 45164 32060 45220
rect 32116 45164 32126 45220
rect 34738 45164 34748 45220
rect 34804 45164 35644 45220
rect 35700 45164 35710 45220
rect 35858 45164 35868 45220
rect 35924 45164 36204 45220
rect 36260 45164 36270 45220
rect 38612 45108 38668 45276
rect 39330 45164 39340 45220
rect 39396 45164 39900 45220
rect 39956 45164 40124 45220
rect 40180 45164 41692 45220
rect 41748 45164 42028 45220
rect 42084 45164 42094 45220
rect 2482 45052 2492 45108
rect 2548 45052 3388 45108
rect 7858 45052 7868 45108
rect 7924 45052 8876 45108
rect 8932 45052 9772 45108
rect 9828 45052 9838 45108
rect 15698 45052 15708 45108
rect 15764 45052 16716 45108
rect 16772 45052 17500 45108
rect 17556 45052 17566 45108
rect 21858 45052 21868 45108
rect 21924 45052 22652 45108
rect 22708 45052 22718 45108
rect 25778 45052 25788 45108
rect 25844 45052 27972 45108
rect 29474 45052 29484 45108
rect 29540 45052 29932 45108
rect 29988 45052 29998 45108
rect 30146 45052 30156 45108
rect 30212 45052 30716 45108
rect 30772 45052 31836 45108
rect 31892 45052 31902 45108
rect 33058 45052 33068 45108
rect 33124 45052 38332 45108
rect 38388 45052 38668 45108
rect 40002 45052 40012 45108
rect 40068 45052 41356 45108
rect 41412 45052 41422 45108
rect 3332 44996 3388 45052
rect 3332 44940 3612 44996
rect 3668 44940 3678 44996
rect 7410 44940 7420 44996
rect 7476 44940 7980 44996
rect 8036 44940 8046 44996
rect 8642 44940 8652 44996
rect 8708 44940 8718 44996
rect 9090 44940 9100 44996
rect 9156 44940 9660 44996
rect 9716 44940 9726 44996
rect 19618 44940 19628 44996
rect 19684 44940 20244 44996
rect 20402 44940 20412 44996
rect 20468 44940 21420 44996
rect 21476 44940 22204 44996
rect 22260 44940 22270 44996
rect 23650 44940 23660 44996
rect 23716 44940 25564 44996
rect 25620 44940 26012 44996
rect 26068 44940 26078 44996
rect 34290 44940 34300 44996
rect 34356 44940 35532 44996
rect 35588 44940 35598 44996
rect 37426 44940 37436 44996
rect 37492 44940 37884 44996
rect 37940 44940 37950 44996
rect 38108 44940 38668 44996
rect 38724 44940 39676 44996
rect 39732 44940 39742 44996
rect 45042 44940 45052 44996
rect 45108 44940 45724 44996
rect 45780 44940 45790 44996
rect 8652 44772 8708 44940
rect 20188 44884 20244 44940
rect 38108 44884 38164 44940
rect 14130 44828 14140 44884
rect 14196 44828 14206 44884
rect 18050 44828 18060 44884
rect 18116 44828 19852 44884
rect 19908 44828 19918 44884
rect 20178 44828 20188 44884
rect 20244 44828 21196 44884
rect 21252 44828 21756 44884
rect 21812 44828 21822 44884
rect 29670 44828 29708 44884
rect 29764 44828 37772 44884
rect 37828 44828 37838 44884
rect 37986 44828 37996 44884
rect 38052 44828 38164 44884
rect 45826 44828 45836 44884
rect 45892 44828 46508 44884
rect 46564 44828 46574 44884
rect 8418 44716 8428 44772
rect 8484 44716 8708 44772
rect 14140 44772 14196 44828
rect 14140 44716 21420 44772
rect 21476 44716 21486 44772
rect 40674 44716 40684 44772
rect 40740 44716 42588 44772
rect 42644 44716 42654 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 8306 44604 8316 44660
rect 8372 44604 8652 44660
rect 8708 44604 8718 44660
rect 14140 44436 14196 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 14578 44604 14588 44660
rect 14644 44604 20188 44660
rect 20244 44604 21532 44660
rect 21588 44604 21598 44660
rect 22306 44604 22316 44660
rect 22372 44604 22428 44660
rect 22484 44604 22494 44660
rect 37762 44604 37772 44660
rect 37828 44604 38108 44660
rect 38164 44604 38174 44660
rect 38434 44604 38444 44660
rect 38500 44604 38668 44660
rect 38724 44604 38734 44660
rect 16594 44492 16604 44548
rect 16660 44492 22372 44548
rect 23090 44492 23100 44548
rect 23156 44492 25116 44548
rect 25172 44492 25182 44548
rect 29698 44492 29708 44548
rect 29764 44492 37996 44548
rect 38052 44492 38062 44548
rect 41458 44492 41468 44548
rect 41524 44492 42588 44548
rect 42644 44492 42654 44548
rect 22316 44436 22372 44492
rect 3910 44380 3948 44436
rect 4004 44380 4014 44436
rect 6290 44380 6300 44436
rect 6356 44380 7644 44436
rect 7700 44380 7710 44436
rect 10434 44380 10444 44436
rect 10500 44380 10892 44436
rect 10948 44380 10958 44436
rect 12012 44380 13916 44436
rect 13972 44380 14196 44436
rect 20402 44380 20412 44436
rect 20468 44380 21532 44436
rect 21588 44380 22092 44436
rect 22148 44380 22158 44436
rect 22316 44380 23548 44436
rect 23604 44380 23996 44436
rect 24052 44380 24062 44436
rect 32386 44380 32396 44436
rect 32452 44380 34300 44436
rect 34356 44380 34366 44436
rect 41570 44380 41580 44436
rect 41636 44380 41748 44436
rect 45938 44380 45948 44436
rect 46004 44380 47068 44436
rect 47124 44380 47134 44436
rect 12012 44324 12068 44380
rect 3714 44268 3724 44324
rect 3780 44268 4172 44324
rect 4228 44268 12068 44324
rect 12898 44268 12908 44324
rect 12964 44268 13580 44324
rect 13636 44268 13646 44324
rect 16370 44268 16380 44324
rect 16436 44268 17052 44324
rect 17108 44268 17118 44324
rect 17826 44268 17836 44324
rect 17892 44268 18732 44324
rect 18788 44268 20300 44324
rect 20356 44268 20366 44324
rect 24658 44268 24668 44324
rect 24724 44268 24892 44324
rect 24948 44268 24958 44324
rect 30706 44268 30716 44324
rect 30772 44268 31948 44324
rect 32004 44268 32014 44324
rect 34402 44268 34412 44324
rect 34468 44268 34972 44324
rect 35028 44268 35038 44324
rect 36418 44268 36428 44324
rect 36484 44268 37100 44324
rect 37156 44268 37166 44324
rect 37874 44268 37884 44324
rect 37940 44268 38668 44324
rect 38724 44268 38734 44324
rect 41234 44268 41244 44324
rect 41300 44268 41356 44324
rect 41412 44268 41422 44324
rect 34972 44212 35028 44268
rect 3378 44156 3388 44212
rect 3444 44156 3948 44212
rect 4004 44156 4014 44212
rect 13794 44156 13804 44212
rect 13860 44156 14588 44212
rect 14644 44156 16828 44212
rect 16884 44156 17500 44212
rect 17556 44156 17566 44212
rect 22418 44156 22428 44212
rect 22484 44156 23884 44212
rect 23940 44156 23950 44212
rect 34972 44156 40684 44212
rect 40740 44156 40750 44212
rect 41010 44156 41020 44212
rect 41076 44156 41086 44212
rect 2594 44044 2604 44100
rect 2660 44044 4060 44100
rect 4116 44044 4126 44100
rect 4722 44044 4732 44100
rect 4788 44044 4956 44100
rect 5012 44044 5022 44100
rect 5506 44044 5516 44100
rect 5572 44044 6524 44100
rect 6580 44044 7084 44100
rect 7140 44044 7150 44100
rect 12338 44044 12348 44100
rect 12404 44044 13356 44100
rect 13412 44044 13422 44100
rect 21410 44044 21420 44100
rect 21476 44044 21756 44100
rect 21812 44044 22204 44100
rect 22260 44044 22988 44100
rect 23044 44044 23054 44100
rect 23538 44044 23548 44100
rect 23604 44044 24108 44100
rect 24164 44044 24174 44100
rect 4732 43988 4788 44044
rect 3602 43932 3612 43988
rect 3668 43932 4788 43988
rect 14466 43932 14476 43988
rect 14532 43932 15036 43988
rect 15092 43932 15102 43988
rect 21970 43932 21980 43988
rect 22036 43932 22764 43988
rect 22820 43932 23324 43988
rect 23380 43932 23390 43988
rect 36082 43932 36092 43988
rect 36148 43932 39900 43988
rect 39956 43932 40796 43988
rect 40852 43932 40862 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 41020 43876 41076 44156
rect 41692 43988 41748 44380
rect 41682 43932 41692 43988
rect 41748 43932 41758 43988
rect 6626 43820 6636 43876
rect 6692 43820 6702 43876
rect 18918 43820 18956 43876
rect 19012 43820 19022 43876
rect 20178 43820 20188 43876
rect 20244 43820 23772 43876
rect 23828 43820 24108 43876
rect 24164 43820 24174 43876
rect 30930 43820 30940 43876
rect 30996 43820 40684 43876
rect 40740 43820 41076 43876
rect 6636 43764 6692 43820
rect 6636 43708 6916 43764
rect 10098 43708 10108 43764
rect 10164 43708 13356 43764
rect 13412 43708 13422 43764
rect 15362 43708 15372 43764
rect 15428 43708 16604 43764
rect 16660 43708 16670 43764
rect 24658 43708 24668 43764
rect 24724 43708 25340 43764
rect 25396 43708 26236 43764
rect 26292 43708 26302 43764
rect 37762 43708 37772 43764
rect 37828 43708 37996 43764
rect 38052 43708 40348 43764
rect 40404 43708 41020 43764
rect 41076 43708 41086 43764
rect 42018 43708 42028 43764
rect 42084 43708 42812 43764
rect 42868 43708 42878 43764
rect 46610 43708 46620 43764
rect 46676 43708 46686 43764
rect 47730 43708 47740 43764
rect 47796 43708 47806 43764
rect 2258 43596 2268 43652
rect 2324 43596 3612 43652
rect 3668 43596 4732 43652
rect 4788 43596 4798 43652
rect 0 43456 800 43568
rect 6860 43540 6916 43708
rect 46620 43652 46676 43708
rect 8978 43596 8988 43652
rect 9044 43596 9324 43652
rect 9380 43596 9390 43652
rect 10994 43596 11004 43652
rect 11060 43596 12012 43652
rect 12068 43596 12078 43652
rect 22726 43596 22764 43652
rect 22820 43596 22830 43652
rect 24210 43596 24220 43652
rect 24276 43596 25116 43652
rect 25172 43596 25182 43652
rect 29698 43596 29708 43652
rect 29764 43596 30044 43652
rect 30100 43596 30110 43652
rect 46620 43596 47404 43652
rect 47460 43596 47470 43652
rect 47740 43540 47796 43708
rect 49200 43540 50000 43568
rect 2370 43484 2380 43540
rect 2436 43484 4620 43540
rect 4676 43484 5852 43540
rect 5908 43484 6636 43540
rect 6692 43484 6702 43540
rect 6860 43484 9100 43540
rect 9156 43484 9166 43540
rect 9538 43484 9548 43540
rect 9604 43484 10556 43540
rect 10612 43484 10622 43540
rect 11666 43484 11676 43540
rect 11732 43484 12796 43540
rect 12852 43484 13468 43540
rect 13524 43484 13534 43540
rect 14018 43484 14028 43540
rect 14084 43484 15260 43540
rect 15316 43484 16828 43540
rect 16884 43484 16894 43540
rect 20748 43484 20972 43540
rect 21028 43484 21038 43540
rect 25554 43484 25564 43540
rect 25620 43484 27020 43540
rect 27076 43484 27086 43540
rect 41570 43484 41580 43540
rect 41636 43484 43036 43540
rect 43092 43484 43102 43540
rect 46610 43484 46620 43540
rect 46676 43484 47180 43540
rect 47236 43484 47246 43540
rect 47740 43484 50000 43540
rect 20748 43428 20804 43484
rect 49200 43456 50000 43484
rect 4722 43372 4732 43428
rect 4788 43372 7084 43428
rect 7140 43372 7150 43428
rect 8530 43372 8540 43428
rect 8596 43372 9660 43428
rect 9716 43372 9726 43428
rect 20738 43372 20748 43428
rect 20804 43372 20814 43428
rect 25330 43372 25340 43428
rect 25396 43372 27244 43428
rect 27300 43372 27310 43428
rect 38994 43372 39004 43428
rect 39060 43372 39900 43428
rect 39956 43372 39966 43428
rect 45266 43372 45276 43428
rect 45332 43372 46508 43428
rect 46564 43372 46574 43428
rect 2930 43260 2940 43316
rect 2996 43260 9436 43316
rect 9492 43260 9502 43316
rect 18610 43260 18620 43316
rect 18676 43260 19180 43316
rect 19236 43260 19852 43316
rect 19908 43260 19918 43316
rect 38658 43260 38668 43316
rect 38724 43260 38762 43316
rect 5058 43148 5068 43204
rect 5124 43148 9548 43204
rect 9604 43148 9614 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 5730 43036 5740 43092
rect 5796 43036 6188 43092
rect 6244 43036 6254 43092
rect 6934 43036 6972 43092
rect 7028 43036 7038 43092
rect 7074 42924 7084 42980
rect 7140 42924 8876 42980
rect 8932 42924 8942 42980
rect 22082 42924 22092 42980
rect 22148 42924 24444 42980
rect 24500 42924 26908 42980
rect 26964 42924 26974 42980
rect 5394 42812 5404 42868
rect 5460 42812 6468 42868
rect 11218 42812 11228 42868
rect 11284 42812 12796 42868
rect 12852 42812 12862 42868
rect 15586 42812 15596 42868
rect 15652 42812 16380 42868
rect 16436 42812 16446 42868
rect 41206 42812 41244 42868
rect 41300 42812 41310 42868
rect 41878 42812 41916 42868
rect 41972 42812 41982 42868
rect 3714 42700 3724 42756
rect 3780 42700 4956 42756
rect 5012 42700 5628 42756
rect 5684 42700 5694 42756
rect 6412 42644 6468 42812
rect 6626 42700 6636 42756
rect 6692 42700 7308 42756
rect 7364 42700 7374 42756
rect 26226 42700 26236 42756
rect 26292 42700 26684 42756
rect 26740 42700 27692 42756
rect 27748 42700 27758 42756
rect 6412 42588 6972 42644
rect 7028 42588 7308 42644
rect 7364 42588 7374 42644
rect 15092 42588 20076 42644
rect 20132 42588 20142 42644
rect 20290 42588 20300 42644
rect 20356 42588 20972 42644
rect 21028 42588 21038 42644
rect 33506 42588 33516 42644
rect 33572 42588 33964 42644
rect 34020 42588 34030 42644
rect 15092 42532 15148 42588
rect 5170 42476 5180 42532
rect 5236 42476 5246 42532
rect 5394 42476 5404 42532
rect 5460 42476 5740 42532
rect 5796 42476 5806 42532
rect 10210 42476 10220 42532
rect 10276 42476 10556 42532
rect 10612 42476 10892 42532
rect 10948 42476 15148 42532
rect 18834 42476 18844 42532
rect 18900 42476 19740 42532
rect 19796 42476 19806 42532
rect 20188 42476 24892 42532
rect 24948 42476 24958 42532
rect 37426 42476 37436 42532
rect 37492 42476 38108 42532
rect 38164 42476 39004 42532
rect 39060 42476 39676 42532
rect 39732 42476 39742 42532
rect 41906 42476 41916 42532
rect 41972 42476 42476 42532
rect 42532 42476 42542 42532
rect 5180 42308 5236 42476
rect 6738 42364 6748 42420
rect 6804 42364 7308 42420
rect 7364 42364 7374 42420
rect 9986 42364 9996 42420
rect 10052 42364 15932 42420
rect 15988 42364 16492 42420
rect 16548 42364 16558 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 5180 42252 15036 42308
rect 15092 42252 15102 42308
rect 15474 42252 15484 42308
rect 15540 42252 16380 42308
rect 16436 42252 16446 42308
rect 20188 42196 20244 42476
rect 24546 42364 24556 42420
rect 24612 42364 25676 42420
rect 25732 42364 28028 42420
rect 28084 42364 41412 42420
rect 41356 42308 41412 42364
rect 36306 42252 36316 42308
rect 36372 42252 36652 42308
rect 36708 42252 36718 42308
rect 41356 42252 44380 42308
rect 44436 42252 44446 42308
rect 11890 42140 11900 42196
rect 11956 42140 20244 42196
rect 33394 42140 33404 42196
rect 33460 42140 39340 42196
rect 39396 42140 39406 42196
rect 45826 42140 45836 42196
rect 45892 42140 45902 42196
rect 45836 42084 45892 42140
rect 11778 42028 11788 42084
rect 11844 42028 12348 42084
rect 12404 42028 12414 42084
rect 12898 42028 12908 42084
rect 12964 42028 16044 42084
rect 16100 42028 16110 42084
rect 31938 42028 31948 42084
rect 32004 42028 33180 42084
rect 33236 42028 33852 42084
rect 33908 42028 34412 42084
rect 34468 42028 34478 42084
rect 36754 42028 36764 42084
rect 36820 42028 38444 42084
rect 38500 42028 38510 42084
rect 40674 42028 40684 42084
rect 40740 42028 40750 42084
rect 45836 42028 46396 42084
rect 46452 42028 46462 42084
rect 40684 41972 40740 42028
rect 3154 41916 3164 41972
rect 3220 41916 5572 41972
rect 7634 41916 7644 41972
rect 7700 41916 8540 41972
rect 8596 41916 8606 41972
rect 18946 41916 18956 41972
rect 19012 41916 19628 41972
rect 19684 41916 20300 41972
rect 20356 41916 20366 41972
rect 21522 41916 21532 41972
rect 21588 41916 21980 41972
rect 22036 41916 22046 41972
rect 22306 41916 22316 41972
rect 22372 41916 22652 41972
rect 22708 41916 22988 41972
rect 23044 41916 23054 41972
rect 24322 41916 24332 41972
rect 24388 41916 25116 41972
rect 25172 41916 25182 41972
rect 26450 41916 26460 41972
rect 26516 41916 26684 41972
rect 26740 41916 26750 41972
rect 27346 41916 27356 41972
rect 27412 41916 29820 41972
rect 29876 41916 29886 41972
rect 31490 41916 31500 41972
rect 31556 41916 32396 41972
rect 32452 41916 32462 41972
rect 32834 41916 32844 41972
rect 32900 41916 33292 41972
rect 33348 41916 33358 41972
rect 33516 41916 35420 41972
rect 35476 41916 35486 41972
rect 36082 41916 36092 41972
rect 36148 41916 37436 41972
rect 37492 41916 37502 41972
rect 39442 41916 39452 41972
rect 39508 41916 40740 41972
rect 44930 41916 44940 41972
rect 44996 41916 46508 41972
rect 46564 41916 46574 41972
rect 5516 41636 5572 41916
rect 33516 41860 33572 41916
rect 8950 41804 8988 41860
rect 9044 41804 9996 41860
rect 10052 41804 10062 41860
rect 15586 41804 15596 41860
rect 15652 41804 16380 41860
rect 16436 41804 16446 41860
rect 20066 41804 20076 41860
rect 20132 41804 21420 41860
rect 21476 41804 21486 41860
rect 24210 41804 24220 41860
rect 24276 41804 24668 41860
rect 24724 41804 24734 41860
rect 25330 41804 25340 41860
rect 25396 41804 27468 41860
rect 27524 41804 27534 41860
rect 29586 41804 29596 41860
rect 29652 41804 31948 41860
rect 32004 41804 32014 41860
rect 33170 41804 33180 41860
rect 33236 41804 33572 41860
rect 34290 41804 34300 41860
rect 34356 41804 38556 41860
rect 38612 41804 38622 41860
rect 16258 41692 16268 41748
rect 16324 41692 21868 41748
rect 21924 41692 21934 41748
rect 22754 41692 22764 41748
rect 22820 41692 23660 41748
rect 23716 41692 23726 41748
rect 34402 41692 34412 41748
rect 34468 41692 35532 41748
rect 35588 41692 35598 41748
rect 45714 41692 45724 41748
rect 45780 41692 46172 41748
rect 46228 41692 46238 41748
rect 5506 41580 5516 41636
rect 5572 41580 6188 41636
rect 6244 41580 7084 41636
rect 7140 41580 22092 41636
rect 22148 41580 22158 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 2706 41356 2716 41412
rect 2772 41356 8428 41412
rect 8484 41356 8494 41412
rect 24770 41356 24780 41412
rect 24836 41356 25452 41412
rect 25508 41356 25518 41412
rect 35074 41356 35084 41412
rect 35140 41356 36204 41412
rect 36260 41356 36270 41412
rect 21756 41244 23772 41300
rect 23828 41244 23838 41300
rect 32386 41244 32396 41300
rect 32452 41244 34972 41300
rect 35028 41244 36092 41300
rect 36148 41244 37324 41300
rect 37380 41244 37390 41300
rect 40002 41244 40012 41300
rect 40068 41244 40572 41300
rect 40628 41244 41580 41300
rect 41636 41244 41646 41300
rect 21756 41188 21812 41244
rect 16370 41132 16380 41188
rect 16436 41132 17276 41188
rect 17332 41132 17342 41188
rect 18918 41132 18956 41188
rect 19012 41132 19022 41188
rect 19170 41132 19180 41188
rect 19236 41132 19628 41188
rect 19684 41132 19694 41188
rect 21746 41132 21756 41188
rect 21812 41132 21822 41188
rect 21970 41132 21980 41188
rect 22036 41132 23436 41188
rect 23492 41132 23502 41188
rect 32946 41132 32956 41188
rect 33012 41132 33964 41188
rect 34020 41132 34524 41188
rect 34580 41132 34590 41188
rect 34748 41132 35756 41188
rect 35812 41132 35822 41188
rect 38882 41132 38892 41188
rect 38948 41132 39788 41188
rect 39844 41132 41244 41188
rect 41300 41132 41310 41188
rect 0 40992 800 41104
rect 34748 41076 34804 41132
rect 49200 41076 50000 41104
rect 2146 41020 2156 41076
rect 2212 41020 3500 41076
rect 3556 41020 3724 41076
rect 3780 41020 3790 41076
rect 5058 41020 5068 41076
rect 5124 41020 6076 41076
rect 6132 41020 6142 41076
rect 6738 41020 6748 41076
rect 6804 41020 6972 41076
rect 7028 41020 7420 41076
rect 7476 41020 7486 41076
rect 16482 41020 16492 41076
rect 16548 41020 20636 41076
rect 20692 41020 21644 41076
rect 21700 41020 21710 41076
rect 22390 41020 22428 41076
rect 22484 41020 22494 41076
rect 22876 41020 23884 41076
rect 23940 41020 23950 41076
rect 22876 40964 22932 41020
rect 26852 40964 26908 41076
rect 26964 41020 31052 41076
rect 31108 41020 31388 41076
rect 31444 41020 31454 41076
rect 33730 41020 33740 41076
rect 33796 41020 34804 41076
rect 35410 41020 35420 41076
rect 35476 41020 36316 41076
rect 36372 41020 36382 41076
rect 41570 41020 41580 41076
rect 41636 41020 42028 41076
rect 42084 41020 42700 41076
rect 42756 41020 42766 41076
rect 45378 41020 45388 41076
rect 45444 41020 46172 41076
rect 46228 41020 46238 41076
rect 48066 41020 48076 41076
rect 48132 41020 50000 41076
rect 49200 40992 50000 41020
rect 2482 40908 2492 40964
rect 2548 40908 3164 40964
rect 3220 40908 3230 40964
rect 8418 40908 8428 40964
rect 8484 40908 9772 40964
rect 9828 40908 9838 40964
rect 15474 40908 15484 40964
rect 15540 40908 22876 40964
rect 22932 40908 22942 40964
rect 23650 40908 23660 40964
rect 23716 40908 24052 40964
rect 24546 40908 24556 40964
rect 24612 40908 26908 40964
rect 34738 40908 34748 40964
rect 34804 40908 36204 40964
rect 36260 40908 36270 40964
rect 38546 40908 38556 40964
rect 38612 40908 39116 40964
rect 39172 40908 39182 40964
rect 7074 40796 7084 40852
rect 7140 40796 7196 40852
rect 7252 40796 7262 40852
rect 17042 40796 17052 40852
rect 17108 40796 18060 40852
rect 18116 40796 18126 40852
rect 22418 40796 22428 40852
rect 22484 40796 23548 40852
rect 23604 40796 23614 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 23996 40740 24052 40908
rect 31378 40796 31388 40852
rect 31444 40796 33516 40852
rect 33572 40796 33582 40852
rect 43586 40796 43596 40852
rect 43652 40796 45164 40852
rect 45220 40796 45230 40852
rect 23996 40684 24556 40740
rect 24612 40684 24622 40740
rect 26450 40684 26460 40740
rect 26516 40684 26526 40740
rect 30146 40684 30156 40740
rect 30212 40684 30940 40740
rect 30996 40684 31612 40740
rect 31668 40684 32396 40740
rect 32452 40684 38668 40740
rect 41234 40684 41244 40740
rect 41300 40684 41916 40740
rect 41972 40684 41982 40740
rect 26460 40628 26516 40684
rect 4722 40572 4732 40628
rect 4788 40572 5516 40628
rect 5572 40572 5582 40628
rect 8530 40572 8540 40628
rect 8596 40572 9660 40628
rect 9716 40572 9726 40628
rect 17490 40572 17500 40628
rect 17556 40572 26516 40628
rect 28662 40572 28700 40628
rect 28756 40572 28766 40628
rect 31938 40572 31948 40628
rect 32004 40572 33180 40628
rect 33236 40572 33246 40628
rect 34748 40572 35084 40628
rect 35140 40572 35150 40628
rect 34748 40516 34804 40572
rect 21522 40460 21532 40516
rect 21588 40460 22988 40516
rect 23044 40460 23054 40516
rect 23314 40460 23324 40516
rect 23380 40460 25396 40516
rect 25554 40460 25564 40516
rect 25620 40460 26460 40516
rect 26516 40460 26526 40516
rect 31164 40460 34804 40516
rect 38612 40516 38668 40684
rect 39106 40572 39116 40628
rect 39172 40572 39340 40628
rect 39396 40572 39788 40628
rect 39844 40572 40684 40628
rect 40740 40572 40750 40628
rect 41682 40572 41692 40628
rect 41748 40572 42252 40628
rect 42308 40572 42318 40628
rect 41692 40516 41748 40572
rect 38612 40460 40236 40516
rect 40292 40460 40302 40516
rect 40786 40460 40796 40516
rect 40852 40460 41748 40516
rect 44482 40460 44492 40516
rect 44548 40460 45388 40516
rect 45444 40460 45454 40516
rect 25340 40404 25396 40460
rect 31164 40404 31220 40460
rect 20178 40348 20188 40404
rect 20244 40348 20972 40404
rect 21028 40348 21038 40404
rect 21410 40348 21420 40404
rect 21476 40348 22652 40404
rect 22708 40348 22718 40404
rect 25330 40348 25340 40404
rect 25396 40348 25406 40404
rect 28690 40348 28700 40404
rect 28756 40348 28766 40404
rect 30818 40348 30828 40404
rect 30884 40348 31164 40404
rect 31220 40348 31230 40404
rect 32386 40348 32396 40404
rect 32452 40348 32732 40404
rect 32788 40348 32798 40404
rect 33170 40348 33180 40404
rect 33236 40348 34468 40404
rect 28700 40292 28756 40348
rect 34412 40292 34468 40348
rect 34748 40292 34804 40460
rect 35522 40348 35532 40404
rect 35588 40348 37436 40404
rect 37492 40348 37502 40404
rect 38882 40348 38892 40404
rect 38948 40348 43708 40404
rect 43764 40348 43932 40404
rect 43988 40348 43998 40404
rect 8306 40236 8316 40292
rect 8372 40236 10108 40292
rect 10164 40236 10174 40292
rect 16482 40236 16492 40292
rect 16548 40236 17500 40292
rect 17556 40236 17566 40292
rect 28700 40236 30380 40292
rect 30436 40236 30446 40292
rect 34402 40236 34412 40292
rect 34468 40236 34478 40292
rect 34626 40236 34636 40292
rect 34692 40236 34804 40292
rect 37538 40236 37548 40292
rect 37604 40236 38220 40292
rect 38276 40236 38556 40292
rect 38612 40236 38622 40292
rect 16146 40124 16156 40180
rect 16212 40124 16604 40180
rect 16660 40124 17276 40180
rect 17332 40124 17342 40180
rect 23650 40124 23660 40180
rect 23716 40124 25116 40180
rect 25172 40124 25182 40180
rect 32274 40124 32284 40180
rect 32340 40124 41580 40180
rect 41636 40124 41646 40180
rect 7522 40012 7532 40068
rect 7588 40012 8204 40068
rect 8260 40012 10556 40068
rect 10612 40012 10622 40068
rect 28662 40012 28700 40068
rect 28756 40012 28766 40068
rect 30370 40012 30380 40068
rect 30436 40012 32396 40068
rect 32452 40012 32462 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 21494 39900 21532 39956
rect 21588 39900 21598 39956
rect 43586 39900 43596 39956
rect 43652 39900 44156 39956
rect 44212 39900 44222 39956
rect 6850 39788 6860 39844
rect 6916 39788 7756 39844
rect 7812 39788 7822 39844
rect 16258 39788 16268 39844
rect 16324 39788 16940 39844
rect 16996 39788 17006 39844
rect 22418 39788 22428 39844
rect 22484 39788 44380 39844
rect 44436 39788 44446 39844
rect 3154 39676 3164 39732
rect 3220 39676 10724 39732
rect 11218 39676 11228 39732
rect 11284 39676 11900 39732
rect 11956 39676 11966 39732
rect 20962 39676 20972 39732
rect 21028 39676 26908 39732
rect 30706 39676 30716 39732
rect 30772 39676 31500 39732
rect 31556 39676 31566 39732
rect 35074 39676 35084 39732
rect 35140 39676 35980 39732
rect 36036 39676 36046 39732
rect 10668 39620 10724 39676
rect 7410 39564 7420 39620
rect 7476 39564 8092 39620
rect 8148 39564 8158 39620
rect 10668 39564 13468 39620
rect 13524 39564 13534 39620
rect 23202 39564 23212 39620
rect 23268 39564 23548 39620
rect 23604 39564 24444 39620
rect 24500 39564 24510 39620
rect 3378 39452 3388 39508
rect 3444 39452 4284 39508
rect 4340 39452 4350 39508
rect 7746 39452 7756 39508
rect 7812 39452 7980 39508
rect 8036 39452 8046 39508
rect 8194 39452 8204 39508
rect 8260 39452 8988 39508
rect 9044 39452 9054 39508
rect 26852 39396 26908 39676
rect 32610 39564 32620 39620
rect 32676 39564 33516 39620
rect 33572 39564 33582 39620
rect 39554 39564 39564 39620
rect 39620 39564 40236 39620
rect 40292 39564 40302 39620
rect 41122 39564 41132 39620
rect 41188 39564 41580 39620
rect 41636 39564 41646 39620
rect 41906 39564 41916 39620
rect 41972 39564 42476 39620
rect 42532 39564 43036 39620
rect 43092 39564 43102 39620
rect 44146 39564 44156 39620
rect 44212 39564 44492 39620
rect 44548 39564 44558 39620
rect 41580 39508 41636 39564
rect 39330 39452 39340 39508
rect 39396 39452 39676 39508
rect 39732 39452 41244 39508
rect 41300 39452 41310 39508
rect 41580 39452 42252 39508
rect 42308 39452 42318 39508
rect 7046 39340 7084 39396
rect 7140 39340 7150 39396
rect 8082 39340 8092 39396
rect 8148 39340 8540 39396
rect 8596 39340 11116 39396
rect 11172 39340 11182 39396
rect 26852 39340 45836 39396
rect 45892 39340 45902 39396
rect 1810 39228 1820 39284
rect 1876 39228 2604 39284
rect 2660 39228 3388 39284
rect 32386 39228 32396 39284
rect 32452 39228 34412 39284
rect 34468 39228 34478 39284
rect 34626 39228 34636 39284
rect 34692 39228 35084 39284
rect 35140 39228 35150 39284
rect 3332 39172 3388 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 3332 39116 12124 39172
rect 12180 39116 12348 39172
rect 12404 39116 12414 39172
rect 24770 39116 24780 39172
rect 24836 39116 25788 39172
rect 25844 39116 25854 39172
rect 35858 39116 35868 39172
rect 35924 39116 36428 39172
rect 36484 39116 36494 39172
rect 3938 39004 3948 39060
rect 4004 39004 4620 39060
rect 4676 39004 4686 39060
rect 14690 39004 14700 39060
rect 14756 39004 16492 39060
rect 16548 39004 16558 39060
rect 20626 39004 20636 39060
rect 20692 39004 21308 39060
rect 21364 39004 22316 39060
rect 22372 39004 22382 39060
rect 40786 39004 40796 39060
rect 40852 39004 41804 39060
rect 41860 39004 41870 39060
rect 3378 38892 3388 38948
rect 3444 38892 4844 38948
rect 4900 38892 5404 38948
rect 5460 38892 7196 38948
rect 7252 38892 7262 38948
rect 8054 38892 8092 38948
rect 8148 38892 8158 38948
rect 13458 38892 13468 38948
rect 13524 38892 15484 38948
rect 15540 38892 15550 38948
rect 24322 38892 24332 38948
rect 24388 38892 24668 38948
rect 24724 38892 25788 38948
rect 25844 38892 25854 38948
rect 26226 38892 26236 38948
rect 26292 38892 26796 38948
rect 26852 38892 26862 38948
rect 29586 38892 29596 38948
rect 29652 38892 30940 38948
rect 30996 38892 31724 38948
rect 31780 38892 31790 38948
rect 34178 38892 34188 38948
rect 34244 38892 34972 38948
rect 35028 38892 39340 38948
rect 39396 38892 39406 38948
rect 41010 38892 41020 38948
rect 41076 38892 41692 38948
rect 41748 38892 41758 38948
rect 43698 38892 43708 38948
rect 43764 38892 44044 38948
rect 44100 38892 44110 38948
rect 7270 38780 7308 38836
rect 7364 38780 7374 38836
rect 7942 38780 7980 38836
rect 8036 38780 8046 38836
rect 8306 38780 8316 38836
rect 8372 38780 8988 38836
rect 9044 38780 9054 38836
rect 15810 38780 15820 38836
rect 15876 38780 15886 38836
rect 22754 38780 22764 38836
rect 22820 38780 23548 38836
rect 23604 38780 23614 38836
rect 25666 38780 25676 38836
rect 25732 38780 26460 38836
rect 26516 38780 26526 38836
rect 34738 38780 34748 38836
rect 34804 38780 35196 38836
rect 35252 38780 37324 38836
rect 37380 38780 37390 38836
rect 37986 38780 37996 38836
rect 38052 38780 38668 38836
rect 38724 38780 40460 38836
rect 40516 38780 40526 38836
rect 15820 38724 15876 38780
rect 1586 38668 1596 38724
rect 1652 38668 2156 38724
rect 2212 38668 2222 38724
rect 7756 38668 7868 38724
rect 7924 38668 7934 38724
rect 15820 38668 16268 38724
rect 16324 38668 24556 38724
rect 24612 38668 24622 38724
rect 35858 38668 35868 38724
rect 35924 38668 36092 38724
rect 36148 38668 36158 38724
rect 48178 38668 48188 38724
rect 48244 38668 48254 38724
rect 0 38612 800 38640
rect 0 38556 1708 38612
rect 1764 38556 1774 38612
rect 3612 38556 4284 38612
rect 4340 38556 4350 38612
rect 0 38528 800 38556
rect 3612 38500 3668 38556
rect 7756 38500 7812 38668
rect 48188 38612 48244 38668
rect 49200 38612 50000 38640
rect 13794 38556 13804 38612
rect 13860 38556 14924 38612
rect 14980 38556 14990 38612
rect 18610 38556 18620 38612
rect 18676 38556 42364 38612
rect 42420 38556 42430 38612
rect 48188 38556 50000 38612
rect 49200 38528 50000 38556
rect 3602 38444 3612 38500
rect 3668 38444 3678 38500
rect 7634 38444 7644 38500
rect 7700 38444 7812 38500
rect 18834 38444 18844 38500
rect 18900 38444 19516 38500
rect 19572 38444 19582 38500
rect 20290 38444 20300 38500
rect 20356 38444 28700 38500
rect 28756 38444 28766 38500
rect 36054 38444 36092 38500
rect 36148 38444 36158 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 8054 38332 8092 38388
rect 8148 38332 8158 38388
rect 23986 38332 23996 38388
rect 24052 38332 24892 38388
rect 24948 38332 24958 38388
rect 28998 38332 29036 38388
rect 29092 38332 29102 38388
rect 8166 38220 8204 38276
rect 8260 38220 8270 38276
rect 20738 38220 20748 38276
rect 20804 38220 28588 38276
rect 28644 38220 28654 38276
rect 28914 38220 28924 38276
rect 28980 38220 29260 38276
rect 29316 38220 29326 38276
rect 2930 38108 2940 38164
rect 2996 38108 8876 38164
rect 8932 38108 9436 38164
rect 9492 38108 9502 38164
rect 28466 38108 28476 38164
rect 28532 38108 31276 38164
rect 31332 38108 31342 38164
rect 24658 37996 24668 38052
rect 24724 37996 25004 38052
rect 25060 37996 26124 38052
rect 26180 37996 26190 38052
rect 27458 37996 27468 38052
rect 27524 37996 28812 38052
rect 28868 37996 28878 38052
rect 29586 37996 29596 38052
rect 29652 37996 30044 38052
rect 30100 37996 30110 38052
rect 38770 37996 38780 38052
rect 38836 37996 39564 38052
rect 39620 37996 39900 38052
rect 39956 37996 39966 38052
rect 29138 37884 29148 37940
rect 29204 37884 29932 37940
rect 29988 37884 29998 37940
rect 3910 37772 3948 37828
rect 4004 37772 4014 37828
rect 24882 37772 24892 37828
rect 24948 37772 25564 37828
rect 25620 37772 25630 37828
rect 29586 37772 29596 37828
rect 29652 37772 30492 37828
rect 30548 37772 30558 37828
rect 7634 37660 7644 37716
rect 7700 37660 7710 37716
rect 2034 37436 2044 37492
rect 2100 37436 3388 37492
rect 3332 37268 3388 37436
rect 7644 37268 7700 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 27794 37548 27804 37604
rect 27860 37548 28252 37604
rect 28308 37548 28318 37604
rect 46050 37548 46060 37604
rect 46116 37548 46844 37604
rect 46900 37548 46910 37604
rect 18050 37436 18060 37492
rect 18116 37436 18508 37492
rect 18564 37436 18574 37492
rect 26562 37436 26572 37492
rect 26628 37436 27244 37492
rect 27300 37436 27310 37492
rect 9426 37324 9436 37380
rect 9492 37324 11564 37380
rect 11620 37324 11630 37380
rect 16258 37324 16268 37380
rect 16324 37324 19068 37380
rect 19124 37324 19404 37380
rect 19460 37324 19516 37380
rect 19572 37324 19582 37380
rect 22642 37324 22652 37380
rect 22708 37324 26684 37380
rect 26740 37324 27020 37380
rect 27076 37324 27086 37380
rect 34738 37324 34748 37380
rect 34804 37324 34972 37380
rect 35028 37324 35038 37380
rect 37538 37324 37548 37380
rect 37604 37324 38108 37380
rect 38164 37324 39788 37380
rect 39844 37324 39854 37380
rect 44258 37324 44268 37380
rect 44324 37324 44828 37380
rect 44884 37324 44894 37380
rect 3332 37212 4396 37268
rect 4452 37212 7644 37268
rect 7700 37212 7710 37268
rect 8194 37212 8204 37268
rect 8260 37212 9548 37268
rect 9604 37212 9614 37268
rect 19842 37212 19852 37268
rect 19908 37212 20300 37268
rect 20356 37212 20366 37268
rect 28018 37212 28028 37268
rect 28084 37212 28094 37268
rect 28578 37212 28588 37268
rect 28644 37212 29596 37268
rect 29652 37212 29662 37268
rect 30818 37212 30828 37268
rect 30884 37212 34748 37268
rect 34804 37212 41132 37268
rect 41188 37212 41804 37268
rect 41860 37212 41870 37268
rect 42130 37212 42140 37268
rect 42196 37212 43036 37268
rect 43092 37212 43484 37268
rect 43540 37212 43550 37268
rect 46050 37212 46060 37268
rect 46116 37212 46844 37268
rect 46900 37212 46910 37268
rect 28028 37156 28084 37212
rect 6514 37100 6524 37156
rect 6580 37100 7532 37156
rect 7588 37100 8316 37156
rect 8372 37100 8382 37156
rect 14242 37100 14252 37156
rect 14308 37100 15036 37156
rect 15092 37100 15372 37156
rect 15428 37100 15438 37156
rect 26114 37100 26124 37156
rect 26180 37100 27356 37156
rect 27412 37100 28084 37156
rect 28354 37100 28364 37156
rect 28420 37100 29260 37156
rect 29316 37100 29484 37156
rect 29540 37100 29550 37156
rect 31042 37100 31052 37156
rect 31108 37100 31948 37156
rect 32004 37100 32014 37156
rect 6636 36988 14588 37044
rect 14644 36988 14654 37044
rect 19954 36988 19964 37044
rect 20020 36988 20860 37044
rect 20916 36988 21868 37044
rect 21924 36988 21934 37044
rect 26562 36988 26572 37044
rect 26628 36988 26684 37044
rect 26740 36988 26750 37044
rect 30146 36988 30156 37044
rect 30212 36988 31500 37044
rect 31556 36988 32060 37044
rect 32116 36988 32620 37044
rect 32676 36988 32686 37044
rect 45938 36988 45948 37044
rect 46004 36988 47852 37044
rect 47908 36988 47918 37044
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 1362 36652 1372 36708
rect 1428 36652 4396 36708
rect 4452 36652 4462 36708
rect 6636 36596 6692 36988
rect 16706 36876 16716 36932
rect 16772 36876 26348 36932
rect 26404 36876 26414 36932
rect 30034 36876 30044 36932
rect 30100 36876 31276 36932
rect 31332 36876 31836 36932
rect 31892 36876 31902 36932
rect 36418 36876 36428 36932
rect 36484 36876 40236 36932
rect 40292 36876 40302 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 17826 36764 17836 36820
rect 17892 36764 23884 36820
rect 23940 36764 23950 36820
rect 40114 36764 40124 36820
rect 40180 36764 41132 36820
rect 41188 36764 41198 36820
rect 6850 36652 6860 36708
rect 6916 36652 22652 36708
rect 22708 36652 23996 36708
rect 24052 36652 24062 36708
rect 30146 36652 30156 36708
rect 30212 36652 37884 36708
rect 37940 36652 37950 36708
rect 2258 36540 2268 36596
rect 2324 36540 6692 36596
rect 7970 36540 7980 36596
rect 8036 36540 8764 36596
rect 8820 36540 8830 36596
rect 11554 36540 11564 36596
rect 11620 36540 12572 36596
rect 12628 36540 12638 36596
rect 22278 36540 22316 36596
rect 22372 36540 22382 36596
rect 23090 36540 23100 36596
rect 23156 36540 23772 36596
rect 23828 36540 23838 36596
rect 32946 36540 32956 36596
rect 33012 36540 43596 36596
rect 43652 36540 43662 36596
rect 22316 36484 22372 36540
rect 1586 36428 1596 36484
rect 1652 36428 12012 36484
rect 12068 36428 12078 36484
rect 19282 36428 19292 36484
rect 19348 36428 19740 36484
rect 19796 36428 21420 36484
rect 21476 36428 21486 36484
rect 22316 36428 25676 36484
rect 25732 36428 25742 36484
rect 27346 36428 27356 36484
rect 27412 36428 27804 36484
rect 27860 36428 27870 36484
rect 38322 36428 38332 36484
rect 38388 36428 39452 36484
rect 39508 36428 39518 36484
rect 41206 36428 41244 36484
rect 41300 36428 41692 36484
rect 41748 36428 41758 36484
rect 45602 36428 45612 36484
rect 45668 36428 46172 36484
rect 46228 36428 46620 36484
rect 46676 36428 46686 36484
rect 3826 36316 3836 36372
rect 3892 36316 5068 36372
rect 5124 36316 6860 36372
rect 6916 36316 6926 36372
rect 19394 36316 19404 36372
rect 19460 36316 19852 36372
rect 19908 36316 19918 36372
rect 23426 36316 23436 36372
rect 23492 36316 28700 36372
rect 28756 36316 28766 36372
rect 37874 36316 37884 36372
rect 37940 36316 39116 36372
rect 39172 36316 39900 36372
rect 39956 36316 39966 36372
rect 5170 36204 5180 36260
rect 5236 36204 6076 36260
rect 6132 36204 6142 36260
rect 18274 36204 18284 36260
rect 18340 36204 19180 36260
rect 19236 36204 19246 36260
rect 39218 36204 39228 36260
rect 39284 36204 39788 36260
rect 39844 36204 39854 36260
rect 0 36148 800 36176
rect 49200 36148 50000 36176
rect 0 36092 1708 36148
rect 1764 36092 1774 36148
rect 39890 36092 39900 36148
rect 39956 36092 40348 36148
rect 40404 36092 40414 36148
rect 48178 36092 48188 36148
rect 48244 36092 50000 36148
rect 0 36064 800 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 49200 36064 50000 36092
rect 9538 35980 9548 36036
rect 9604 35980 11788 36036
rect 11844 35980 19684 36036
rect 24210 35980 24220 36036
rect 24276 35980 24556 36036
rect 24612 35980 24622 36036
rect 19628 35924 19684 35980
rect 17490 35868 17500 35924
rect 17556 35868 17566 35924
rect 18806 35868 18844 35924
rect 18900 35868 18910 35924
rect 19628 35868 20972 35924
rect 21028 35868 22764 35924
rect 22820 35868 22830 35924
rect 17500 35700 17556 35868
rect 17938 35756 17948 35812
rect 18004 35756 19292 35812
rect 19348 35756 19358 35812
rect 19730 35756 19740 35812
rect 19796 35756 20412 35812
rect 20468 35756 20478 35812
rect 28466 35756 28476 35812
rect 28532 35756 29932 35812
rect 29988 35756 29998 35812
rect 33282 35756 33292 35812
rect 33348 35756 34412 35812
rect 34468 35756 35532 35812
rect 35588 35756 35598 35812
rect 41122 35756 41132 35812
rect 41188 35756 42364 35812
rect 42420 35756 42430 35812
rect 17500 35644 17724 35700
rect 17780 35644 17790 35700
rect 21634 35644 21644 35700
rect 21700 35644 23548 35700
rect 23604 35644 23614 35700
rect 23874 35644 23884 35700
rect 23940 35644 26908 35700
rect 26964 35644 27804 35700
rect 27860 35644 27870 35700
rect 29474 35644 29484 35700
rect 29540 35644 30044 35700
rect 30100 35644 30716 35700
rect 30772 35644 30782 35700
rect 32722 35644 32732 35700
rect 32788 35644 34860 35700
rect 34916 35644 38444 35700
rect 38500 35644 38510 35700
rect 38612 35644 39004 35700
rect 39060 35644 39070 35700
rect 39778 35644 39788 35700
rect 39844 35644 40236 35700
rect 40292 35644 40572 35700
rect 40628 35644 40638 35700
rect 38612 35588 38668 35644
rect 2258 35532 2268 35588
rect 2324 35532 4956 35588
rect 5012 35532 5022 35588
rect 17826 35532 17836 35588
rect 17892 35532 19068 35588
rect 19124 35532 19134 35588
rect 20626 35532 20636 35588
rect 20692 35532 21308 35588
rect 21364 35532 21374 35588
rect 24210 35532 24220 35588
rect 24276 35532 26796 35588
rect 26852 35532 26862 35588
rect 37762 35532 37772 35588
rect 37828 35532 38668 35588
rect 45602 35532 45612 35588
rect 45668 35532 46172 35588
rect 46228 35532 46238 35588
rect 18386 35420 18396 35476
rect 18452 35420 19404 35476
rect 19460 35420 19470 35476
rect 21410 35420 21420 35476
rect 21476 35420 21756 35476
rect 21812 35420 21822 35476
rect 26226 35420 26236 35476
rect 26292 35420 26908 35476
rect 30006 35420 30044 35476
rect 30100 35420 30110 35476
rect 37426 35420 37436 35476
rect 37492 35420 38108 35476
rect 38164 35420 39004 35476
rect 39060 35420 39070 35476
rect 41682 35420 41692 35476
rect 41748 35420 43148 35476
rect 43204 35420 43214 35476
rect 26852 35364 26908 35420
rect 4946 35308 4956 35364
rect 5012 35308 5628 35364
rect 5684 35308 5694 35364
rect 8876 35308 8988 35364
rect 9044 35308 9054 35364
rect 17042 35308 17052 35364
rect 17108 35308 19180 35364
rect 19236 35308 19246 35364
rect 20402 35308 20412 35364
rect 20468 35308 21196 35364
rect 21252 35308 21262 35364
rect 22082 35308 22092 35364
rect 22148 35308 23100 35364
rect 23156 35308 26572 35364
rect 26628 35308 26638 35364
rect 26852 35308 27356 35364
rect 27412 35308 28252 35364
rect 28308 35308 28318 35364
rect 29670 35308 29708 35364
rect 29764 35308 29774 35364
rect 30156 35308 34972 35364
rect 35028 35308 35038 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 8866 35252 8876 35308
rect 8932 35252 8942 35308
rect 30156 35252 30212 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 6850 35196 6860 35252
rect 6916 35196 7420 35252
rect 7476 35196 7486 35252
rect 24546 35196 24556 35252
rect 24612 35196 30212 35252
rect 30930 35196 30940 35252
rect 30996 35196 32060 35252
rect 32116 35196 32126 35252
rect 38546 35196 38556 35252
rect 38612 35196 39340 35252
rect 39396 35196 39406 35252
rect 29922 35084 29932 35140
rect 29988 35084 30492 35140
rect 30548 35084 31836 35140
rect 31892 35084 31902 35140
rect 35252 35084 41692 35140
rect 41748 35084 41758 35140
rect 35252 35028 35308 35084
rect 3714 34972 3724 35028
rect 3780 34972 4060 35028
rect 4116 34972 4126 35028
rect 5058 34972 5068 35028
rect 5124 34972 7644 35028
rect 7700 34972 7710 35028
rect 16706 34972 16716 35028
rect 16772 34972 17836 35028
rect 17892 34972 17902 35028
rect 27122 34972 27132 35028
rect 27188 34972 27692 35028
rect 27748 34972 27758 35028
rect 29026 34972 29036 35028
rect 29092 34972 35308 35028
rect 4274 34860 4284 34916
rect 4340 34860 5964 34916
rect 6020 34860 6972 34916
rect 7028 34860 7038 34916
rect 16034 34860 16044 34916
rect 16100 34860 17948 34916
rect 18004 34860 18014 34916
rect 18610 34860 18620 34916
rect 18676 34860 18956 34916
rect 19012 34860 19022 34916
rect 21970 34860 21980 34916
rect 22036 34860 22988 34916
rect 23044 34860 25900 34916
rect 25956 34860 25966 34916
rect 31042 34860 31052 34916
rect 31108 34860 31836 34916
rect 31892 34860 31902 34916
rect 34178 34860 34188 34916
rect 34244 34860 35196 34916
rect 35252 34860 35262 34916
rect 37762 34860 37772 34916
rect 37828 34860 38332 34916
rect 38388 34860 38398 34916
rect 41234 34860 41244 34916
rect 41300 34860 42476 34916
rect 42532 34860 42542 34916
rect 4386 34748 4396 34804
rect 4452 34748 6748 34804
rect 6804 34748 7756 34804
rect 7812 34748 7822 34804
rect 15922 34748 15932 34804
rect 15988 34748 20188 34804
rect 20244 34748 21308 34804
rect 21364 34748 21868 34804
rect 21924 34748 21934 34804
rect 27010 34748 27020 34804
rect 27076 34748 28364 34804
rect 28420 34748 29484 34804
rect 29540 34748 29820 34804
rect 29876 34748 38668 34804
rect 39666 34748 39676 34804
rect 39732 34748 40908 34804
rect 40964 34748 40974 34804
rect 5730 34636 5740 34692
rect 5796 34636 7420 34692
rect 7476 34636 7532 34692
rect 7588 34636 7598 34692
rect 12450 34636 12460 34692
rect 12516 34636 17388 34692
rect 17444 34636 18508 34692
rect 18564 34636 18574 34692
rect 34738 34636 34748 34692
rect 34804 34636 36204 34692
rect 36260 34636 37100 34692
rect 37156 34636 37166 34692
rect 6178 34524 6188 34580
rect 6244 34524 9772 34580
rect 9828 34524 9838 34580
rect 27906 34524 27916 34580
rect 27972 34524 28476 34580
rect 28532 34524 29036 34580
rect 29092 34524 29260 34580
rect 29316 34524 35812 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 34636 34412 35532 34468
rect 35588 34412 35598 34468
rect 3602 34300 3612 34356
rect 3668 34300 4620 34356
rect 4676 34300 5068 34356
rect 5124 34300 6188 34356
rect 6244 34300 6254 34356
rect 7970 34300 7980 34356
rect 8036 34300 8540 34356
rect 8596 34300 9100 34356
rect 9156 34300 9324 34356
rect 9380 34300 9390 34356
rect 14354 34300 14364 34356
rect 14420 34300 14700 34356
rect 14756 34300 14766 34356
rect 17714 34300 17724 34356
rect 17780 34300 18620 34356
rect 18676 34300 18686 34356
rect 21410 34300 21420 34356
rect 21476 34300 22204 34356
rect 22260 34300 22270 34356
rect 24882 34300 24892 34356
rect 24948 34300 26460 34356
rect 26516 34300 26526 34356
rect 34636 34244 34692 34412
rect 35756 34356 35812 34524
rect 38612 34468 38668 34748
rect 46246 34524 46284 34580
rect 46340 34524 46350 34580
rect 38612 34412 46620 34468
rect 46676 34412 47740 34468
rect 47796 34412 47806 34468
rect 35298 34300 35308 34356
rect 35364 34300 35374 34356
rect 35756 34300 47068 34356
rect 47124 34300 47134 34356
rect 4274 34188 4284 34244
rect 4340 34188 5180 34244
rect 5236 34188 6412 34244
rect 6468 34188 6478 34244
rect 12674 34188 12684 34244
rect 12740 34188 13916 34244
rect 13972 34188 16492 34244
rect 16548 34188 16558 34244
rect 18834 34188 18844 34244
rect 18900 34188 18910 34244
rect 33730 34188 33740 34244
rect 33796 34188 34636 34244
rect 34692 34188 34702 34244
rect 2258 34076 2268 34132
rect 2324 34076 12236 34132
rect 12292 34076 12302 34132
rect 14354 34076 14364 34132
rect 14420 34076 16268 34132
rect 16324 34076 16334 34132
rect 2678 33964 2716 34020
rect 2772 33964 2782 34020
rect 3332 33908 3388 34020
rect 3444 33964 3836 34020
rect 3892 33964 4732 34020
rect 4788 33964 15148 34020
rect 15810 33964 15820 34020
rect 15876 33964 16380 34020
rect 16436 33964 16446 34020
rect 15092 33908 15148 33964
rect 18844 33908 18900 34188
rect 19954 34076 19964 34132
rect 20020 34076 25452 34132
rect 25508 34076 25518 34132
rect 35308 34020 35364 34300
rect 35522 34188 35532 34244
rect 35588 34188 35868 34244
rect 35924 34188 40348 34244
rect 40404 34188 40414 34244
rect 45042 34188 45052 34244
rect 45108 34188 45724 34244
rect 45780 34188 45790 34244
rect 46470 34076 46508 34132
rect 46564 34076 46574 34132
rect 19282 33964 19292 34020
rect 19348 33964 21084 34020
rect 21140 33964 30156 34020
rect 30212 33964 30222 34020
rect 34402 33964 34412 34020
rect 34468 33964 35364 34020
rect 38994 33964 39004 34020
rect 39060 33964 39676 34020
rect 39732 33964 39742 34020
rect 2146 33852 2156 33908
rect 2212 33852 2940 33908
rect 2996 33852 3388 33908
rect 6514 33852 6524 33908
rect 6580 33852 8428 33908
rect 8484 33852 8494 33908
rect 15092 33852 18900 33908
rect 25890 33852 25900 33908
rect 25956 33852 25966 33908
rect 34850 33852 34860 33908
rect 34916 33852 35756 33908
rect 35812 33852 35822 33908
rect 40450 33852 40460 33908
rect 40516 33852 40908 33908
rect 40964 33852 40974 33908
rect 46610 33852 46620 33908
rect 46676 33852 47292 33908
rect 47348 33852 47358 33908
rect 14914 33740 14924 33796
rect 14980 33740 17388 33796
rect 17444 33740 17454 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 25900 33684 25956 33852
rect 47058 33740 47068 33796
rect 47124 33740 47628 33796
rect 47684 33740 48300 33796
rect 48356 33740 48366 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 49200 33684 50000 33712
rect 0 33628 1708 33684
rect 1764 33628 1876 33684
rect 2034 33628 2044 33684
rect 2100 33628 2110 33684
rect 14130 33628 14140 33684
rect 14196 33628 16828 33684
rect 16884 33628 16894 33684
rect 18694 33628 18732 33684
rect 18788 33628 18798 33684
rect 25900 33628 31052 33684
rect 31108 33628 31118 33684
rect 37538 33628 37548 33684
rect 37604 33628 38332 33684
rect 38388 33628 38398 33684
rect 41234 33628 41244 33684
rect 41300 33628 42028 33684
rect 42084 33628 42924 33684
rect 42980 33628 42990 33684
rect 48178 33628 48188 33684
rect 48244 33628 50000 33684
rect 0 33600 800 33628
rect 1820 33124 1876 33628
rect 2044 33572 2100 33628
rect 49200 33600 50000 33628
rect 2044 33516 2380 33572
rect 2436 33516 3388 33572
rect 3444 33516 3454 33572
rect 6962 33516 6972 33572
rect 7028 33516 10332 33572
rect 10388 33516 10398 33572
rect 14018 33516 14028 33572
rect 14084 33516 14700 33572
rect 14756 33516 14766 33572
rect 18162 33516 18172 33572
rect 18228 33516 19068 33572
rect 19124 33516 19628 33572
rect 19684 33516 19694 33572
rect 4274 33404 4284 33460
rect 4340 33404 6300 33460
rect 6356 33404 6366 33460
rect 8642 33404 8652 33460
rect 8708 33404 12572 33460
rect 12628 33404 14476 33460
rect 14532 33404 15484 33460
rect 15540 33404 15550 33460
rect 37090 33404 37100 33460
rect 37156 33404 37884 33460
rect 37940 33404 37950 33460
rect 8082 33292 8092 33348
rect 8148 33292 9548 33348
rect 9604 33292 9614 33348
rect 11890 33292 11900 33348
rect 11956 33292 12236 33348
rect 12292 33292 12684 33348
rect 12740 33292 13132 33348
rect 13188 33292 13198 33348
rect 18498 33292 18508 33348
rect 18564 33292 18732 33348
rect 18788 33292 21308 33348
rect 21364 33292 21374 33348
rect 42690 33292 42700 33348
rect 42756 33292 43596 33348
rect 43652 33292 43662 33348
rect 46162 33292 46172 33348
rect 46228 33292 46508 33348
rect 46564 33292 46574 33348
rect 4834 33180 4844 33236
rect 4900 33180 5740 33236
rect 5796 33180 5806 33236
rect 8194 33180 8204 33236
rect 8260 33180 9324 33236
rect 9380 33180 9996 33236
rect 10052 33180 10062 33236
rect 10322 33180 10332 33236
rect 10388 33180 13580 33236
rect 13636 33180 13646 33236
rect 14802 33180 14812 33236
rect 14868 33180 16044 33236
rect 16100 33180 16110 33236
rect 19618 33180 19628 33236
rect 19684 33180 20524 33236
rect 20580 33180 21532 33236
rect 21588 33180 21598 33236
rect 21942 33180 21980 33236
rect 22036 33180 22046 33236
rect 39778 33180 39788 33236
rect 39844 33180 41132 33236
rect 41188 33180 41198 33236
rect 1820 33068 1932 33124
rect 1988 33068 1998 33124
rect 9538 33068 9548 33124
rect 9604 33068 10220 33124
rect 10276 33068 10286 33124
rect 10658 33068 10668 33124
rect 10724 33068 11676 33124
rect 11732 33068 12124 33124
rect 12180 33068 12190 33124
rect 17826 33068 17836 33124
rect 17892 33068 17948 33124
rect 18004 33068 18396 33124
rect 18452 33068 18462 33124
rect 19394 33068 19404 33124
rect 19460 33068 19852 33124
rect 19908 33068 19918 33124
rect 20290 33068 20300 33124
rect 20356 33068 21308 33124
rect 21364 33068 21374 33124
rect 32050 33068 32060 33124
rect 32116 33068 37212 33124
rect 37268 33068 37278 33124
rect 39554 33068 39564 33124
rect 39620 33068 40124 33124
rect 40180 33068 40190 33124
rect 41346 33068 41356 33124
rect 41412 33068 42476 33124
rect 42532 33068 42542 33124
rect 41682 32956 41692 33012
rect 41748 32956 43036 33012
rect 43092 32956 43102 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 7410 32844 7420 32900
rect 7476 32844 7644 32900
rect 7700 32844 8652 32900
rect 8708 32844 8718 32900
rect 23314 32844 23324 32900
rect 23380 32844 38668 32900
rect 39778 32844 39788 32900
rect 39844 32844 40012 32900
rect 40068 32844 44044 32900
rect 44100 32844 44110 32900
rect 38612 32788 38668 32844
rect 2482 32732 2492 32788
rect 2548 32732 2828 32788
rect 2884 32732 3388 32788
rect 3444 32732 4284 32788
rect 4340 32732 4350 32788
rect 7746 32732 7756 32788
rect 7812 32732 8092 32788
rect 8148 32732 10108 32788
rect 10164 32732 10174 32788
rect 22082 32732 22092 32788
rect 22148 32732 28252 32788
rect 28308 32732 28318 32788
rect 34178 32732 34188 32788
rect 34244 32732 34972 32788
rect 35028 32732 35038 32788
rect 38612 32732 40460 32788
rect 40516 32732 40526 32788
rect 40898 32732 40908 32788
rect 40964 32732 41692 32788
rect 41748 32732 41758 32788
rect 6290 32620 6300 32676
rect 6356 32620 8428 32676
rect 8484 32620 9548 32676
rect 9604 32620 9614 32676
rect 10994 32620 11004 32676
rect 11060 32620 11452 32676
rect 11508 32620 11518 32676
rect 19954 32620 19964 32676
rect 20020 32620 20412 32676
rect 20468 32620 20972 32676
rect 21028 32620 21038 32676
rect 36530 32620 36540 32676
rect 36596 32620 37212 32676
rect 37268 32620 37278 32676
rect 40338 32620 40348 32676
rect 40404 32620 41244 32676
rect 41300 32620 41310 32676
rect 46050 32620 46060 32676
rect 46116 32620 46732 32676
rect 46788 32620 46798 32676
rect 2930 32508 2940 32564
rect 2996 32508 3836 32564
rect 3892 32508 3902 32564
rect 6066 32508 6076 32564
rect 6132 32508 6142 32564
rect 7196 32508 7980 32564
rect 8036 32508 8046 32564
rect 9650 32508 9660 32564
rect 9716 32508 10668 32564
rect 10724 32508 10734 32564
rect 12338 32508 12348 32564
rect 12404 32508 12572 32564
rect 12628 32508 12638 32564
rect 20738 32508 20748 32564
rect 20804 32508 21868 32564
rect 21924 32508 22764 32564
rect 22820 32508 22830 32564
rect 29250 32508 29260 32564
rect 29316 32508 31052 32564
rect 31108 32508 32060 32564
rect 32116 32508 32126 32564
rect 34710 32508 34748 32564
rect 34804 32508 34814 32564
rect 36418 32508 36428 32564
rect 36484 32508 37436 32564
rect 37492 32508 38556 32564
rect 38612 32508 38622 32564
rect 6076 32452 6132 32508
rect 7196 32452 7252 32508
rect 3332 32396 6132 32452
rect 6514 32396 6524 32452
rect 6580 32396 7196 32452
rect 7252 32396 7262 32452
rect 7634 32396 7644 32452
rect 7700 32396 24668 32452
rect 24724 32396 25228 32452
rect 25284 32396 25294 32452
rect 3332 32340 3388 32396
rect 2034 32284 2044 32340
rect 2100 32284 3388 32340
rect 5954 32284 5964 32340
rect 6020 32284 8540 32340
rect 8596 32284 8606 32340
rect 10210 32284 10220 32340
rect 10276 32284 11228 32340
rect 11284 32284 11294 32340
rect 17042 32284 17052 32340
rect 17108 32284 18956 32340
rect 19012 32284 23996 32340
rect 24052 32284 24062 32340
rect 27458 32284 27468 32340
rect 27524 32284 36876 32340
rect 36932 32284 36942 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 2678 32060 2716 32116
rect 2772 32060 2782 32116
rect 14242 32060 14252 32116
rect 14308 32060 14588 32116
rect 14644 32060 14654 32116
rect 3826 31948 3836 32004
rect 3892 31948 6748 32004
rect 6804 31948 6814 32004
rect 9986 31948 9996 32004
rect 10052 31948 10892 32004
rect 10948 31948 11116 32004
rect 11172 31948 11182 32004
rect 12338 31948 12348 32004
rect 12404 31948 13356 32004
rect 13412 31948 14700 32004
rect 14756 31948 14766 32004
rect 31500 31948 32004 32004
rect 31500 31892 31556 31948
rect 31948 31892 32004 31948
rect 6850 31836 6860 31892
rect 6916 31836 7532 31892
rect 7588 31836 9100 31892
rect 9156 31836 9166 31892
rect 15698 31836 15708 31892
rect 15764 31836 16156 31892
rect 16212 31836 16222 31892
rect 23314 31836 23324 31892
rect 23380 31836 31556 31892
rect 31686 31836 31724 31892
rect 31780 31836 31790 31892
rect 31948 31836 32956 31892
rect 33012 31836 33022 31892
rect 34402 31836 34412 31892
rect 34468 31836 35644 31892
rect 35700 31836 35710 31892
rect 41346 31836 41356 31892
rect 41412 31836 41916 31892
rect 41972 31836 41982 31892
rect 42578 31836 42588 31892
rect 42644 31836 43708 31892
rect 43764 31836 43774 31892
rect 46274 31836 46284 31892
rect 46340 31836 47516 31892
rect 47572 31836 47582 31892
rect 7074 31724 7084 31780
rect 7140 31724 8092 31780
rect 8148 31724 8158 31780
rect 8316 31724 13468 31780
rect 13524 31724 13534 31780
rect 14914 31724 14924 31780
rect 14980 31724 15372 31780
rect 15428 31724 15438 31780
rect 22530 31724 22540 31780
rect 22596 31724 23548 31780
rect 23604 31724 23614 31780
rect 29922 31724 29932 31780
rect 29988 31724 30716 31780
rect 30772 31724 31612 31780
rect 31668 31724 31678 31780
rect 34514 31724 34524 31780
rect 34580 31724 35532 31780
rect 35588 31724 35598 31780
rect 8316 31668 8372 31724
rect 1922 31612 1932 31668
rect 1988 31612 2492 31668
rect 2548 31612 3388 31668
rect 3826 31612 3836 31668
rect 3892 31612 8372 31668
rect 9538 31612 9548 31668
rect 9604 31612 11116 31668
rect 11172 31612 11182 31668
rect 12786 31612 12796 31668
rect 12852 31612 14700 31668
rect 14756 31612 27020 31668
rect 27076 31612 27244 31668
rect 27300 31612 27468 31668
rect 27524 31612 27534 31668
rect 28578 31612 28588 31668
rect 28644 31612 29484 31668
rect 29540 31612 29550 31668
rect 34626 31612 34636 31668
rect 34692 31612 35980 31668
rect 36036 31612 37436 31668
rect 37492 31612 37502 31668
rect 38770 31612 38780 31668
rect 38836 31612 39788 31668
rect 39844 31612 39854 31668
rect 3332 31556 3388 31612
rect 3332 31500 6076 31556
rect 6132 31500 7420 31556
rect 7476 31500 7486 31556
rect 8642 31500 8652 31556
rect 8708 31500 8876 31556
rect 8932 31500 9996 31556
rect 10052 31500 10062 31556
rect 22306 31500 22316 31556
rect 22372 31500 22540 31556
rect 22596 31500 23772 31556
rect 23828 31500 23838 31556
rect 38546 31500 38556 31556
rect 38612 31500 40684 31556
rect 40740 31500 40750 31556
rect 42466 31500 42476 31556
rect 42532 31500 42542 31556
rect 42476 31444 42532 31500
rect 4610 31388 4620 31444
rect 4676 31388 4956 31444
rect 5012 31388 5022 31444
rect 5730 31388 5740 31444
rect 5796 31388 6188 31444
rect 6244 31388 6524 31444
rect 6580 31388 6590 31444
rect 14802 31388 14812 31444
rect 14868 31388 15316 31444
rect 21746 31388 21756 31444
rect 21812 31388 22876 31444
rect 22932 31388 22942 31444
rect 42018 31388 42028 31444
rect 42084 31388 42532 31444
rect 15260 31332 15316 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 14998 31276 15036 31332
rect 15092 31276 15102 31332
rect 15250 31276 15260 31332
rect 15316 31276 15326 31332
rect 21858 31276 21868 31332
rect 21924 31276 24780 31332
rect 24836 31276 24846 31332
rect 31490 31276 31500 31332
rect 31556 31276 31724 31332
rect 31780 31276 31790 31332
rect 0 31220 800 31248
rect 49200 31220 50000 31248
rect 0 31164 1932 31220
rect 1988 31164 1998 31220
rect 8082 31164 8092 31220
rect 8148 31164 9660 31220
rect 9716 31164 9726 31220
rect 28802 31164 28812 31220
rect 28868 31164 31948 31220
rect 32004 31164 32014 31220
rect 48178 31164 48188 31220
rect 48244 31164 50000 31220
rect 0 31136 800 31164
rect 49200 31136 50000 31164
rect 7186 31052 7196 31108
rect 7252 31052 7588 31108
rect 7746 31052 7756 31108
rect 7812 31052 10108 31108
rect 10164 31052 10174 31108
rect 16034 31052 16044 31108
rect 16100 31052 17500 31108
rect 17556 31052 17566 31108
rect 7532 30996 7588 31052
rect 4834 30940 4844 30996
rect 4900 30940 6412 30996
rect 6468 30940 7308 30996
rect 7364 30940 7374 30996
rect 7532 30940 8316 30996
rect 8372 30940 9548 30996
rect 9604 30940 9614 30996
rect 9874 30940 9884 30996
rect 9940 30940 12124 30996
rect 12180 30940 12190 30996
rect 14018 30940 14028 30996
rect 14084 30940 15652 30996
rect 16370 30940 16380 30996
rect 16436 30940 17388 30996
rect 17444 30940 17454 30996
rect 18386 30940 18396 30996
rect 18452 30940 20076 30996
rect 20132 30940 22540 30996
rect 22596 30940 22606 30996
rect 29026 30940 29036 30996
rect 29092 30940 29820 30996
rect 29876 30940 29886 30996
rect 30818 30940 30828 30996
rect 30884 30940 31388 30996
rect 31444 30940 31454 30996
rect 15596 30884 15652 30940
rect 2930 30828 2940 30884
rect 2996 30828 4956 30884
rect 5012 30828 5022 30884
rect 7858 30828 7868 30884
rect 7924 30828 8652 30884
rect 8708 30828 8718 30884
rect 10770 30828 10780 30884
rect 10836 30828 11788 30884
rect 11844 30828 11854 30884
rect 15092 30828 15372 30884
rect 15428 30828 15438 30884
rect 15596 30828 16268 30884
rect 16324 30828 16334 30884
rect 16706 30828 16716 30884
rect 16772 30828 18284 30884
rect 18340 30828 18350 30884
rect 20514 30828 20524 30884
rect 20580 30828 23212 30884
rect 23268 30828 23884 30884
rect 23940 30828 23950 30884
rect 28466 30828 28476 30884
rect 28532 30828 29932 30884
rect 29988 30828 31948 30884
rect 32004 30828 32014 30884
rect 5478 30604 5516 30660
rect 5572 30604 5582 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 15092 30436 15148 30828
rect 32050 30716 32060 30772
rect 32116 30716 33292 30772
rect 33348 30716 35308 30772
rect 35364 30716 35374 30772
rect 41234 30716 41244 30772
rect 41300 30716 42252 30772
rect 42308 30716 42318 30772
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 14018 30380 14028 30436
rect 14084 30380 28700 30436
rect 28756 30380 28766 30436
rect 44342 30380 44380 30436
rect 44436 30380 44446 30436
rect 1922 30268 1932 30324
rect 1988 30268 3276 30324
rect 3332 30268 3342 30324
rect 7746 30268 7756 30324
rect 7812 30268 8428 30324
rect 8484 30268 8494 30324
rect 14130 30268 14140 30324
rect 14196 30268 14644 30324
rect 15138 30268 15148 30324
rect 15204 30268 16380 30324
rect 16436 30268 16446 30324
rect 5170 30156 5180 30212
rect 5236 30156 5964 30212
rect 6020 30156 6030 30212
rect 14326 30156 14364 30212
rect 14420 30156 14430 30212
rect 8866 30044 8876 30100
rect 8932 30044 11340 30100
rect 11396 30044 11406 30100
rect 14588 29988 14644 30268
rect 14802 30156 14812 30212
rect 14868 30156 15596 30212
rect 15652 30156 16716 30212
rect 16772 30156 16782 30212
rect 20738 30156 20748 30212
rect 20804 30156 21196 30212
rect 21252 30156 23548 30212
rect 23604 30156 23614 30212
rect 23986 30156 23996 30212
rect 24052 30156 27020 30212
rect 27076 30156 27244 30212
rect 27300 30156 27310 30212
rect 28028 30100 28084 30380
rect 28242 30156 28252 30212
rect 28308 30156 29260 30212
rect 29316 30156 29326 30212
rect 34738 30156 34748 30212
rect 34804 30156 35420 30212
rect 35476 30156 35486 30212
rect 36194 30156 36204 30212
rect 36260 30156 36988 30212
rect 37044 30156 37054 30212
rect 41122 30156 41132 30212
rect 41188 30156 42364 30212
rect 42420 30156 42430 30212
rect 42578 30156 42588 30212
rect 42644 30156 43484 30212
rect 43540 30156 45724 30212
rect 45780 30156 45790 30212
rect 17378 30044 17388 30100
rect 17444 30044 18060 30100
rect 18116 30044 18620 30100
rect 18676 30044 18686 30100
rect 28018 30044 28028 30100
rect 28084 30044 28094 30100
rect 28466 30044 28476 30100
rect 28532 30044 29372 30100
rect 29428 30044 30044 30100
rect 30100 30044 30110 30100
rect 34514 30044 34524 30100
rect 34580 30044 35868 30100
rect 35924 30044 35934 30100
rect 40338 30044 40348 30100
rect 40404 30044 41356 30100
rect 41412 30044 41422 30100
rect 1698 29932 1708 29988
rect 1764 29932 2268 29988
rect 2324 29932 2334 29988
rect 11414 29932 11452 29988
rect 11508 29932 11518 29988
rect 14578 29932 14588 29988
rect 14644 29932 15036 29988
rect 15092 29932 15102 29988
rect 17602 29932 17612 29988
rect 17668 29932 19292 29988
rect 19348 29932 19358 29988
rect 21858 29932 21868 29988
rect 21924 29932 23548 29988
rect 33842 29932 33852 29988
rect 33908 29932 35980 29988
rect 36036 29932 36046 29988
rect 36194 29932 36204 29988
rect 36260 29932 37100 29988
rect 37156 29932 37166 29988
rect 23492 29876 23548 29932
rect 36204 29876 36260 29932
rect 5730 29820 5740 29876
rect 5796 29820 6076 29876
rect 6132 29820 6636 29876
rect 6692 29820 16324 29876
rect 16594 29820 16604 29876
rect 16660 29820 18172 29876
rect 18228 29820 18956 29876
rect 19012 29820 19022 29876
rect 23492 29820 26908 29876
rect 29558 29820 29596 29876
rect 29652 29820 29662 29876
rect 33954 29820 33964 29876
rect 34020 29820 36260 29876
rect 36316 29820 38444 29876
rect 38500 29820 39116 29876
rect 39172 29820 39564 29876
rect 39620 29820 39630 29876
rect 16268 29764 16324 29820
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 26852 29764 26908 29820
rect 36316 29764 36372 29820
rect 16268 29708 18508 29764
rect 18564 29708 18574 29764
rect 26852 29708 36372 29764
rect 38612 29708 40012 29764
rect 40068 29708 40572 29764
rect 40628 29708 40908 29764
rect 40964 29708 40974 29764
rect 38612 29652 38668 29708
rect 40348 29652 40404 29708
rect 4386 29596 4396 29652
rect 4452 29596 5404 29652
rect 5460 29596 7532 29652
rect 7588 29596 7598 29652
rect 10546 29596 10556 29652
rect 10612 29596 16604 29652
rect 16660 29596 16670 29652
rect 20178 29596 20188 29652
rect 20244 29596 20636 29652
rect 20692 29596 21644 29652
rect 21700 29596 21710 29652
rect 24658 29596 24668 29652
rect 24724 29596 24892 29652
rect 24948 29596 25452 29652
rect 25508 29596 26236 29652
rect 26292 29596 26302 29652
rect 29670 29596 29708 29652
rect 29764 29596 29774 29652
rect 35074 29596 35084 29652
rect 35140 29596 38668 29652
rect 40338 29596 40348 29652
rect 40404 29596 40414 29652
rect 43474 29596 43484 29652
rect 43540 29596 43932 29652
rect 43988 29596 44604 29652
rect 44660 29596 47180 29652
rect 47236 29596 47246 29652
rect 14700 29540 14756 29596
rect 5506 29484 5516 29540
rect 5572 29484 5740 29540
rect 5796 29484 5806 29540
rect 11218 29484 11228 29540
rect 11284 29484 11788 29540
rect 14690 29484 14700 29540
rect 14756 29484 14766 29540
rect 17266 29484 17276 29540
rect 17332 29484 18396 29540
rect 18452 29484 18844 29540
rect 18900 29484 19404 29540
rect 19460 29484 19470 29540
rect 25554 29484 25564 29540
rect 25620 29484 27356 29540
rect 27412 29484 27422 29540
rect 11732 29428 11788 29484
rect 11732 29372 11900 29428
rect 11956 29372 14364 29428
rect 14420 29372 14430 29428
rect 26786 29372 26796 29428
rect 26852 29372 29484 29428
rect 29540 29372 29550 29428
rect 31938 29372 31948 29428
rect 32004 29372 32732 29428
rect 32788 29372 32798 29428
rect 40674 29372 40684 29428
rect 40740 29372 41468 29428
rect 41524 29372 41534 29428
rect 42690 29372 42700 29428
rect 42756 29372 43596 29428
rect 43652 29372 43932 29428
rect 43988 29372 43998 29428
rect 1810 29260 1820 29316
rect 1876 29260 4844 29316
rect 4900 29260 4910 29316
rect 29586 29260 29596 29316
rect 29652 29260 30156 29316
rect 30212 29260 30222 29316
rect 39554 29260 39564 29316
rect 39620 29260 39900 29316
rect 39956 29260 39966 29316
rect 40226 29260 40236 29316
rect 40292 29260 40460 29316
rect 40516 29260 40526 29316
rect 8978 29148 8988 29204
rect 9044 29148 9772 29204
rect 9828 29148 9838 29204
rect 11414 29148 11452 29204
rect 11508 29148 11518 29204
rect 26338 29148 26348 29204
rect 26404 29148 26852 29204
rect 38966 29148 39004 29204
rect 39060 29148 39070 29204
rect 26796 29092 26852 29148
rect 5730 29036 5740 29092
rect 5796 29036 6076 29092
rect 6132 29036 6142 29092
rect 26786 29036 26796 29092
rect 26852 29036 26862 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 40450 28924 40460 28980
rect 40516 28924 41244 28980
rect 41300 28924 41310 28980
rect 25442 28812 25452 28868
rect 25508 28812 26012 28868
rect 26068 28812 27580 28868
rect 27636 28812 27646 28868
rect 35074 28812 35084 28868
rect 35140 28812 35308 28868
rect 35364 28812 35374 28868
rect 39442 28812 39452 28868
rect 39508 28812 43372 28868
rect 43428 28812 45164 28868
rect 45220 28812 45948 28868
rect 46004 28812 46014 28868
rect 0 28756 800 28784
rect 49200 28756 50000 28784
rect 0 28700 1820 28756
rect 1876 28700 1886 28756
rect 4610 28700 4620 28756
rect 4676 28700 5852 28756
rect 5908 28700 5918 28756
rect 9426 28700 9436 28756
rect 9492 28700 11228 28756
rect 11284 28700 11294 28756
rect 15586 28700 15596 28756
rect 15652 28700 16380 28756
rect 16436 28700 17052 28756
rect 17108 28700 17118 28756
rect 18498 28700 18508 28756
rect 18564 28700 19852 28756
rect 19908 28700 19918 28756
rect 21074 28700 21084 28756
rect 21140 28700 24220 28756
rect 24276 28700 24286 28756
rect 38098 28700 38108 28756
rect 38164 28700 43484 28756
rect 43540 28700 43550 28756
rect 45266 28700 45276 28756
rect 45332 28700 46620 28756
rect 46676 28700 46686 28756
rect 48188 28700 50000 28756
rect 0 28672 800 28700
rect 1698 28588 1708 28644
rect 1764 28588 2604 28644
rect 2660 28588 5068 28644
rect 5124 28588 5134 28644
rect 10770 28588 10780 28644
rect 10836 28588 11564 28644
rect 11620 28588 11630 28644
rect 19170 28588 19180 28644
rect 19236 28588 21532 28644
rect 21588 28588 22652 28644
rect 22708 28588 22718 28644
rect 27010 28588 27020 28644
rect 27076 28588 27580 28644
rect 27636 28588 28252 28644
rect 28308 28588 28318 28644
rect 35410 28588 35420 28644
rect 35476 28588 35980 28644
rect 36036 28588 36046 28644
rect 37090 28588 37100 28644
rect 37156 28588 39116 28644
rect 39172 28588 39182 28644
rect 43698 28588 43708 28644
rect 43764 28588 43774 28644
rect 43708 28532 43764 28588
rect 48188 28532 48244 28700
rect 49200 28672 50000 28700
rect 9874 28476 9884 28532
rect 9940 28476 10668 28532
rect 10724 28476 11116 28532
rect 11172 28476 11182 28532
rect 14662 28476 14700 28532
rect 14756 28476 14766 28532
rect 21634 28476 21644 28532
rect 21700 28476 22092 28532
rect 22148 28476 22158 28532
rect 31602 28476 31612 28532
rect 31668 28476 31948 28532
rect 32004 28476 32620 28532
rect 32676 28476 32686 28532
rect 34962 28476 34972 28532
rect 35028 28476 35196 28532
rect 35252 28476 35868 28532
rect 35924 28476 35934 28532
rect 37650 28476 37660 28532
rect 37716 28476 38668 28532
rect 38724 28476 38734 28532
rect 38994 28476 39004 28532
rect 39060 28476 39340 28532
rect 39396 28476 39406 28532
rect 43708 28476 45388 28532
rect 45444 28476 45454 28532
rect 48178 28476 48188 28532
rect 48244 28476 48254 28532
rect 14914 28364 14924 28420
rect 14980 28364 15260 28420
rect 15316 28364 15326 28420
rect 26982 28364 27020 28420
rect 27076 28364 27086 28420
rect 28018 28364 28028 28420
rect 28084 28364 30828 28420
rect 30884 28364 32060 28420
rect 32116 28364 32126 28420
rect 38770 28364 38780 28420
rect 38836 28364 39452 28420
rect 39508 28364 39518 28420
rect 10780 28252 11004 28308
rect 11060 28252 11070 28308
rect 10780 28196 10836 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 10770 28140 10780 28196
rect 10836 28140 10846 28196
rect 11004 28140 11564 28196
rect 11620 28140 12236 28196
rect 12292 28140 12796 28196
rect 12852 28140 12862 28196
rect 13990 28140 14028 28196
rect 14084 28140 14094 28196
rect 11004 28084 11060 28140
rect 10994 28028 11004 28084
rect 11060 28028 11070 28084
rect 11778 28028 11788 28084
rect 11844 28028 12348 28084
rect 12404 28028 12414 28084
rect 20514 28028 20524 28084
rect 20580 28028 32060 28084
rect 32116 28028 32126 28084
rect 37538 28028 37548 28084
rect 37604 28028 39004 28084
rect 39060 28028 39070 28084
rect 39330 28028 39340 28084
rect 39396 28028 40236 28084
rect 40292 28028 40302 28084
rect 13570 27916 13580 27972
rect 13636 27916 14476 27972
rect 14532 27916 14542 27972
rect 21522 27916 21532 27972
rect 21588 27916 22764 27972
rect 22820 27916 22830 27972
rect 23398 27916 23436 27972
rect 23492 27916 23502 27972
rect 28466 27916 28476 27972
rect 28532 27916 29708 27972
rect 29764 27916 29774 27972
rect 35298 27916 35308 27972
rect 35364 27916 35868 27972
rect 35924 27916 35934 27972
rect 39554 27916 39564 27972
rect 39620 27916 40124 27972
rect 40180 27916 40190 27972
rect 2258 27804 2268 27860
rect 2324 27804 2940 27860
rect 2996 27804 3612 27860
rect 3668 27804 3678 27860
rect 10098 27804 10108 27860
rect 10164 27804 12012 27860
rect 12068 27804 12348 27860
rect 12404 27804 12414 27860
rect 15250 27804 15260 27860
rect 15316 27804 15820 27860
rect 15876 27804 15886 27860
rect 17714 27804 17724 27860
rect 17780 27804 19404 27860
rect 19460 27804 19470 27860
rect 21942 27804 21980 27860
rect 22036 27804 22046 27860
rect 38546 27804 38556 27860
rect 38612 27804 40348 27860
rect 40404 27804 40414 27860
rect 12450 27692 12460 27748
rect 12516 27692 13244 27748
rect 13300 27692 13804 27748
rect 13860 27692 13870 27748
rect 20514 27692 20524 27748
rect 20580 27692 29708 27748
rect 29764 27692 29774 27748
rect 30594 27692 30604 27748
rect 30660 27692 31388 27748
rect 31444 27692 31454 27748
rect 11778 27580 11788 27636
rect 11844 27580 12796 27636
rect 12852 27580 12862 27636
rect 17042 27580 17052 27636
rect 17108 27580 18060 27636
rect 18116 27580 18126 27636
rect 23090 27580 23100 27636
rect 23156 27580 23996 27636
rect 24052 27580 24062 27636
rect 30258 27580 30268 27636
rect 30324 27580 31612 27636
rect 31668 27580 33180 27636
rect 33236 27580 33246 27636
rect 35634 27580 35644 27636
rect 35700 27580 36092 27636
rect 36148 27580 40236 27636
rect 40292 27580 40302 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 37660 27356 38332 27412
rect 38388 27356 38398 27412
rect 39778 27356 39788 27412
rect 39844 27356 41020 27412
rect 41076 27356 41086 27412
rect 37660 27300 37716 27356
rect 6738 27244 6748 27300
rect 6804 27244 7420 27300
rect 7476 27244 19404 27300
rect 19460 27244 20412 27300
rect 20468 27244 20478 27300
rect 20626 27244 20636 27300
rect 20692 27244 21868 27300
rect 21924 27244 21934 27300
rect 32722 27244 32732 27300
rect 32788 27244 35308 27300
rect 35364 27244 35374 27300
rect 37622 27244 37660 27300
rect 37716 27244 37726 27300
rect 37986 27244 37996 27300
rect 38052 27244 38780 27300
rect 38836 27244 38846 27300
rect 41234 27244 41244 27300
rect 41300 27244 46284 27300
rect 46340 27244 46350 27300
rect 8194 27132 8204 27188
rect 8260 27132 8876 27188
rect 8932 27132 8942 27188
rect 11106 27132 11116 27188
rect 11172 27132 12012 27188
rect 12068 27132 12078 27188
rect 12338 27132 12348 27188
rect 12404 27132 13020 27188
rect 13076 27132 13086 27188
rect 13580 27132 14700 27188
rect 14756 27132 14766 27188
rect 21634 27132 21644 27188
rect 21700 27132 22764 27188
rect 22820 27132 23772 27188
rect 23828 27132 23838 27188
rect 25554 27132 25564 27188
rect 25620 27132 36988 27188
rect 37044 27132 37054 27188
rect 13580 27076 13636 27132
rect 2594 27020 2604 27076
rect 2660 27020 3276 27076
rect 3332 27020 3342 27076
rect 12684 27020 13580 27076
rect 13636 27020 13646 27076
rect 13906 27020 13916 27076
rect 13972 27020 15932 27076
rect 15988 27020 15998 27076
rect 16594 27020 16604 27076
rect 16660 27020 16940 27076
rect 16996 27020 17612 27076
rect 17668 27020 17678 27076
rect 17826 27020 17836 27076
rect 17892 27020 17930 27076
rect 20738 27020 20748 27076
rect 20804 27020 24220 27076
rect 24276 27020 24286 27076
rect 32050 27020 32060 27076
rect 32116 27020 32844 27076
rect 32900 27020 32910 27076
rect 33058 27020 33068 27076
rect 33124 27020 33628 27076
rect 33684 27020 33694 27076
rect 38658 27020 38668 27076
rect 38724 27020 39900 27076
rect 39956 27020 39966 27076
rect 12684 26964 12740 27020
rect 2930 26908 2940 26964
rect 2996 26908 4060 26964
rect 4116 26908 4126 26964
rect 4946 26908 4956 26964
rect 5012 26908 5852 26964
rect 5908 26908 5918 26964
rect 10994 26908 11004 26964
rect 11060 26908 12180 26964
rect 12674 26908 12684 26964
rect 12740 26908 12750 26964
rect 13010 26908 13020 26964
rect 13076 26908 13636 26964
rect 14466 26908 14476 26964
rect 14532 26908 17724 26964
rect 17780 26908 17790 26964
rect 21858 26908 21868 26964
rect 21924 26908 22764 26964
rect 22820 26908 23100 26964
rect 23156 26908 23166 26964
rect 30828 26908 31500 26964
rect 31556 26908 31566 26964
rect 45154 26908 45164 26964
rect 45220 26908 45724 26964
rect 45780 26908 45790 26964
rect 12114 26852 12124 26908
rect 12180 26852 12190 26908
rect 13580 26852 13636 26908
rect 30818 26852 30828 26908
rect 30884 26852 30894 26908
rect 12534 26796 12572 26852
rect 12628 26796 12638 26852
rect 13570 26796 13580 26852
rect 13636 26796 13646 26852
rect 16146 26796 16156 26852
rect 16212 26796 18508 26852
rect 18564 26796 18574 26852
rect 27682 26796 27692 26852
rect 27748 26796 28028 26852
rect 28084 26796 28094 26852
rect 31686 26796 31724 26852
rect 31780 26796 31790 26852
rect 17602 26684 17612 26740
rect 17668 26684 18284 26740
rect 18340 26684 18350 26740
rect 26982 26684 27020 26740
rect 27076 26684 27086 26740
rect 30930 26684 30940 26740
rect 30996 26684 31006 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 30940 26628 30996 26684
rect 9986 26572 9996 26628
rect 10052 26572 10332 26628
rect 10388 26572 10398 26628
rect 30940 26572 31164 26628
rect 31220 26572 31230 26628
rect 34710 26572 34748 26628
rect 34804 26572 34814 26628
rect 16482 26460 16492 26516
rect 16548 26460 16716 26516
rect 16772 26460 16782 26516
rect 22082 26460 22092 26516
rect 22148 26460 22158 26516
rect 33506 26460 33516 26516
rect 33572 26460 39004 26516
rect 39060 26460 39070 26516
rect 46610 26460 46620 26516
rect 46676 26460 47404 26516
rect 47460 26460 47470 26516
rect 0 26292 800 26320
rect 22092 26292 22148 26460
rect 28690 26348 28700 26404
rect 28756 26348 28924 26404
rect 28980 26348 28990 26404
rect 31266 26348 31276 26404
rect 31332 26348 31342 26404
rect 31276 26292 31332 26348
rect 49200 26292 50000 26320
rect 0 26236 1708 26292
rect 1764 26236 1774 26292
rect 5058 26236 5068 26292
rect 5124 26236 5628 26292
rect 5684 26236 8988 26292
rect 9044 26236 9054 26292
rect 22092 26236 23772 26292
rect 23828 26236 23838 26292
rect 27906 26236 27916 26292
rect 27972 26236 29148 26292
rect 29204 26236 29214 26292
rect 31276 26236 31612 26292
rect 31668 26236 31678 26292
rect 32610 26236 32620 26292
rect 32676 26236 33852 26292
rect 33908 26236 33918 26292
rect 38612 26236 46732 26292
rect 46788 26236 46798 26292
rect 48178 26236 48188 26292
rect 48244 26236 50000 26292
rect 0 26208 800 26236
rect 38612 26180 38668 26236
rect 49200 26208 50000 26236
rect 9762 26124 9772 26180
rect 9828 26124 10556 26180
rect 10612 26124 10622 26180
rect 16370 26124 16380 26180
rect 16436 26124 18284 26180
rect 18340 26124 18350 26180
rect 24994 26124 25004 26180
rect 25060 26124 38668 26180
rect 44146 26124 44156 26180
rect 44212 26124 44828 26180
rect 44884 26124 45164 26180
rect 45220 26124 45230 26180
rect 15810 26012 15820 26068
rect 15876 26012 16492 26068
rect 16548 26012 16558 26068
rect 27458 26012 27468 26068
rect 27524 26012 44044 26068
rect 44100 26012 44110 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 18694 25788 18732 25844
rect 18788 25788 18798 25844
rect 14242 25676 14252 25732
rect 14308 25676 15148 25732
rect 15204 25676 15708 25732
rect 15764 25676 15774 25732
rect 5842 25564 5852 25620
rect 5908 25564 6748 25620
rect 6804 25564 7756 25620
rect 7812 25564 7822 25620
rect 18722 25564 18732 25620
rect 18788 25564 20748 25620
rect 20804 25564 21532 25620
rect 21588 25564 21598 25620
rect 45378 25564 45388 25620
rect 45444 25564 46284 25620
rect 46340 25564 46350 25620
rect 4610 25452 4620 25508
rect 4676 25452 5292 25508
rect 5348 25452 5628 25508
rect 5684 25452 5694 25508
rect 14326 25452 14364 25508
rect 14420 25452 14430 25508
rect 18274 25452 18284 25508
rect 18340 25452 20636 25508
rect 20692 25452 20702 25508
rect 27122 25452 27132 25508
rect 27188 25452 27468 25508
rect 27524 25452 28028 25508
rect 28084 25452 29036 25508
rect 29092 25452 29102 25508
rect 46386 25452 46396 25508
rect 46452 25452 46620 25508
rect 46676 25452 46686 25508
rect 8978 25340 8988 25396
rect 9044 25340 11788 25396
rect 11844 25340 11854 25396
rect 18956 25340 21420 25396
rect 21476 25340 21486 25396
rect 46470 25340 46508 25396
rect 46564 25340 46574 25396
rect 18956 25284 19012 25340
rect 5842 25228 5852 25284
rect 5908 25228 7420 25284
rect 7476 25228 7486 25284
rect 8306 25228 8316 25284
rect 8372 25228 9100 25284
rect 9156 25228 9166 25284
rect 10882 25228 10892 25284
rect 10948 25228 12460 25284
rect 12516 25228 12526 25284
rect 14214 25228 14252 25284
rect 14308 25228 14700 25284
rect 14756 25228 14766 25284
rect 18498 25228 18508 25284
rect 18564 25228 19012 25284
rect 20066 25228 20076 25284
rect 20132 25228 21196 25284
rect 21252 25228 21262 25284
rect 42130 25228 42140 25284
rect 42196 25228 42476 25284
rect 42532 25228 42542 25284
rect 18956 25172 19012 25228
rect 4274 25116 4284 25172
rect 4340 25116 5180 25172
rect 5236 25116 5246 25172
rect 14998 25116 15036 25172
rect 15092 25116 15102 25172
rect 18946 25116 18956 25172
rect 19012 25116 19022 25172
rect 38770 25116 38780 25172
rect 38836 25116 39564 25172
rect 39620 25116 39630 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 4834 25004 4844 25060
rect 4900 25004 6076 25060
rect 6132 25004 6860 25060
rect 6916 25004 6926 25060
rect 25218 25004 25228 25060
rect 25284 25004 25900 25060
rect 25956 25004 25966 25060
rect 37958 25004 37996 25060
rect 38052 25004 38444 25060
rect 38500 25004 38510 25060
rect 39442 25004 39452 25060
rect 39508 25004 39900 25060
rect 39956 25004 39966 25060
rect 11106 24892 11116 24948
rect 11172 24892 11788 24948
rect 11844 24892 11882 24948
rect 26338 24892 26348 24948
rect 26404 24892 27692 24948
rect 27748 24892 27758 24948
rect 31826 24892 31836 24948
rect 31892 24892 33964 24948
rect 34020 24892 34030 24948
rect 37202 24892 37212 24948
rect 37268 24892 37884 24948
rect 37940 24892 37950 24948
rect 4722 24780 4732 24836
rect 4788 24780 6412 24836
rect 6468 24780 6478 24836
rect 19954 24780 19964 24836
rect 20020 24780 20860 24836
rect 20916 24780 20926 24836
rect 26450 24780 26460 24836
rect 26516 24780 27132 24836
rect 27188 24780 27198 24836
rect 40002 24780 40012 24836
rect 40068 24780 41132 24836
rect 41188 24780 41692 24836
rect 41748 24780 41758 24836
rect 41906 24780 41916 24836
rect 41972 24780 42588 24836
rect 42644 24780 43148 24836
rect 43204 24780 43214 24836
rect 17266 24668 17276 24724
rect 17332 24668 18060 24724
rect 18116 24668 20300 24724
rect 20356 24668 20366 24724
rect 25442 24668 25452 24724
rect 25508 24668 29148 24724
rect 29204 24668 29214 24724
rect 33506 24668 33516 24724
rect 33572 24668 33964 24724
rect 34020 24668 34030 24724
rect 39778 24668 39788 24724
rect 39844 24668 40348 24724
rect 40404 24668 41020 24724
rect 41076 24668 41086 24724
rect 41570 24668 41580 24724
rect 41636 24668 42924 24724
rect 42980 24668 42990 24724
rect 43586 24668 43596 24724
rect 43652 24668 44044 24724
rect 44100 24668 44110 24724
rect 44818 24668 44828 24724
rect 44884 24668 45388 24724
rect 45444 24668 45454 24724
rect 23398 24556 23436 24612
rect 23492 24556 23502 24612
rect 28578 24556 28588 24612
rect 28644 24556 29708 24612
rect 29764 24556 29774 24612
rect 35858 24556 35868 24612
rect 35924 24556 37660 24612
rect 37716 24556 37726 24612
rect 42690 24556 42700 24612
rect 42756 24556 43036 24612
rect 43092 24556 43708 24612
rect 43764 24556 43774 24612
rect 11106 24444 11116 24500
rect 11172 24444 11452 24500
rect 11508 24444 11518 24500
rect 43810 24444 43820 24500
rect 43876 24444 45052 24500
rect 45108 24444 45118 24500
rect 13990 24332 14028 24388
rect 14084 24332 14094 24388
rect 24098 24332 24108 24388
rect 24164 24332 25676 24388
rect 25732 24332 25742 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 29698 24220 29708 24276
rect 29764 24220 29774 24276
rect 29708 24164 29764 24220
rect 29708 24108 46732 24164
rect 46788 24108 46798 24164
rect 1586 23996 1596 24052
rect 1652 23996 2268 24052
rect 2324 23996 2334 24052
rect 12226 23996 12236 24052
rect 12292 23996 12572 24052
rect 12628 23996 12638 24052
rect 26114 23996 26124 24052
rect 26180 23996 26460 24052
rect 26516 23996 26526 24052
rect 44370 23996 44380 24052
rect 44436 23996 44940 24052
rect 44996 23996 45006 24052
rect 10098 23884 10108 23940
rect 10164 23884 10780 23940
rect 10836 23884 10846 23940
rect 12114 23884 12124 23940
rect 12180 23884 12796 23940
rect 12852 23884 12862 23940
rect 23202 23884 23212 23940
rect 23268 23884 25452 23940
rect 25508 23884 25518 23940
rect 31602 23884 31612 23940
rect 31668 23884 31948 23940
rect 32004 23884 32014 23940
rect 0 23828 800 23856
rect 49200 23828 50000 23856
rect 0 23772 1708 23828
rect 1764 23772 1774 23828
rect 18498 23772 18508 23828
rect 18564 23772 20188 23828
rect 20244 23772 20254 23828
rect 22866 23772 22876 23828
rect 22932 23772 23548 23828
rect 23604 23772 23614 23828
rect 25106 23772 25116 23828
rect 25172 23772 34076 23828
rect 34132 23772 34142 23828
rect 48066 23772 48076 23828
rect 48132 23772 50000 23828
rect 0 23744 800 23772
rect 49200 23744 50000 23772
rect 10770 23660 10780 23716
rect 10836 23660 11340 23716
rect 11396 23660 11406 23716
rect 19282 23660 19292 23716
rect 19348 23660 19852 23716
rect 19908 23660 21420 23716
rect 21476 23660 21486 23716
rect 23986 23660 23996 23716
rect 24052 23660 26348 23716
rect 26404 23660 26414 23716
rect 29558 23660 29596 23716
rect 29652 23660 29662 23716
rect 33058 23660 33068 23716
rect 33124 23660 33964 23716
rect 34020 23660 34030 23716
rect 37650 23660 37660 23716
rect 37716 23660 38668 23716
rect 38612 23604 38668 23660
rect 3602 23548 3612 23604
rect 3668 23548 6412 23604
rect 6468 23548 6478 23604
rect 13794 23548 13804 23604
rect 13860 23548 14588 23604
rect 14644 23548 14654 23604
rect 15474 23548 15484 23604
rect 15540 23548 16716 23604
rect 16772 23548 16782 23604
rect 22978 23548 22988 23604
rect 23044 23548 24220 23604
rect 24276 23548 24286 23604
rect 38612 23548 42700 23604
rect 42756 23548 42766 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 17378 23436 17388 23492
rect 17444 23436 18732 23492
rect 18788 23436 18798 23492
rect 28130 23436 28140 23492
rect 28196 23436 28868 23492
rect 37398 23436 37436 23492
rect 37492 23436 37502 23492
rect 39778 23436 39788 23492
rect 39844 23436 40236 23492
rect 40292 23436 40908 23492
rect 40964 23436 41580 23492
rect 41636 23436 41646 23492
rect 28812 23380 28868 23436
rect 5842 23324 5852 23380
rect 5908 23324 6860 23380
rect 6916 23324 6926 23380
rect 27570 23324 27580 23380
rect 27636 23324 28532 23380
rect 28802 23324 28812 23380
rect 28868 23324 29932 23380
rect 29988 23324 45500 23380
rect 45556 23324 45566 23380
rect 45826 23324 45836 23380
rect 45892 23324 46172 23380
rect 46228 23324 46238 23380
rect 10322 23212 10332 23268
rect 10388 23212 11340 23268
rect 11396 23212 11406 23268
rect 13122 23212 13132 23268
rect 13188 23212 13916 23268
rect 13972 23212 13982 23268
rect 15586 23212 15596 23268
rect 15652 23212 16156 23268
rect 16212 23212 16222 23268
rect 28476 23156 28532 23324
rect 33842 23212 33852 23268
rect 33908 23212 35532 23268
rect 35588 23212 35598 23268
rect 38322 23212 38332 23268
rect 38388 23212 39396 23268
rect 39340 23156 39396 23212
rect 10210 23100 10220 23156
rect 10276 23100 11676 23156
rect 11732 23100 12796 23156
rect 12852 23100 12862 23156
rect 26674 23100 26684 23156
rect 26740 23100 27580 23156
rect 27636 23100 27646 23156
rect 28466 23100 28476 23156
rect 28532 23100 29148 23156
rect 29204 23100 38668 23156
rect 39330 23100 39340 23156
rect 39396 23100 39406 23156
rect 38612 23044 38668 23100
rect 6178 22988 6188 23044
rect 6244 22988 7644 23044
rect 7700 22988 7710 23044
rect 10770 22988 10780 23044
rect 10836 22988 12684 23044
rect 12740 22988 12750 23044
rect 14578 22988 14588 23044
rect 14644 22988 14924 23044
rect 14980 22988 14990 23044
rect 25778 22988 25788 23044
rect 25844 22988 33852 23044
rect 33908 22988 33918 23044
rect 34066 22988 34076 23044
rect 34132 22988 34972 23044
rect 35028 22988 35308 23044
rect 35364 22988 35374 23044
rect 38612 22988 45388 23044
rect 45444 22988 45454 23044
rect 14354 22876 14364 22932
rect 14420 22876 14812 22932
rect 14868 22876 14878 22932
rect 38630 22764 38668 22820
rect 38724 22764 38734 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14998 22652 15036 22708
rect 15092 22652 15102 22708
rect 19394 22652 19404 22708
rect 19460 22652 20188 22708
rect 20244 22652 29372 22708
rect 29428 22652 29438 22708
rect 14690 22540 14700 22596
rect 14756 22540 15708 22596
rect 15764 22540 15774 22596
rect 17602 22540 17612 22596
rect 17668 22540 25900 22596
rect 25956 22540 26124 22596
rect 26180 22540 26190 22596
rect 39414 22540 39452 22596
rect 39508 22540 39518 22596
rect 7634 22428 7644 22484
rect 7700 22428 8540 22484
rect 8596 22428 9996 22484
rect 10052 22428 10062 22484
rect 11106 22428 11116 22484
rect 11172 22428 11788 22484
rect 11844 22428 11854 22484
rect 14578 22428 14588 22484
rect 14644 22428 15484 22484
rect 15540 22428 15550 22484
rect 19730 22428 19740 22484
rect 19796 22428 22092 22484
rect 22148 22428 22158 22484
rect 28802 22428 28812 22484
rect 28868 22428 29260 22484
rect 29316 22428 29326 22484
rect 40002 22428 40012 22484
rect 40068 22428 40572 22484
rect 40628 22428 40638 22484
rect 41458 22428 41468 22484
rect 41524 22428 42252 22484
rect 42308 22428 42318 22484
rect 8418 22316 8428 22372
rect 8484 22316 9772 22372
rect 9828 22316 9838 22372
rect 11890 22316 11900 22372
rect 11956 22316 13356 22372
rect 13412 22316 13422 22372
rect 20486 22316 20524 22372
rect 20580 22316 20590 22372
rect 21298 22316 21308 22372
rect 21364 22316 22204 22372
rect 22260 22316 22270 22372
rect 26226 22316 26236 22372
rect 26292 22316 27244 22372
rect 27300 22316 27310 22372
rect 37874 22316 37884 22372
rect 37940 22316 38556 22372
rect 38612 22316 38622 22372
rect 46162 22316 46172 22372
rect 46228 22316 47068 22372
rect 47124 22316 47134 22372
rect 18722 22204 18732 22260
rect 18788 22204 21084 22260
rect 21140 22204 21150 22260
rect 37426 22204 37436 22260
rect 37492 22204 38332 22260
rect 38388 22204 38398 22260
rect 45938 22204 45948 22260
rect 46004 22204 46844 22260
rect 46900 22204 46910 22260
rect 16818 22092 16828 22148
rect 16884 22092 18172 22148
rect 18228 22092 18238 22148
rect 20066 22092 20076 22148
rect 20132 22092 21532 22148
rect 21588 22092 22204 22148
rect 22260 22092 22270 22148
rect 26898 22092 26908 22148
rect 26964 22092 27244 22148
rect 27300 22092 27310 22148
rect 45266 22092 45276 22148
rect 45332 22092 46956 22148
rect 47012 22092 47022 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 13906 21868 13916 21924
rect 13972 21868 14700 21924
rect 14756 21868 18844 21924
rect 18900 21868 18910 21924
rect 20972 21812 21028 22092
rect 37426 21868 37436 21924
rect 37492 21868 39340 21924
rect 39396 21868 39406 21924
rect 45378 21868 45388 21924
rect 45444 21868 46396 21924
rect 46452 21868 46462 21924
rect 2258 21756 2268 21812
rect 2324 21756 6972 21812
rect 7028 21756 7038 21812
rect 9874 21756 9884 21812
rect 9940 21756 10892 21812
rect 10948 21756 11452 21812
rect 11508 21756 11518 21812
rect 14914 21756 14924 21812
rect 14980 21756 17276 21812
rect 17332 21756 17342 21812
rect 17938 21756 17948 21812
rect 18004 21756 18284 21812
rect 18340 21756 18350 21812
rect 20962 21756 20972 21812
rect 21028 21756 21038 21812
rect 42690 21756 42700 21812
rect 42756 21756 43260 21812
rect 43316 21756 43326 21812
rect 1250 21644 1260 21700
rect 1316 21644 26124 21700
rect 26180 21644 26190 21700
rect 5058 21532 5068 21588
rect 5124 21532 5628 21588
rect 5684 21532 8316 21588
rect 8372 21532 8382 21588
rect 15026 21532 15036 21588
rect 15092 21532 15820 21588
rect 15876 21532 15886 21588
rect 17602 21532 17612 21588
rect 17668 21532 18060 21588
rect 18116 21532 18228 21588
rect 20178 21532 20188 21588
rect 20244 21532 20636 21588
rect 20692 21532 20702 21588
rect 29698 21532 29708 21588
rect 29764 21532 30268 21588
rect 30324 21532 30334 21588
rect 0 21364 800 21392
rect 15484 21364 15540 21532
rect 0 21308 1708 21364
rect 1764 21308 1774 21364
rect 15474 21308 15484 21364
rect 15540 21308 15550 21364
rect 17154 21308 17164 21364
rect 17220 21308 17724 21364
rect 17780 21308 17790 21364
rect 0 21280 800 21308
rect 18172 21252 18228 21532
rect 49200 21364 50000 21392
rect 19506 21308 19516 21364
rect 19572 21308 20524 21364
rect 20580 21308 20590 21364
rect 48066 21308 48076 21364
rect 48132 21308 50000 21364
rect 49200 21280 50000 21308
rect 14802 21196 14812 21252
rect 14868 21196 17948 21252
rect 18004 21196 18014 21252
rect 18172 21196 20300 21252
rect 20356 21196 20366 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 15138 21084 15148 21140
rect 15204 21084 15708 21140
rect 15764 21084 15774 21140
rect 26226 20972 26236 21028
rect 26292 20972 26572 21028
rect 26628 20972 26638 21028
rect 26852 20916 26908 21140
rect 26964 21084 27244 21140
rect 27300 21084 28028 21140
rect 28084 21084 28588 21140
rect 28644 21084 28654 21140
rect 27010 20972 27020 21028
rect 27076 20972 27086 21028
rect 28802 20972 28812 21028
rect 28868 20972 33852 21028
rect 33908 20972 33918 21028
rect 12674 20860 12684 20916
rect 12740 20860 17836 20916
rect 17892 20860 17902 20916
rect 25218 20860 25228 20916
rect 25284 20860 25788 20916
rect 25844 20860 26908 20916
rect 27020 20804 27076 20972
rect 31714 20860 31724 20916
rect 31780 20860 32284 20916
rect 32340 20860 32620 20916
rect 32676 20860 33740 20916
rect 33796 20860 33806 20916
rect 39106 20860 39116 20916
rect 39172 20860 39788 20916
rect 39844 20860 39854 20916
rect 4050 20748 4060 20804
rect 4116 20748 5964 20804
rect 6020 20748 6030 20804
rect 16930 20748 16940 20804
rect 16996 20748 17724 20804
rect 17780 20748 17790 20804
rect 19282 20748 19292 20804
rect 19348 20748 21420 20804
rect 21476 20748 21486 20804
rect 26114 20748 26124 20804
rect 26180 20748 27076 20804
rect 30034 20748 30044 20804
rect 30100 20748 30716 20804
rect 30772 20748 30782 20804
rect 33282 20748 33292 20804
rect 33348 20748 46732 20804
rect 46788 20748 46798 20804
rect 19292 20692 19348 20748
rect 15586 20636 15596 20692
rect 15652 20636 19348 20692
rect 20178 20636 20188 20692
rect 20244 20636 20748 20692
rect 20804 20636 21196 20692
rect 21252 20636 21262 20692
rect 27346 20636 27356 20692
rect 27412 20636 28140 20692
rect 28196 20636 28588 20692
rect 28644 20636 44828 20692
rect 44884 20636 44894 20692
rect 11218 20524 11228 20580
rect 11284 20524 12124 20580
rect 12180 20524 12190 20580
rect 20066 20524 20076 20580
rect 20132 20524 20412 20580
rect 20468 20524 20478 20580
rect 25666 20524 25676 20580
rect 25732 20524 27804 20580
rect 27860 20524 27870 20580
rect 16706 20412 16716 20468
rect 16772 20412 17276 20468
rect 17332 20412 17342 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 17042 20300 17052 20356
rect 17108 20300 18844 20356
rect 18900 20300 18910 20356
rect 34290 20300 34300 20356
rect 34356 20300 34860 20356
rect 34916 20300 35196 20356
rect 35252 20300 36092 20356
rect 36148 20300 36158 20356
rect 39778 20300 39788 20356
rect 39844 20300 41020 20356
rect 41076 20300 41086 20356
rect 1138 20188 1148 20244
rect 1204 20188 22092 20244
rect 22148 20188 22540 20244
rect 22596 20188 22606 20244
rect 31602 20188 31612 20244
rect 31668 20188 31948 20244
rect 32004 20188 32396 20244
rect 32452 20188 33292 20244
rect 33348 20188 33358 20244
rect 34738 20188 34748 20244
rect 34804 20188 36428 20244
rect 36484 20188 36494 20244
rect 10994 20076 11004 20132
rect 11060 20076 12796 20132
rect 12852 20076 12862 20132
rect 17154 20076 17164 20132
rect 17220 20076 17948 20132
rect 18004 20076 18014 20132
rect 21522 20076 21532 20132
rect 21588 20076 22316 20132
rect 22372 20076 22382 20132
rect 23202 20076 23212 20132
rect 23268 20076 24220 20132
rect 24276 20076 24892 20132
rect 24948 20076 24958 20132
rect 25554 20076 25564 20132
rect 25620 20076 27244 20132
rect 27300 20076 27310 20132
rect 30818 20076 30828 20132
rect 30884 20076 31164 20132
rect 31220 20076 31230 20132
rect 31490 20076 31500 20132
rect 31556 20076 33068 20132
rect 33124 20076 33134 20132
rect 37314 20076 37324 20132
rect 37380 20076 38108 20132
rect 38164 20076 38174 20132
rect 38612 20076 39900 20132
rect 39956 20076 39966 20132
rect 3938 19964 3948 20020
rect 4004 19964 11396 20020
rect 14018 19964 14028 20020
rect 14084 19964 17276 20020
rect 17332 19964 17342 20020
rect 19730 19964 19740 20020
rect 19796 19964 21868 20020
rect 21924 19964 21934 20020
rect 30146 19964 30156 20020
rect 30212 19964 31388 20020
rect 31444 19964 31454 20020
rect 37874 19964 37884 20020
rect 37940 19964 38220 20020
rect 38276 19964 38556 20020
rect 38612 19964 38668 20076
rect 38770 19964 38780 20020
rect 38836 19964 40236 20020
rect 40292 19964 40302 20020
rect 11340 19908 11396 19964
rect 9874 19852 9884 19908
rect 9940 19852 11116 19908
rect 11172 19852 11182 19908
rect 11340 19852 25228 19908
rect 25284 19852 25294 19908
rect 27906 19852 27916 19908
rect 27972 19852 29036 19908
rect 29092 19852 30940 19908
rect 30996 19852 31006 19908
rect 35074 19852 35084 19908
rect 35140 19852 36316 19908
rect 36372 19852 36382 19908
rect 36642 19852 36652 19908
rect 36708 19852 37548 19908
rect 37604 19852 37614 19908
rect 47170 19852 47180 19908
rect 47236 19852 47628 19908
rect 47684 19852 47694 19908
rect 9986 19740 9996 19796
rect 10052 19740 10556 19796
rect 10612 19740 10622 19796
rect 18722 19740 18732 19796
rect 18788 19740 19628 19796
rect 19684 19740 19694 19796
rect 26852 19740 37100 19796
rect 37156 19740 37996 19796
rect 38052 19740 38062 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 26852 19572 26908 19740
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 21970 19516 21980 19572
rect 22036 19516 26908 19572
rect 27020 19516 30940 19572
rect 30996 19516 31006 19572
rect 36866 19516 36876 19572
rect 36932 19516 37548 19572
rect 37604 19516 37614 19572
rect 27020 19460 27076 19516
rect 15138 19404 15148 19460
rect 15204 19404 15484 19460
rect 15540 19404 27076 19460
rect 32732 19404 44492 19460
rect 44548 19404 44558 19460
rect 14998 19292 15036 19348
rect 15092 19292 15102 19348
rect 23986 19292 23996 19348
rect 24052 19292 28700 19348
rect 28756 19292 28766 19348
rect 32732 19236 32788 19404
rect 33058 19292 33068 19348
rect 33124 19292 33740 19348
rect 33796 19292 33806 19348
rect 36194 19292 36204 19348
rect 36260 19292 37212 19348
rect 37268 19292 37278 19348
rect 39554 19292 39564 19348
rect 39620 19292 40236 19348
rect 40292 19292 41020 19348
rect 41076 19292 41086 19348
rect 41570 19292 41580 19348
rect 41636 19292 42140 19348
rect 42196 19292 42206 19348
rect 10434 19180 10444 19236
rect 10500 19180 11564 19236
rect 11620 19180 12012 19236
rect 12068 19180 12078 19236
rect 25442 19180 25452 19236
rect 25508 19180 26124 19236
rect 26180 19180 32788 19236
rect 33618 19180 33628 19236
rect 33684 19180 35084 19236
rect 35140 19180 35150 19236
rect 35970 19180 35980 19236
rect 36036 19180 36316 19236
rect 36372 19180 36988 19236
rect 37044 19180 37054 19236
rect 38322 19180 38332 19236
rect 38388 19180 39676 19236
rect 39732 19180 39742 19236
rect 39890 19180 39900 19236
rect 39956 19180 40908 19236
rect 40964 19180 40974 19236
rect 44594 19180 44604 19236
rect 44660 19180 45388 19236
rect 45444 19180 45454 19236
rect 11330 19068 11340 19124
rect 11396 19068 13468 19124
rect 13524 19068 13534 19124
rect 48066 19068 48076 19124
rect 48132 19068 48142 19124
rect 11442 18956 11452 19012
rect 11508 18956 12124 19012
rect 12180 18956 12190 19012
rect 12562 18956 12572 19012
rect 12628 18956 13692 19012
rect 13748 18956 13758 19012
rect 21858 18956 21868 19012
rect 21924 18956 22204 19012
rect 22260 18956 22270 19012
rect 38182 18956 38220 19012
rect 38276 18956 38286 19012
rect 0 18816 800 18928
rect 48076 18900 48132 19068
rect 49200 18900 50000 18928
rect 23426 18844 23436 18900
rect 23492 18844 47068 18900
rect 47124 18844 47134 18900
rect 48076 18844 50000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 49200 18816 50000 18844
rect 31154 18732 31164 18788
rect 31220 18732 31948 18788
rect 32004 18732 32014 18788
rect 37538 18732 37548 18788
rect 37604 18732 38220 18788
rect 38276 18732 38286 18788
rect 10434 18620 10444 18676
rect 10500 18620 12908 18676
rect 12964 18620 27468 18676
rect 27524 18620 27534 18676
rect 31724 18620 37436 18676
rect 37492 18620 37660 18676
rect 37716 18620 37726 18676
rect 37874 18620 37884 18676
rect 37940 18620 38332 18676
rect 38388 18620 38398 18676
rect 38630 18620 38668 18676
rect 38724 18620 39228 18676
rect 39284 18620 39294 18676
rect 31724 18564 31780 18620
rect 9874 18508 9884 18564
rect 9940 18508 10836 18564
rect 10994 18508 11004 18564
rect 11060 18508 11900 18564
rect 11956 18508 11966 18564
rect 12226 18508 12236 18564
rect 12292 18508 12796 18564
rect 12852 18508 12862 18564
rect 14578 18508 14588 18564
rect 14644 18508 17164 18564
rect 17220 18508 17230 18564
rect 31714 18508 31724 18564
rect 31780 18508 31790 18564
rect 36642 18508 36652 18564
rect 36708 18508 37100 18564
rect 37156 18508 37166 18564
rect 40338 18508 40348 18564
rect 40404 18508 41692 18564
rect 41748 18508 41758 18564
rect 9202 18396 9212 18452
rect 9268 18396 9772 18452
rect 9828 18396 10332 18452
rect 10388 18396 10398 18452
rect 10780 18340 10836 18508
rect 11106 18396 11116 18452
rect 11172 18396 13244 18452
rect 13300 18396 13310 18452
rect 14354 18396 14364 18452
rect 14420 18396 14924 18452
rect 14980 18396 14990 18452
rect 17826 18396 17836 18452
rect 17892 18396 18508 18452
rect 18564 18396 18574 18452
rect 24322 18396 24332 18452
rect 24388 18396 25228 18452
rect 25284 18396 25294 18452
rect 26226 18396 26236 18452
rect 26292 18396 26796 18452
rect 26852 18396 26862 18452
rect 28802 18396 28812 18452
rect 28868 18396 36540 18452
rect 36596 18396 36606 18452
rect 38098 18396 38108 18452
rect 38164 18396 39004 18452
rect 39060 18396 39452 18452
rect 39508 18396 39518 18452
rect 12236 18340 12292 18396
rect 10780 18284 11004 18340
rect 11060 18284 11070 18340
rect 12226 18284 12236 18340
rect 12292 18284 12302 18340
rect 19170 18284 19180 18340
rect 19236 18284 20076 18340
rect 20132 18284 20524 18340
rect 20580 18284 20590 18340
rect 22642 18284 22652 18340
rect 22708 18284 25340 18340
rect 25396 18284 25406 18340
rect 27458 18284 27468 18340
rect 27524 18284 29932 18340
rect 29988 18284 29998 18340
rect 38770 18284 38780 18340
rect 38836 18284 40124 18340
rect 40180 18284 40190 18340
rect 40338 18284 40348 18340
rect 40404 18284 41804 18340
rect 41860 18284 43484 18340
rect 43540 18284 43550 18340
rect 11330 18172 11340 18228
rect 11396 18172 12460 18228
rect 12516 18172 12526 18228
rect 16258 18172 16268 18228
rect 16324 18172 16604 18228
rect 16660 18172 16670 18228
rect 37202 18172 37212 18228
rect 37268 18172 38668 18228
rect 38724 18172 38734 18228
rect 6402 18060 6412 18116
rect 6468 18060 21420 18116
rect 21476 18060 21486 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 38546 17948 38556 18004
rect 38612 17948 38668 18172
rect 30930 17836 30940 17892
rect 30996 17836 38892 17892
rect 38948 17836 38958 17892
rect 14130 17724 14140 17780
rect 14196 17724 14588 17780
rect 14644 17724 15036 17780
rect 15092 17724 15102 17780
rect 24994 17724 25004 17780
rect 25060 17724 29372 17780
rect 29428 17724 31164 17780
rect 31220 17724 31230 17780
rect 31714 17724 31724 17780
rect 31780 17724 32284 17780
rect 32340 17724 32350 17780
rect 39218 17724 39228 17780
rect 39284 17724 39676 17780
rect 39732 17724 40124 17780
rect 40180 17724 40190 17780
rect 13682 17612 13692 17668
rect 13748 17612 14476 17668
rect 14532 17612 14542 17668
rect 15092 17612 24444 17668
rect 24500 17612 25116 17668
rect 25172 17612 25564 17668
rect 25620 17612 25630 17668
rect 38770 17612 38780 17668
rect 38836 17612 39004 17668
rect 39060 17612 39452 17668
rect 39508 17612 39518 17668
rect 41570 17612 41580 17668
rect 41636 17612 42028 17668
rect 42084 17612 42094 17668
rect 13692 17556 13748 17612
rect 9538 17500 9548 17556
rect 9604 17500 11116 17556
rect 11172 17500 13748 17556
rect 14662 17500 14700 17556
rect 14756 17500 14766 17556
rect 15092 17444 15148 17612
rect 15922 17500 15932 17556
rect 15988 17500 16716 17556
rect 16772 17500 16782 17556
rect 19058 17500 19068 17556
rect 19124 17500 19964 17556
rect 20020 17500 20030 17556
rect 36194 17500 36204 17556
rect 36260 17500 37884 17556
rect 37940 17500 37950 17556
rect 5506 17388 5516 17444
rect 5572 17388 15148 17444
rect 15250 17388 15260 17444
rect 15316 17388 15820 17444
rect 15876 17388 15886 17444
rect 29922 17388 29932 17444
rect 29988 17388 30492 17444
rect 30548 17388 31164 17444
rect 31220 17388 31230 17444
rect 38322 17388 38332 17444
rect 38388 17388 38556 17444
rect 38612 17388 38622 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 26226 17052 26236 17108
rect 26292 17052 28588 17108
rect 28644 17052 28654 17108
rect 33618 17052 33628 17108
rect 33684 17052 34188 17108
rect 34244 17052 38780 17108
rect 38836 17052 38846 17108
rect 21410 16940 21420 16996
rect 21476 16940 22204 16996
rect 22260 16940 34524 16996
rect 34580 16940 34590 16996
rect 35970 16940 35980 16996
rect 36036 16940 36046 16996
rect 11666 16828 11676 16884
rect 11732 16828 12348 16884
rect 12404 16828 14140 16884
rect 14196 16828 14206 16884
rect 14466 16828 14476 16884
rect 14532 16828 15484 16884
rect 15540 16828 15708 16884
rect 15764 16828 15774 16884
rect 16258 16828 16268 16884
rect 16324 16828 18732 16884
rect 18788 16828 21084 16884
rect 21140 16828 21150 16884
rect 29362 16828 29372 16884
rect 29428 16828 29932 16884
rect 29988 16828 29998 16884
rect 31154 16828 31164 16884
rect 31220 16828 32060 16884
rect 32116 16828 32126 16884
rect 14242 16716 14252 16772
rect 14308 16716 14588 16772
rect 14644 16716 14654 16772
rect 14130 16604 14140 16660
rect 14196 16604 14700 16660
rect 14756 16604 18732 16660
rect 18788 16604 18798 16660
rect 35980 16548 36036 16940
rect 35970 16492 35980 16548
rect 36036 16492 36046 16548
rect 0 16352 800 16464
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 49200 16436 50000 16464
rect 47730 16380 47740 16436
rect 47796 16380 50000 16436
rect 49200 16352 50000 16380
rect 24658 16268 24668 16324
rect 24724 16268 25788 16324
rect 25844 16268 25854 16324
rect 14354 16156 14364 16212
rect 14420 16156 15260 16212
rect 15316 16156 15326 16212
rect 20178 16156 20188 16212
rect 20244 16156 20860 16212
rect 20916 16156 22092 16212
rect 22148 16156 23100 16212
rect 23156 16156 23166 16212
rect 24882 16156 24892 16212
rect 24948 16156 25900 16212
rect 25956 16156 25966 16212
rect 29698 16156 29708 16212
rect 29764 16156 30716 16212
rect 30772 16156 31276 16212
rect 31332 16156 31342 16212
rect 43026 16156 43036 16212
rect 43092 16156 44828 16212
rect 44884 16156 44894 16212
rect 47058 16156 47068 16212
rect 47124 16156 47628 16212
rect 47684 16156 47694 16212
rect 8978 16044 8988 16100
rect 9044 16044 10444 16100
rect 10500 16044 10510 16100
rect 19170 16044 19180 16100
rect 19236 16044 19964 16100
rect 20020 16044 21980 16100
rect 22036 16044 22046 16100
rect 29810 16044 29820 16100
rect 29876 16044 29886 16100
rect 30370 16044 30380 16100
rect 30436 16044 32060 16100
rect 32116 16044 32844 16100
rect 32900 16044 32910 16100
rect 19254 15932 19292 15988
rect 19348 15932 19358 15988
rect 10994 15820 11004 15876
rect 11060 15820 12348 15876
rect 12404 15820 12414 15876
rect 22306 15820 22316 15876
rect 22372 15820 23436 15876
rect 23492 15820 23502 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 29820 15652 29876 16044
rect 43698 15820 43708 15876
rect 43764 15820 45724 15876
rect 45780 15820 45790 15876
rect 45042 15708 45052 15764
rect 45108 15708 45500 15764
rect 45556 15708 45566 15764
rect 11330 15596 11340 15652
rect 11396 15596 12348 15652
rect 12404 15596 13132 15652
rect 13188 15596 13198 15652
rect 29810 15596 29820 15652
rect 29876 15596 29886 15652
rect 11554 15484 11564 15540
rect 11620 15484 11900 15540
rect 11956 15484 12572 15540
rect 12628 15484 12638 15540
rect 15698 15484 15708 15540
rect 15764 15484 16156 15540
rect 16212 15484 16222 15540
rect 21522 15484 21532 15540
rect 21588 15484 22316 15540
rect 22372 15484 22382 15540
rect 24434 15484 24444 15540
rect 24500 15484 25340 15540
rect 25396 15484 26908 15540
rect 27906 15484 27916 15540
rect 27972 15484 37548 15540
rect 37604 15484 37614 15540
rect 37986 15484 37996 15540
rect 38052 15484 38220 15540
rect 38276 15484 38286 15540
rect 26852 15428 26908 15484
rect 11442 15372 11452 15428
rect 11508 15372 13020 15428
rect 13076 15372 13086 15428
rect 22530 15372 22540 15428
rect 22596 15372 22876 15428
rect 22932 15372 22942 15428
rect 26852 15372 29932 15428
rect 29988 15372 38556 15428
rect 38612 15372 38622 15428
rect 23314 15260 23324 15316
rect 23380 15260 24108 15316
rect 24164 15260 24174 15316
rect 25778 15260 25788 15316
rect 25844 15260 35868 15316
rect 35924 15260 35934 15316
rect 36082 15260 36092 15316
rect 36148 15260 36764 15316
rect 36820 15260 37436 15316
rect 37492 15260 37502 15316
rect 37762 15260 37772 15316
rect 37828 15260 38780 15316
rect 38836 15260 38846 15316
rect 35868 15204 35924 15260
rect 35868 15148 36988 15204
rect 37044 15148 37054 15204
rect 26450 15092 26460 15148
rect 26516 15092 26526 15148
rect 19618 15036 19628 15092
rect 19684 15036 21196 15092
rect 21252 15036 21262 15092
rect 25890 15036 25900 15092
rect 25956 15036 26516 15092
rect 29586 15036 29596 15092
rect 29652 15036 30156 15092
rect 30212 15036 30492 15092
rect 30548 15036 30558 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 31042 14812 31052 14868
rect 31108 14812 35028 14868
rect 34972 14756 35028 14812
rect 30482 14700 30492 14756
rect 30548 14700 32060 14756
rect 32116 14700 32126 14756
rect 34972 14700 46732 14756
rect 46788 14700 46798 14756
rect 14466 14588 14476 14644
rect 14532 14588 14700 14644
rect 14756 14588 15708 14644
rect 15764 14588 15774 14644
rect 16706 14588 16716 14644
rect 16772 14588 21588 14644
rect 28914 14588 28924 14644
rect 28980 14588 29260 14644
rect 29316 14588 29708 14644
rect 29764 14588 29774 14644
rect 30594 14588 30604 14644
rect 30660 14588 31052 14644
rect 31108 14588 31118 14644
rect 31892 14588 33292 14644
rect 33348 14588 35868 14644
rect 35924 14588 38332 14644
rect 38388 14588 38398 14644
rect 40450 14588 40460 14644
rect 40516 14588 40908 14644
rect 40964 14588 40974 14644
rect 43586 14588 43596 14644
rect 43652 14588 44828 14644
rect 44884 14588 44894 14644
rect 21532 14532 21588 14588
rect 31892 14532 31948 14588
rect 12562 14476 12572 14532
rect 12628 14476 17836 14532
rect 17892 14476 17902 14532
rect 21522 14476 21532 14532
rect 21588 14476 23548 14532
rect 23604 14476 23614 14532
rect 25554 14476 25564 14532
rect 25620 14476 31948 14532
rect 36866 14476 36876 14532
rect 36932 14476 37212 14532
rect 37268 14476 37278 14532
rect 39106 14476 39116 14532
rect 39172 14476 40124 14532
rect 40180 14476 41132 14532
rect 41188 14476 41198 14532
rect 43474 14476 43484 14532
rect 43540 14476 44044 14532
rect 44100 14476 44110 14532
rect 44258 14476 44268 14532
rect 44324 14476 45388 14532
rect 45444 14476 45454 14532
rect 13570 14364 13580 14420
rect 13636 14364 14588 14420
rect 14644 14364 14654 14420
rect 15362 14364 15372 14420
rect 15428 14364 16604 14420
rect 16660 14364 16670 14420
rect 17042 14364 17052 14420
rect 17108 14364 22652 14420
rect 22708 14364 22718 14420
rect 25666 14364 25676 14420
rect 25732 14364 26572 14420
rect 26628 14364 26638 14420
rect 26898 14364 26908 14420
rect 26964 14364 32732 14420
rect 32788 14364 35420 14420
rect 35476 14364 38220 14420
rect 38276 14364 38286 14420
rect 11890 14252 11900 14308
rect 11956 14252 13020 14308
rect 13076 14252 17388 14308
rect 17444 14252 17454 14308
rect 22082 14252 22092 14308
rect 22148 14252 24668 14308
rect 24724 14252 32396 14308
rect 32452 14252 32462 14308
rect 35522 14252 35532 14308
rect 35588 14252 36876 14308
rect 36932 14252 36942 14308
rect 13804 14084 13860 14252
rect 31892 14140 36092 14196
rect 36148 14140 37100 14196
rect 37156 14140 37166 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 31892 14084 31948 14140
rect 13794 14028 13804 14084
rect 13860 14028 13870 14084
rect 29138 14028 29148 14084
rect 29204 14028 31948 14084
rect 0 13888 800 14000
rect 49200 13972 50000 14000
rect 12898 13916 12908 13972
rect 12964 13916 16716 13972
rect 16772 13916 16782 13972
rect 18722 13916 18732 13972
rect 18788 13916 19628 13972
rect 19684 13916 19694 13972
rect 31052 13916 31836 13972
rect 31892 13916 32284 13972
rect 32340 13916 32350 13972
rect 37426 13916 37436 13972
rect 37492 13916 38220 13972
rect 38276 13916 38286 13972
rect 48066 13916 48076 13972
rect 48132 13916 50000 13972
rect 31052 13860 31108 13916
rect 49200 13888 50000 13916
rect 13346 13804 13356 13860
rect 13412 13804 14476 13860
rect 14532 13804 14542 13860
rect 15138 13804 15148 13860
rect 15204 13804 15484 13860
rect 15540 13804 15550 13860
rect 23986 13804 23996 13860
rect 24052 13804 25228 13860
rect 25284 13804 25294 13860
rect 30482 13804 30492 13860
rect 30548 13804 31052 13860
rect 31108 13804 31118 13860
rect 37538 13804 37548 13860
rect 37604 13804 38108 13860
rect 38164 13804 38174 13860
rect 43922 13804 43932 13860
rect 43988 13804 46620 13860
rect 46676 13804 46686 13860
rect 20626 13692 20636 13748
rect 20692 13692 22204 13748
rect 22260 13692 22270 13748
rect 23426 13692 23436 13748
rect 23492 13692 24108 13748
rect 24164 13692 24556 13748
rect 24612 13692 24622 13748
rect 38770 13692 38780 13748
rect 38836 13692 39452 13748
rect 39508 13692 39518 13748
rect 12338 13580 12348 13636
rect 12404 13580 13468 13636
rect 13524 13580 13534 13636
rect 15922 13580 15932 13636
rect 15988 13580 21084 13636
rect 21140 13580 21756 13636
rect 21812 13580 21822 13636
rect 26852 13580 27132 13636
rect 27188 13580 27198 13636
rect 38434 13580 38444 13636
rect 38500 13580 39060 13636
rect 26852 13524 26908 13580
rect 39004 13524 39060 13580
rect 14438 13468 14476 13524
rect 14532 13468 14542 13524
rect 17602 13468 17612 13524
rect 17668 13468 19292 13524
rect 19348 13468 19358 13524
rect 23426 13468 23436 13524
rect 23492 13468 26908 13524
rect 38994 13468 39004 13524
rect 39060 13468 39900 13524
rect 39956 13468 39966 13524
rect 14354 13356 14364 13412
rect 14420 13356 15820 13412
rect 15876 13356 15886 13412
rect 36194 13356 36204 13412
rect 36260 13356 36652 13412
rect 36708 13356 37100 13412
rect 37156 13356 38668 13412
rect 38724 13356 38734 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 15586 13244 15596 13300
rect 15652 13244 15932 13300
rect 15988 13244 15998 13300
rect 14914 13020 14924 13076
rect 14980 13020 15932 13076
rect 15988 13020 15998 13076
rect 19618 13020 19628 13076
rect 19684 13020 20076 13076
rect 20132 13020 20412 13076
rect 20468 13020 20524 13076
rect 20580 13020 20590 13076
rect 43250 13020 43260 13076
rect 43316 13020 45052 13076
rect 45108 13020 45118 13076
rect 12226 12908 12236 12964
rect 12292 12908 12796 12964
rect 12852 12908 13692 12964
rect 13748 12908 13758 12964
rect 30818 12908 30828 12964
rect 30884 12908 32060 12964
rect 32116 12908 32126 12964
rect 39330 12908 39340 12964
rect 39396 12908 39788 12964
rect 39844 12908 39854 12964
rect 13570 12796 13580 12852
rect 13636 12796 14028 12852
rect 14084 12796 15372 12852
rect 15428 12796 15438 12852
rect 19058 12796 19068 12852
rect 19124 12796 19628 12852
rect 19684 12796 19694 12852
rect 39890 12796 39900 12852
rect 39956 12796 41692 12852
rect 41748 12796 42252 12852
rect 42308 12796 42318 12852
rect 18610 12684 18620 12740
rect 18676 12684 19740 12740
rect 19796 12684 19806 12740
rect 22530 12684 22540 12740
rect 22596 12684 25340 12740
rect 25396 12684 26908 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 26852 12404 26908 12684
rect 12674 12348 12684 12404
rect 12740 12348 13356 12404
rect 13412 12348 13422 12404
rect 15362 12348 15372 12404
rect 15428 12348 16604 12404
rect 16660 12348 16670 12404
rect 25442 12348 25452 12404
rect 25508 12348 26348 12404
rect 26404 12348 26414 12404
rect 26852 12348 28252 12404
rect 28308 12348 28318 12404
rect 27794 12236 27804 12292
rect 27860 12236 35532 12292
rect 35588 12236 35598 12292
rect 15138 12124 15148 12180
rect 15204 12124 15820 12180
rect 15876 12124 15886 12180
rect 26226 12124 26236 12180
rect 26292 12124 27468 12180
rect 27524 12124 27534 12180
rect 28466 12124 28476 12180
rect 28532 12124 46732 12180
rect 46788 12124 46798 12180
rect 13682 12012 13692 12068
rect 13748 12012 14252 12068
rect 14308 12012 14318 12068
rect 41458 12012 41468 12068
rect 41524 12012 42364 12068
rect 42420 12012 42430 12068
rect 19068 11900 19292 11956
rect 19348 11900 19358 11956
rect 38770 11900 38780 11956
rect 38836 11900 41692 11956
rect 41748 11900 42588 11956
rect 42644 11900 42654 11956
rect 19068 11844 19124 11900
rect 12226 11788 12236 11844
rect 12292 11788 13916 11844
rect 13972 11788 13982 11844
rect 15026 11788 15036 11844
rect 15092 11788 15596 11844
rect 15652 11788 15662 11844
rect 19058 11788 19068 11844
rect 19124 11788 19134 11844
rect 23762 11788 23772 11844
rect 23828 11788 25004 11844
rect 25060 11788 26236 11844
rect 26292 11788 26302 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 11218 11676 11228 11732
rect 11284 11676 12348 11732
rect 12404 11676 13020 11732
rect 13076 11676 13086 11732
rect 22754 11676 22764 11732
rect 22820 11676 23660 11732
rect 23716 11676 23726 11732
rect 0 11424 800 11536
rect 49200 11508 50000 11536
rect 29138 11452 29148 11508
rect 29204 11452 29820 11508
rect 29876 11452 29886 11508
rect 33282 11452 33292 11508
rect 33348 11452 34188 11508
rect 34244 11452 34254 11508
rect 47730 11452 47740 11508
rect 47796 11452 50000 11508
rect 49200 11424 50000 11452
rect 28242 11340 28252 11396
rect 28308 11340 31948 11396
rect 32946 11340 32956 11396
rect 33012 11340 33740 11396
rect 33796 11340 33806 11396
rect 36306 11340 36316 11396
rect 36372 11340 37324 11396
rect 37380 11340 38220 11396
rect 38276 11340 38286 11396
rect 31892 11284 31948 11340
rect 11330 11228 11340 11284
rect 11396 11228 12460 11284
rect 12516 11228 12526 11284
rect 28018 11228 28028 11284
rect 28084 11228 28588 11284
rect 28644 11228 28654 11284
rect 29250 11228 29260 11284
rect 29316 11228 30268 11284
rect 30324 11228 30334 11284
rect 31892 11228 36204 11284
rect 36260 11228 36270 11284
rect 29260 11172 29316 11228
rect 12786 11116 12796 11172
rect 12852 11116 18172 11172
rect 18228 11116 18956 11172
rect 19012 11116 19022 11172
rect 24546 11116 24556 11172
rect 24612 11116 25116 11172
rect 25172 11116 29316 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 24770 10780 24780 10836
rect 24836 10780 26012 10836
rect 26068 10780 26078 10836
rect 21522 10668 21532 10724
rect 21588 10668 22764 10724
rect 22820 10668 22830 10724
rect 34962 10668 34972 10724
rect 35028 10668 35644 10724
rect 35700 10668 35710 10724
rect 43474 10668 43484 10724
rect 43540 10668 44380 10724
rect 44436 10668 44446 10724
rect 18610 10556 18620 10612
rect 18676 10556 19628 10612
rect 19684 10556 19694 10612
rect 20066 10556 20076 10612
rect 20132 10556 20748 10612
rect 20804 10556 21868 10612
rect 21924 10556 21934 10612
rect 35522 10556 35532 10612
rect 35588 10556 37548 10612
rect 37604 10556 37614 10612
rect 43250 10556 43260 10612
rect 43316 10556 44044 10612
rect 44100 10556 44110 10612
rect 34178 10444 34188 10500
rect 34244 10444 34972 10500
rect 35028 10444 35420 10500
rect 35476 10444 36764 10500
rect 36820 10444 36830 10500
rect 27010 10332 27020 10388
rect 27076 10332 27692 10388
rect 27748 10332 27758 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 26450 10108 26460 10164
rect 26516 10108 27356 10164
rect 27412 10108 27422 10164
rect 42802 10108 42812 10164
rect 42868 10108 44044 10164
rect 44100 10108 44110 10164
rect 13234 9996 13244 10052
rect 13300 9996 15708 10052
rect 15764 9996 16604 10052
rect 16660 9996 16670 10052
rect 29474 9996 29484 10052
rect 29540 9996 30716 10052
rect 30772 9996 30782 10052
rect 15810 9884 15820 9940
rect 15876 9884 16268 9940
rect 16324 9884 17164 9940
rect 17220 9884 25564 9940
rect 25620 9884 25630 9940
rect 33618 9884 33628 9940
rect 33684 9884 46732 9940
rect 46788 9884 46798 9940
rect 12002 9772 12012 9828
rect 12068 9772 15596 9828
rect 15652 9772 15662 9828
rect 19170 9772 19180 9828
rect 19236 9772 20188 9828
rect 20244 9772 20254 9828
rect 37986 9772 37996 9828
rect 38052 9772 38668 9828
rect 38724 9772 38734 9828
rect 42130 9772 42140 9828
rect 42196 9772 42924 9828
rect 42980 9772 42990 9828
rect 18722 9660 18732 9716
rect 18788 9660 19628 9716
rect 19684 9660 19694 9716
rect 20850 9660 20860 9716
rect 20916 9660 21644 9716
rect 21700 9660 21710 9716
rect 27010 9660 27020 9716
rect 27076 9660 27580 9716
rect 27636 9660 37436 9716
rect 37492 9660 37772 9716
rect 37828 9660 38108 9716
rect 38164 9660 38174 9716
rect 38322 9660 38332 9716
rect 38388 9660 39340 9716
rect 39396 9660 39406 9716
rect 14354 9548 14364 9604
rect 14420 9548 17724 9604
rect 17780 9548 18396 9604
rect 18452 9548 18462 9604
rect 40114 9548 40124 9604
rect 40180 9548 40908 9604
rect 40964 9548 40974 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 37650 9212 37660 9268
rect 37716 9212 38668 9268
rect 38724 9212 38734 9268
rect 13906 9100 13916 9156
rect 13972 9100 14924 9156
rect 14980 9100 14990 9156
rect 31154 9100 31164 9156
rect 31220 9100 31724 9156
rect 31780 9100 31790 9156
rect 0 8960 800 9072
rect 49200 9044 50000 9072
rect 28466 8988 28476 9044
rect 28532 8988 33516 9044
rect 33572 8988 33582 9044
rect 36530 8988 36540 9044
rect 36596 8988 37212 9044
rect 37268 8988 38444 9044
rect 38500 8988 38510 9044
rect 43362 8988 43372 9044
rect 43428 8988 44044 9044
rect 44100 8988 44110 9044
rect 48066 8988 48076 9044
rect 48132 8988 50000 9044
rect 49200 8960 50000 8988
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 34514 8428 34524 8484
rect 34580 8428 35084 8484
rect 35140 8428 35150 8484
rect 15474 8316 15484 8372
rect 15540 8316 16492 8372
rect 16548 8316 17948 8372
rect 18004 8316 18014 8372
rect 21746 8316 21756 8372
rect 21812 8316 22428 8372
rect 22484 8316 22494 8372
rect 15698 8204 15708 8260
rect 15764 8204 16604 8260
rect 16660 8204 17724 8260
rect 17780 8204 17790 8260
rect 22306 8204 22316 8260
rect 22372 8204 23772 8260
rect 23828 8204 23838 8260
rect 34402 8204 34412 8260
rect 34468 8204 35084 8260
rect 35140 8204 35150 8260
rect 17378 8092 17388 8148
rect 17444 8092 18620 8148
rect 18676 8092 18686 8148
rect 19506 8092 19516 8148
rect 19572 8092 20412 8148
rect 20468 8092 20478 8148
rect 31892 8092 41132 8148
rect 41188 8092 41198 8148
rect 31892 8036 31948 8092
rect 20066 7980 20076 8036
rect 20132 7980 20636 8036
rect 20692 7980 20702 8036
rect 22866 7980 22876 8036
rect 22932 7980 23660 8036
rect 23716 7980 23726 8036
rect 27906 7980 27916 8036
rect 27972 7980 31948 8036
rect 33394 7980 33404 8036
rect 33460 7980 34636 8036
rect 34692 7980 34702 8036
rect 26898 7868 26908 7924
rect 26964 7868 27468 7924
rect 27524 7868 28252 7924
rect 28308 7868 28318 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 26226 7756 26236 7812
rect 26292 7756 27132 7812
rect 27188 7756 27804 7812
rect 27860 7756 27870 7812
rect 28018 7644 28028 7700
rect 28084 7644 28700 7700
rect 28756 7644 28766 7700
rect 20962 7532 20972 7588
rect 21028 7532 21868 7588
rect 21924 7532 21934 7588
rect 24098 7420 24108 7476
rect 24164 7420 25788 7476
rect 25844 7420 25854 7476
rect 31602 7420 31612 7476
rect 31668 7420 32956 7476
rect 33012 7420 33022 7476
rect 34962 7420 34972 7476
rect 35028 7420 35532 7476
rect 35588 7420 35598 7476
rect 41906 7420 41916 7476
rect 41972 7420 42476 7476
rect 42532 7420 42542 7476
rect 41458 7196 41468 7252
rect 41524 7196 42812 7252
rect 42868 7196 42878 7252
rect 29810 7084 29820 7140
rect 29876 7084 30268 7140
rect 30324 7084 30334 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 24322 6860 24332 6916
rect 24388 6860 25228 6916
rect 25284 6860 25294 6916
rect 26898 6860 26908 6916
rect 26964 6860 27356 6916
rect 27412 6860 27422 6916
rect 36082 6748 36092 6804
rect 36148 6748 36764 6804
rect 36820 6748 36830 6804
rect 37762 6748 37772 6804
rect 37828 6748 38780 6804
rect 38836 6748 38846 6804
rect 31266 6636 31276 6692
rect 31332 6636 32396 6692
rect 32452 6636 34412 6692
rect 34468 6636 34478 6692
rect 0 6496 800 6608
rect 49200 6580 50000 6608
rect 31378 6524 31388 6580
rect 31444 6524 33180 6580
rect 33236 6524 33852 6580
rect 33908 6524 34636 6580
rect 34692 6524 34702 6580
rect 48066 6524 48076 6580
rect 48132 6524 50000 6580
rect 49200 6496 50000 6524
rect 31892 6412 35420 6468
rect 35476 6412 35486 6468
rect 31892 6356 31948 6412
rect 29810 6300 29820 6356
rect 29876 6300 30380 6356
rect 30436 6300 31948 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 18834 6076 18844 6132
rect 18900 6076 20300 6132
rect 20356 6076 20366 6132
rect 26562 6076 26572 6132
rect 26628 6076 33180 6132
rect 33236 6076 33852 6132
rect 33908 6076 36428 6132
rect 36484 6076 37324 6132
rect 37380 6076 37884 6132
rect 37940 6076 37950 6132
rect 38882 6076 38892 6132
rect 38948 6076 39564 6132
rect 39620 6076 39630 6132
rect 18386 5964 18396 6020
rect 18452 5964 19180 6020
rect 19236 5964 19246 6020
rect 33628 5964 37548 6020
rect 37604 5964 37614 6020
rect 40898 5964 40908 6020
rect 40964 5964 41580 6020
rect 41636 5964 42364 6020
rect 42420 5964 42430 6020
rect 33628 5908 33684 5964
rect 13458 5852 13468 5908
rect 13524 5852 14364 5908
rect 14420 5852 14430 5908
rect 16258 5852 16268 5908
rect 16324 5852 16716 5908
rect 16772 5852 17724 5908
rect 17780 5852 17790 5908
rect 19058 5852 19068 5908
rect 19124 5852 19852 5908
rect 19908 5852 20860 5908
rect 20916 5852 20926 5908
rect 24546 5852 24556 5908
rect 24612 5852 33628 5908
rect 33684 5852 33694 5908
rect 35522 5852 35532 5908
rect 35588 5852 36092 5908
rect 36148 5852 36158 5908
rect 15026 5740 15036 5796
rect 15092 5740 15708 5796
rect 15764 5740 15774 5796
rect 35634 5740 35644 5796
rect 35700 5740 37436 5796
rect 37492 5740 37996 5796
rect 38052 5740 38062 5796
rect 14578 5628 14588 5684
rect 14644 5628 17276 5684
rect 17332 5628 17342 5684
rect 20290 5628 20300 5684
rect 20356 5628 22316 5684
rect 22372 5628 22382 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19394 5292 19404 5348
rect 19460 5292 20524 5348
rect 20580 5292 20590 5348
rect 24994 5292 25004 5348
rect 25060 5292 28700 5348
rect 28756 5292 31948 5348
rect 17938 5180 17948 5236
rect 18004 5180 24332 5236
rect 24388 5180 24398 5236
rect 25330 5180 25340 5236
rect 25396 5180 26012 5236
rect 26068 5180 26078 5236
rect 20738 5068 20748 5124
rect 20804 5068 21532 5124
rect 21588 5068 22316 5124
rect 22372 5068 22382 5124
rect 22642 5068 22652 5124
rect 22708 5068 23828 5124
rect 29362 5068 29372 5124
rect 29428 5068 30044 5124
rect 30100 5068 30604 5124
rect 30660 5068 30670 5124
rect 23772 5012 23828 5068
rect 31892 5012 31948 5292
rect 37884 5068 39284 5124
rect 37884 5012 37940 5068
rect 39228 5012 39284 5068
rect 23762 4956 23772 5012
rect 23828 4956 25340 5012
rect 25396 4956 25406 5012
rect 31892 4956 37940 5012
rect 38098 4956 38108 5012
rect 38164 4956 39004 5012
rect 39060 4956 39070 5012
rect 39228 4956 41132 5012
rect 41188 4956 41198 5012
rect 28018 4844 28028 4900
rect 28084 4844 39452 4900
rect 39508 4844 40460 4900
rect 40516 4844 40526 4900
rect 40226 4732 40236 4788
rect 40292 4732 44604 4788
rect 44660 4732 44670 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 28466 4508 28476 4564
rect 28532 4508 31948 4564
rect 31892 4452 31948 4508
rect 14690 4396 14700 4452
rect 14756 4396 19012 4452
rect 29922 4396 29932 4452
rect 29988 4396 30492 4452
rect 30548 4396 30558 4452
rect 31892 4396 46620 4452
rect 46676 4396 46686 4452
rect 11330 4172 11340 4228
rect 11396 4172 13468 4228
rect 13524 4172 13534 4228
rect 0 4032 800 4144
rect 18956 4116 19012 4396
rect 23538 4284 23548 4340
rect 23604 4284 25900 4340
rect 25956 4284 25966 4340
rect 27458 4284 27468 4340
rect 27524 4284 30604 4340
rect 30660 4284 31500 4340
rect 31556 4284 31566 4340
rect 49200 4116 50000 4144
rect 18946 4060 18956 4116
rect 19012 4060 19404 4116
rect 19460 4060 45276 4116
rect 45332 4060 45342 4116
rect 48066 4060 48076 4116
rect 48132 4060 50000 4116
rect 49200 4032 50000 4060
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 22978 3612 22988 3668
rect 23044 3612 24892 3668
rect 24948 3612 24958 3668
rect 40674 3612 40684 3668
rect 40740 3612 44044 3668
rect 44100 3612 44110 3668
rect 26898 3500 26908 3556
rect 26964 3500 46060 3556
rect 46116 3500 46126 3556
rect 7298 3388 7308 3444
rect 7364 3388 8764 3444
rect 8820 3388 8830 3444
rect 14802 3388 14812 3444
rect 14868 3388 15372 3444
rect 15428 3388 15438 3444
rect 21522 3388 21532 3444
rect 21588 3388 31220 3444
rect 31164 3332 31220 3388
rect 31154 3276 31164 3332
rect 31220 3276 31230 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 1568 800 1680
rect 49200 1652 50000 1680
rect 47730 1596 47740 1652
rect 47796 1596 50000 1652
rect 49200 1568 50000 1596
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 22092 76300 22148 76356
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 7084 69132 7140 69188
rect 34972 69132 35028 69188
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 7644 67900 7700 67956
rect 19292 67564 19348 67620
rect 31388 67564 31444 67620
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 12236 66108 12292 66164
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 15484 64428 15540 64484
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 12236 64092 12292 64148
rect 19068 63644 19124 63700
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 7196 63084 7252 63140
rect 7644 63084 7700 63140
rect 33404 62972 33460 63028
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 7196 62300 7252 62356
rect 31724 62300 31780 62356
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 18956 61516 19012 61572
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 19068 61068 19124 61124
rect 33404 60508 33460 60564
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19292 60060 19348 60116
rect 18956 59948 19012 60004
rect 31388 59612 31444 59668
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 15484 59052 15540 59108
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 9212 58604 9268 58660
rect 37996 58156 38052 58212
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 10668 57932 10724 57988
rect 15260 57932 15316 57988
rect 17948 57932 18004 57988
rect 11452 57708 11508 57764
rect 10780 57596 10836 57652
rect 15708 57596 15764 57652
rect 44604 57596 44660 57652
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 8988 57148 9044 57204
rect 15932 57036 15988 57092
rect 40796 56812 40852 56868
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 23324 56364 23380 56420
rect 28476 56252 28532 56308
rect 13804 56028 13860 56084
rect 41020 55916 41076 55972
rect 44604 55916 44660 55972
rect 18732 55804 18788 55860
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 25676 55356 25732 55412
rect 22316 55244 22372 55300
rect 25452 55244 25508 55300
rect 33404 54908 33460 54964
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 14476 54796 14532 54852
rect 41692 54684 41748 54740
rect 13804 54572 13860 54628
rect 16156 54572 16212 54628
rect 39228 54236 39284 54292
rect 41244 54124 41300 54180
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 28140 54012 28196 54068
rect 6076 53900 6132 53956
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 13804 53004 13860 53060
rect 10668 52892 10724 52948
rect 22652 52892 22708 52948
rect 40908 52892 40964 52948
rect 41244 52780 41300 52836
rect 15260 52668 15316 52724
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 41132 52332 41188 52388
rect 41692 52332 41748 52388
rect 16156 52220 16212 52276
rect 15708 51996 15764 52052
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 23324 51324 23380 51380
rect 40796 51660 40852 51716
rect 28812 51100 28868 51156
rect 40908 51100 40964 51156
rect 18732 50988 18788 51044
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 35756 50876 35812 50932
rect 41580 50764 41636 50820
rect 28140 50652 28196 50708
rect 6076 50540 6132 50596
rect 37660 50540 37716 50596
rect 10780 50204 10836 50260
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 11452 49980 11508 50036
rect 17948 49980 18004 50036
rect 25452 49980 25508 50036
rect 22316 49868 22372 49924
rect 10780 49644 10836 49700
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 15932 49308 15988 49364
rect 9212 48972 9268 49028
rect 26684 48972 26740 49028
rect 33404 48748 33460 48804
rect 39228 48748 39284 48804
rect 14476 48636 14532 48692
rect 35756 48636 35812 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 41132 48524 41188 48580
rect 7084 48412 7140 48468
rect 8988 48188 9044 48244
rect 41020 48076 41076 48132
rect 10780 47964 10836 48020
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 25676 47516 25732 47572
rect 7644 47180 7700 47236
rect 26796 47180 26852 47236
rect 22652 47068 22708 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 26572 46844 26628 46900
rect 34748 46620 34804 46676
rect 26684 46396 26740 46452
rect 34636 46396 34692 46452
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 37548 46172 37604 46228
rect 22764 45948 22820 46004
rect 26796 45948 26852 46004
rect 21532 45612 21588 45668
rect 29260 45612 29316 45668
rect 41916 45612 41972 45668
rect 29036 45500 29092 45556
rect 41244 45500 41300 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 24668 45388 24724 45444
rect 38668 45388 38724 45444
rect 19404 45276 19460 45332
rect 30940 45276 30996 45332
rect 7980 44940 8036 44996
rect 29708 44828 29764 44884
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 22316 44604 22372 44660
rect 3948 44380 4004 44436
rect 41244 44268 41300 44324
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 18956 43820 19012 43876
rect 30940 43820 30996 43876
rect 22764 43596 22820 43652
rect 30044 43596 30100 43652
rect 38668 43260 38724 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 6972 43036 7028 43092
rect 41244 42812 41300 42868
rect 41916 42812 41972 42868
rect 7308 42588 7364 42644
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 8988 41804 9044 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 36092 41244 36148 41300
rect 18956 41132 19012 41188
rect 6972 41020 7028 41076
rect 7420 41020 7476 41076
rect 22428 41020 22484 41076
rect 7084 40796 7140 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 28700 40572 28756 40628
rect 8204 40012 8260 40068
rect 28700 40012 28756 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 21532 39900 21588 39956
rect 22428 39788 22484 39844
rect 40236 39564 40292 39620
rect 7084 39340 7140 39396
rect 34636 39228 34692 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 8092 38892 8148 38948
rect 7308 38780 7364 38836
rect 7980 38780 8036 38836
rect 36092 38444 36148 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 8092 38332 8148 38388
rect 29036 38332 29092 38388
rect 8204 38220 8260 38276
rect 29260 38220 29316 38276
rect 24668 37996 24724 38052
rect 3948 37772 4004 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 19404 37324 19460 37380
rect 34748 37324 34804 37380
rect 37548 37324 37604 37380
rect 26572 36988 26628 37044
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 22316 36540 22372 36596
rect 41244 36428 41300 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 18844 35868 18900 35924
rect 30044 35420 30100 35476
rect 8988 35308 9044 35364
rect 29708 35308 29764 35364
rect 34972 35308 35028 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 7420 34636 7476 34692
rect 37100 34636 37156 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 14700 34300 14756 34356
rect 46284 34524 46340 34580
rect 18844 34188 18900 34244
rect 2716 33964 2772 34020
rect 46508 34076 46564 34132
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 18732 33628 18788 33684
rect 31052 33628 31108 33684
rect 21980 33180 22036 33236
rect 17836 33068 17892 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 7644 32844 7700 32900
rect 22092 32732 22148 32788
rect 12572 32508 12628 32564
rect 34748 32508 34804 32564
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 2716 32060 2772 32116
rect 14252 32060 14308 32116
rect 31724 31836 31780 31892
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 15036 31276 15092 31332
rect 31724 31276 31780 31332
rect 5516 30604 5572 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 44380 30380 44436 30436
rect 14364 30156 14420 30212
rect 11452 29932 11508 29988
rect 15036 29932 15092 29988
rect 29596 29820 29652 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 29708 29596 29764 29652
rect 5516 29484 5572 29540
rect 14364 29372 14420 29428
rect 40236 29260 40292 29316
rect 11452 29148 11508 29204
rect 39004 29148 39060 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 37100 28588 37156 28644
rect 14700 28476 14756 28532
rect 27020 28364 27076 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 14028 28140 14084 28196
rect 39004 28028 39060 28084
rect 23436 27916 23492 27972
rect 21980 27804 22036 27860
rect 11788 27580 11844 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 37660 27244 37716 27300
rect 46284 27244 46340 27300
rect 17836 27020 17892 27076
rect 12572 26796 12628 26852
rect 31724 26796 31780 26852
rect 27020 26684 27076 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 34748 26572 34804 26628
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 18732 25788 18788 25844
rect 14364 25452 14420 25508
rect 46508 25340 46564 25396
rect 14252 25228 14308 25284
rect 15036 25116 15092 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 37996 25004 38052 25060
rect 11788 24892 11844 24948
rect 23436 24556 23492 24612
rect 29708 24556 29764 24612
rect 14028 24332 14084 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 12572 23996 12628 24052
rect 44380 23996 44436 24052
rect 29596 23660 29652 23716
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 37436 23436 37492 23492
rect 41580 23436 41636 23492
rect 16156 23212 16212 23268
rect 38668 22764 38724 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 15036 22652 15092 22708
rect 39452 22540 39508 22596
rect 20524 22316 20580 22372
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 14700 21868 14756 21924
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 28812 20972 28868 21028
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 30940 19516 30996 19572
rect 15036 19292 15092 19348
rect 38220 18956 38276 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 38668 18620 38724 18676
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 39452 17612 39508 17668
rect 14700 17500 14756 17556
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19292 15932 19348 15988
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 16156 15484 16212 15540
rect 38220 15484 38276 15540
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 31052 14812 31108 14868
rect 14476 14588 14532 14644
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 37436 13916 37492 13972
rect 14476 13468 14532 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 20524 13020 20580 13076
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 19292 11900 19348 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 28476 4508 28532 4564
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 7084 69188 7140 69198
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 6076 53956 6132 53966
rect 6076 50596 6132 53900
rect 6076 50530 6132 50540
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 7084 48468 7140 69132
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 7644 67956 7700 67966
rect 7196 63140 7252 63150
rect 7196 62356 7252 63084
rect 7644 63140 7700 67900
rect 19292 67620 19348 67630
rect 12236 66164 12292 66174
rect 12236 64148 12292 66108
rect 12236 64082 12292 64092
rect 15484 64484 15540 64494
rect 7644 63074 7700 63084
rect 7196 62290 7252 62300
rect 15484 59108 15540 64428
rect 19068 63700 19124 63710
rect 18956 61572 19012 61582
rect 18956 60004 19012 61516
rect 19068 61124 19124 63644
rect 19068 61058 19124 61068
rect 19292 60116 19348 67564
rect 19292 60050 19348 60060
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 18956 59938 19012 59948
rect 15484 59042 15540 59052
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 9212 58660 9268 58670
rect 7084 48402 7140 48412
rect 8988 57204 9044 57214
rect 8988 48244 9044 57148
rect 9212 49028 9268 58604
rect 19808 58044 20128 59556
rect 10668 57988 10724 57998
rect 10668 52948 10724 57932
rect 15260 57988 15316 57998
rect 11452 57764 11508 57774
rect 10668 52882 10724 52892
rect 10780 57652 10836 57662
rect 10780 50260 10836 57596
rect 10780 50194 10836 50204
rect 11452 50036 11508 57708
rect 13804 56084 13860 56094
rect 13804 54628 13860 56028
rect 13804 53060 13860 54572
rect 13804 52994 13860 53004
rect 14476 54852 14532 54862
rect 11452 49970 11508 49980
rect 9212 48962 9268 48972
rect 10780 49700 10836 49710
rect 8988 48178 9044 48188
rect 10780 48020 10836 49644
rect 14476 48692 14532 54796
rect 15260 52724 15316 57932
rect 17948 57988 18004 57998
rect 15260 52658 15316 52668
rect 15708 57652 15764 57662
rect 15708 52052 15764 57596
rect 15708 51986 15764 51996
rect 15932 57092 15988 57102
rect 15932 49364 15988 57036
rect 16156 54628 16212 54638
rect 16156 52276 16212 54572
rect 16156 52210 16212 52220
rect 17948 50036 18004 57932
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 18732 55860 18788 55870
rect 18732 51044 18788 55804
rect 18732 50978 18788 50988
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 17948 49970 18004 49980
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 15932 49298 15988 49308
rect 14476 48626 14532 48636
rect 19808 48636 20128 50148
rect 10780 47954 10836 47964
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 3948 44436 4004 44446
rect 3948 37828 4004 44380
rect 3948 37762 4004 37772
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 7644 47236 7700 47246
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 6972 43092 7028 43102
rect 6972 41076 7028 43036
rect 6972 41010 7028 41020
rect 7308 42644 7364 42654
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 7084 40852 7140 40862
rect 7084 39396 7140 40796
rect 7084 39330 7140 39340
rect 7308 38836 7364 42588
rect 7308 38770 7364 38780
rect 7420 41076 7476 41086
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 2716 34020 2772 34030
rect 2716 32116 2772 33964
rect 2716 32050 2772 32060
rect 4448 33740 4768 35252
rect 7420 34692 7476 41020
rect 7420 34626 7476 34636
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 7644 32900 7700 47180
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 22092 76356 22148 76366
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19404 45332 19460 45342
rect 7980 44996 8036 45006
rect 7980 38836 8036 44940
rect 18956 43876 19012 43886
rect 8988 41860 9044 41870
rect 8204 40068 8260 40078
rect 7980 38770 8036 38780
rect 8092 38948 8148 38958
rect 8092 38388 8148 38892
rect 8092 38322 8148 38332
rect 8204 38276 8260 40012
rect 8204 38210 8260 38220
rect 8988 35364 9044 41804
rect 18956 41188 19012 43820
rect 18956 41122 19012 41132
rect 19404 37380 19460 45276
rect 19404 37314 19460 37324
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 21532 45668 21588 45678
rect 21532 39956 21588 45612
rect 21532 39890 21588 39900
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 8988 35298 9044 35308
rect 18844 35924 18900 35934
rect 7644 32834 7700 32844
rect 14700 34356 14756 34366
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 12572 32564 12628 32574
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 5516 30660 5572 30670
rect 5516 29540 5572 30604
rect 5516 29474 5572 29484
rect 11452 29988 11508 29998
rect 11452 29204 11508 29932
rect 11452 29138 11508 29148
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 11788 27636 11844 27646
rect 11788 24948 11844 27580
rect 11788 24882 11844 24892
rect 12572 26852 12628 32508
rect 14252 32116 14308 32126
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 12572 24052 12628 26796
rect 14028 28196 14084 28206
rect 14028 24388 14084 28140
rect 14252 25284 14308 32060
rect 14364 30212 14420 30222
rect 14364 29428 14420 30156
rect 14364 25508 14420 29372
rect 14700 28532 14756 34300
rect 18844 34244 18900 35868
rect 18844 34178 18900 34188
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 18732 33684 18788 33694
rect 17836 33124 17892 33134
rect 14700 28466 14756 28476
rect 15036 31332 15092 31342
rect 15036 29988 15092 31276
rect 14364 25442 14420 25452
rect 14252 25218 14308 25228
rect 15036 25172 15092 29932
rect 17836 27076 17892 33068
rect 17836 27010 17892 27020
rect 18732 25844 18788 33628
rect 18732 25778 18788 25788
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 21980 33236 22036 33246
rect 21980 27860 22036 33180
rect 22092 32788 22148 76300
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 34972 69188 35028 69198
rect 31388 67620 31444 67630
rect 31388 59668 31444 67564
rect 33404 63028 33460 63038
rect 31388 59602 31444 59612
rect 31724 62356 31780 62366
rect 23324 56420 23380 56430
rect 22316 55300 22372 55310
rect 22316 49924 22372 55244
rect 22316 49858 22372 49868
rect 22652 52948 22708 52958
rect 22652 47124 22708 52892
rect 23324 51380 23380 56364
rect 28476 56308 28532 56318
rect 25676 55412 25732 55422
rect 23324 51314 23380 51324
rect 25452 55300 25508 55310
rect 25452 50036 25508 55244
rect 25452 49970 25508 49980
rect 25676 47572 25732 55356
rect 28140 54068 28196 54078
rect 28140 50708 28196 54012
rect 28140 50642 28196 50652
rect 25676 47506 25732 47516
rect 26684 49028 26740 49038
rect 22652 47058 22708 47068
rect 26572 46900 26628 46910
rect 22764 46004 22820 46014
rect 22316 44660 22372 44670
rect 22316 36596 22372 44604
rect 22764 43652 22820 45948
rect 22764 43586 22820 43596
rect 24668 45444 24724 45454
rect 22428 41076 22484 41086
rect 22428 39844 22484 41020
rect 22428 39778 22484 39788
rect 24668 38052 24724 45388
rect 24668 37986 24724 37996
rect 26572 37044 26628 46844
rect 26684 46452 26740 48972
rect 26684 46386 26740 46396
rect 26796 47236 26852 47246
rect 26796 46004 26852 47180
rect 26796 45938 26852 45948
rect 26572 36978 26628 36988
rect 22316 36530 22372 36540
rect 22092 32722 22148 32732
rect 27020 28420 27076 28430
rect 21980 27794 22036 27804
rect 23436 27972 23492 27982
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 15036 25106 15092 25116
rect 19808 25116 20128 26628
rect 14028 24322 14084 24332
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 12572 23986 12628 23996
rect 19808 23548 20128 25060
rect 23436 24612 23492 27916
rect 27020 26740 27076 28364
rect 27020 26674 27076 26684
rect 23436 24546 23492 24556
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 16156 23268 16212 23278
rect 4448 21196 4768 22708
rect 15036 22708 15092 22718
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 14700 21924 14756 21934
rect 14700 17556 14756 21868
rect 15036 19348 15092 22652
rect 15036 19282 15092 19292
rect 14700 17490 14756 17500
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 16156 15540 16212 23212
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 16156 15474 16212 15484
rect 19292 15988 19348 15998
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 14476 14644 14532 14654
rect 14476 13524 14532 14588
rect 14476 13458 14532 13468
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 19292 11956 19348 15932
rect 19292 11890 19348 11900
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 20524 22372 20580 22382
rect 20524 13076 20580 22316
rect 20524 13010 20580 13020
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 28476 4564 28532 56252
rect 28812 51156 28868 51166
rect 28700 40628 28756 40638
rect 28700 40068 28756 40572
rect 28700 40002 28756 40012
rect 28812 21028 28868 51100
rect 29260 45668 29316 45678
rect 29036 45556 29092 45566
rect 29036 38388 29092 45500
rect 29036 38322 29092 38332
rect 29260 38276 29316 45612
rect 30940 45332 30996 45342
rect 29260 38210 29316 38220
rect 29708 44884 29764 44894
rect 29708 35364 29764 44828
rect 30940 43876 30996 45276
rect 30044 43652 30100 43662
rect 30044 35476 30100 43596
rect 30044 35410 30100 35420
rect 29708 35298 29764 35308
rect 29596 29876 29652 29886
rect 29596 23716 29652 29820
rect 29708 29652 29764 29662
rect 29708 24612 29764 29596
rect 29708 24546 29764 24556
rect 29596 23650 29652 23660
rect 28812 20962 28868 20972
rect 30940 19572 30996 43820
rect 30940 19506 30996 19516
rect 31052 33684 31108 33694
rect 31052 14868 31108 33628
rect 31724 31892 31780 62300
rect 33404 60564 33460 62972
rect 33404 60498 33460 60508
rect 33404 54964 33460 54974
rect 33404 48804 33460 54908
rect 33404 48738 33460 48748
rect 34748 46676 34804 46686
rect 34636 46452 34692 46462
rect 34636 39284 34692 46396
rect 34636 39218 34692 39228
rect 34748 37380 34804 46620
rect 34748 37314 34804 37324
rect 34972 35364 35028 69132
rect 34972 35298 35028 35308
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 37996 58212 38052 58222
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35756 50932 35812 50942
rect 35756 48692 35812 50876
rect 35756 48626 35812 48636
rect 37660 50596 37716 50606
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 37548 46228 37604 46238
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 36092 41300 36148 41310
rect 36092 38500 36148 41244
rect 36092 38434 36148 38444
rect 35168 36876 35488 38388
rect 37548 37380 37604 46172
rect 37548 37314 37604 37324
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 31724 31826 31780 31836
rect 34748 32564 34804 32574
rect 31724 31332 31780 31342
rect 31724 26852 31780 31276
rect 31724 26786 31780 26796
rect 34748 26628 34804 32508
rect 34748 26562 34804 26572
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 37100 34692 37156 34702
rect 37100 28644 37156 34636
rect 37100 28578 37156 28588
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 31052 14802 31108 14812
rect 35168 25900 35488 27412
rect 37660 27300 37716 50540
rect 37660 27234 37716 27244
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 37996 25060 38052 58156
rect 44604 57652 44660 57662
rect 40796 56868 40852 56878
rect 39228 54292 39284 54302
rect 39228 48804 39284 54236
rect 40796 51716 40852 56812
rect 41020 55972 41076 55982
rect 40796 51650 40852 51660
rect 40908 52948 40964 52958
rect 40908 51156 40964 52892
rect 40908 51090 40964 51100
rect 39228 48738 39284 48748
rect 41020 48132 41076 55916
rect 44604 55972 44660 57596
rect 44604 55906 44660 55916
rect 41692 54740 41748 54750
rect 41244 54180 41300 54190
rect 41244 52836 41300 54124
rect 41244 52770 41300 52780
rect 41132 52388 41188 52398
rect 41132 48580 41188 52332
rect 41692 52388 41748 54684
rect 41692 52322 41748 52332
rect 41132 48514 41188 48524
rect 41580 50820 41636 50830
rect 41020 48066 41076 48076
rect 41244 45556 41300 45566
rect 38668 45444 38724 45454
rect 38668 43316 38724 45388
rect 38668 43250 38724 43260
rect 41244 44324 41300 45500
rect 41244 42868 41300 44268
rect 40236 39620 40292 39630
rect 40236 29316 40292 39564
rect 41244 36484 41300 42812
rect 41244 36418 41300 36428
rect 40236 29250 40292 29260
rect 39004 29204 39060 29214
rect 39004 28084 39060 29148
rect 39004 28018 39060 28028
rect 37996 24994 38052 25004
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 28476 4498 28532 4508
rect 35168 13356 35488 14868
rect 37436 23492 37492 23502
rect 37436 13972 37492 23436
rect 41580 23492 41636 50764
rect 41916 45668 41972 45678
rect 41916 42868 41972 45612
rect 41916 42802 41972 42812
rect 46284 34580 46340 34590
rect 44380 30436 44436 30446
rect 44380 24052 44436 30380
rect 46284 27300 46340 34524
rect 46284 27234 46340 27244
rect 46508 34132 46564 34142
rect 46508 25396 46564 34076
rect 46508 25330 46564 25340
rect 44380 23986 44436 23996
rect 41580 23426 41636 23436
rect 38668 22820 38724 22830
rect 38220 19012 38276 19022
rect 38220 15540 38276 18956
rect 38668 18676 38724 22764
rect 38668 18610 38724 18620
rect 39452 22596 39508 22606
rect 39452 17668 39508 22540
rect 39452 17602 39508 17612
rect 38220 15474 38276 15484
rect 37436 13906 37492 13916
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1463_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14224 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1465_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1466_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1467_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1468_
timestamp 1698431365
transform 1 0 21728 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1469_
timestamp 1698431365
transform -1 0 24864 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1470_
timestamp 1698431365
transform -1 0 24640 0 -1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1471_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22176 0 1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1472_
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1473_
timestamp 1698431365
transform 1 0 18592 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1474_
timestamp 1698431365
transform -1 0 20944 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1475_
timestamp 1698431365
transform 1 0 18144 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1476_
timestamp 1698431365
transform 1 0 19264 0 1 70560
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1477_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6832 0 1 68992
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1478_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1479_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 -1 72128
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1480_
timestamp 1698431365
transform 1 0 21504 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1481_
timestamp 1698431365
transform 1 0 22848 0 -1 70560
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1482_
timestamp 1698431365
transform 1 0 23408 0 1 72128
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1483_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26320 0 1 70560
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1484_
timestamp 1698431365
transform 1 0 17248 0 1 70560
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1485_
timestamp 1698431365
transform 1 0 18256 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1486_
timestamp 1698431365
transform 1 0 19488 0 -1 73696
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1487_
timestamp 1698431365
transform 1 0 17024 0 1 73696
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1488_
timestamp 1698431365
transform -1 0 22064 0 -1 72128
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1489_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6832 0 1 68992
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1490_
timestamp 1698431365
transform 1 0 8176 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1491_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8512 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1492_
timestamp 1698431365
transform -1 0 7392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1493_
timestamp 1698431365
transform -1 0 7056 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1494_
timestamp 1698431365
transform 1 0 5376 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1495_
timestamp 1698431365
transform 1 0 8176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1496_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8064 0 1 70560
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1497_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 70560
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1498_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5712 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11760 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1500_
timestamp 1698431365
transform 1 0 10976 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1501_
timestamp 1698431365
transform 1 0 20048 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1502_
timestamp 1698431365
transform -1 0 21504 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1503_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23520 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1504_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1505_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27216 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1506_
timestamp 1698431365
transform 1 0 39088 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1507_
timestamp 1698431365
transform -1 0 40432 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1508_
timestamp 1698431365
transform -1 0 39424 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1509_
timestamp 1698431365
transform -1 0 36512 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1510_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1511_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21840 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1512_
timestamp 1698431365
transform 1 0 22176 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1513_
timestamp 1698431365
transform 1 0 23296 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1514_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1515_
timestamp 1698431365
transform 1 0 32256 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1516_
timestamp 1698431365
transform -1 0 33152 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1517_
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1518_
timestamp 1698431365
transform -1 0 19040 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1519_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1520_
timestamp 1698431365
transform -1 0 21728 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1521_
timestamp 1698431365
transform -1 0 21616 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1522_
timestamp 1698431365
transform 1 0 22624 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1523_
timestamp 1698431365
transform 1 0 8288 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1524_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 54880
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1525_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25872 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1526_
timestamp 1698431365
transform 1 0 11088 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1698431365
transform 1 0 9744 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1528_
timestamp 1698431365
transform 1 0 10192 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1529_
timestamp 1698431365
transform 1 0 39760 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1530_
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1531_
timestamp 1698431365
transform -1 0 38864 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1532_
timestamp 1698431365
transform -1 0 28448 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1533_
timestamp 1698431365
transform 1 0 31360 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1534_
timestamp 1698431365
transform 1 0 33152 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1535_
timestamp 1698431365
transform -1 0 33152 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1536_
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1537_
timestamp 1698431365
transform 1 0 23408 0 1 56448
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1538_
timestamp 1698431365
transform 1 0 26320 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1539_
timestamp 1698431365
transform 1 0 29792 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1540_
timestamp 1698431365
transform 1 0 31584 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1541_
timestamp 1698431365
transform 1 0 19712 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1542_
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1543_
timestamp 1698431365
transform 1 0 41328 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1544_
timestamp 1698431365
transform 1 0 40880 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1545_
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1546_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23520 0 1 51744
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1698431365
transform 1 0 10528 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1548_
timestamp 1698431365
transform 1 0 12544 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1549_
timestamp 1698431365
transform 1 0 16464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1550_
timestamp 1698431365
transform 1 0 26656 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1551_
timestamp 1698431365
transform -1 0 29568 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1552_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 -1 51744
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1553_
timestamp 1698431365
transform -1 0 31584 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1554_
timestamp 1698431365
transform -1 0 30912 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1555_
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1556_
timestamp 1698431365
transform -1 0 41440 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1557_
timestamp 1698431365
transform 1 0 9632 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1558_
timestamp 1698431365
transform 1 0 23520 0 1 50176
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1559_
timestamp 1698431365
transform -1 0 14896 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1560_
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1561_
timestamp 1698431365
transform 1 0 27328 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1562_
timestamp 1698431365
transform 1 0 25760 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1563_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1564_
timestamp 1698431365
transform -1 0 14672 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1565_
timestamp 1698431365
transform 1 0 14784 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1566_
timestamp 1698431365
transform 1 0 14112 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1567_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15344 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1568_
timestamp 1698431365
transform -1 0 40320 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1569_
timestamp 1698431365
transform -1 0 39984 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1570_
timestamp 1698431365
transform 1 0 26320 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1571_
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1572_
timestamp 1698431365
transform -1 0 31696 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1573_
timestamp 1698431365
transform 1 0 23072 0 1 48608
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1574_
timestamp 1698431365
transform 1 0 26320 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1575_
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1576_
timestamp 1698431365
transform 1 0 17136 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1577_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20608 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1578_
timestamp 1698431365
transform -1 0 18592 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1579_
timestamp 1698431365
transform 1 0 18480 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1580_
timestamp 1698431365
transform 1 0 19488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1582_
timestamp 1698431365
transform -1 0 40544 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1583_
timestamp 1698431365
transform 1 0 30128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1584_
timestamp 1698431365
transform -1 0 31472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1585_
timestamp 1698431365
transform -1 0 30128 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1586_
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1587_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1588_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22960 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1589_
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1590_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1591_
timestamp 1698431365
transform 1 0 18032 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform 1 0 21056 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1593_
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1594_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1595_
timestamp 1698431365
transform 1 0 36960 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1596_
timestamp 1698431365
transform 1 0 37072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1597_
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1598_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1599_
timestamp 1698431365
transform -1 0 4144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1600_
timestamp 1698431365
transform -1 0 20944 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1601_
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_4  _1602_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23296 0 1 36064
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1603_
timestamp 1698431365
transform -1 0 47936 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1604_
timestamp 1698431365
transform 1 0 19488 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1605_
timestamp 1698431365
transform 1 0 21056 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1606_
timestamp 1698431365
transform 1 0 22512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1607_
timestamp 1698431365
transform -1 0 28112 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1608_
timestamp 1698431365
transform 1 0 25648 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_4  _1609_
timestamp 1698431365
transform 1 0 21840 0 1 34496
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1610_
timestamp 1698431365
transform -1 0 47936 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1611_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1612_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1613_
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1614_
timestamp 1698431365
transform -1 0 6384 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1615_
timestamp 1698431365
transform -1 0 20832 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _1616_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1617_
timestamp 1698431365
transform -1 0 47936 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1618_
timestamp 1698431365
transform -1 0 17920 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1619_
timestamp 1698431365
transform -1 0 22736 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1620_
timestamp 1698431365
transform -1 0 20384 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1621_
timestamp 1698431365
transform -1 0 18928 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1622_
timestamp 1698431365
transform -1 0 18816 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1623_
timestamp 1698431365
transform 1 0 18592 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1624_
timestamp 1698431365
transform 1 0 18368 0 -1 54880
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1625_
timestamp 1698431365
transform -1 0 17696 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1626_
timestamp 1698431365
transform -1 0 18816 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1698431365
transform -1 0 17808 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1628_
timestamp 1698431365
transform -1 0 19152 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1629_
timestamp 1698431365
transform 1 0 16464 0 1 54880
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1630_
timestamp 1698431365
transform -1 0 17360 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1698431365
transform -1 0 17024 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1632_
timestamp 1698431365
transform -1 0 18480 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1633_
timestamp 1698431365
transform 1 0 17808 0 -1 59584
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1634_
timestamp 1698431365
transform -1 0 19152 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform -1 0 17808 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1636_
timestamp 1698431365
transform 1 0 18816 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1637_
timestamp 1698431365
transform -1 0 19376 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1638_
timestamp 1698431365
transform 1 0 16464 0 1 56448
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1639_
timestamp 1698431365
transform -1 0 24864 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1640_
timestamp 1698431365
transform 1 0 17696 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1641_
timestamp 1698431365
transform 1 0 21616 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1642_
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1643_
timestamp 1698431365
transform -1 0 23520 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1698431365
transform 1 0 20496 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1645_
timestamp 1698431365
transform 1 0 22288 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1646_
timestamp 1698431365
transform 1 0 21280 0 1 53312
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1647_
timestamp 1698431365
transform 1 0 20384 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1648_
timestamp 1698431365
transform 1 0 20384 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1649_
timestamp 1698431365
transform 1 0 19712 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1650_
timestamp 1698431365
transform 1 0 20384 0 -1 58016
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1651_
timestamp 1698431365
transform 1 0 11424 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1652_
timestamp 1698431365
transform 1 0 11760 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1653_
timestamp 1698431365
transform 1 0 17248 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_4  _1654_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9072 0 -1 68992
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1655_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1656_
timestamp 1698431365
transform 1 0 7168 0 1 67424
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1657_
timestamp 1698431365
transform 1 0 7504 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1658_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1659_
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1660_
timestamp 1698431365
transform -1 0 4032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1661_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 -1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1662_
timestamp 1698431365
transform -1 0 8624 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1663_
timestamp 1698431365
transform -1 0 4368 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1664_
timestamp 1698431365
transform 1 0 7280 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1665_
timestamp 1698431365
transform -1 0 11536 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1666_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1667_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8400 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1668_
timestamp 1698431365
transform -1 0 7280 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_4  _1669_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 -1 54880
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1670_
timestamp 1698431365
transform -1 0 9184 0 -1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1671_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 1 51744
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__and3_4  _1672_
timestamp 1698431365
transform -1 0 5264 0 1 50176
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1673_
timestamp 1698431365
transform -1 0 7056 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1674_
timestamp 1698431365
transform -1 0 9184 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1675_
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1676_
timestamp 1698431365
transform -1 0 8288 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1677_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1678_
timestamp 1698431365
transform -1 0 9184 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1679_
timestamp 1698431365
transform 1 0 6384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1680_
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1681_
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1682_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7280 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1683_
timestamp 1698431365
transform -1 0 6384 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1684_
timestamp 1698431365
transform -1 0 7392 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1685_
timestamp 1698431365
transform -1 0 7056 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1686_
timestamp 1698431365
transform -1 0 8512 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1687_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7728 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1688_
timestamp 1698431365
transform 1 0 15344 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1690_
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1691_
timestamp 1698431365
transform 1 0 30464 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1692_
timestamp 1698431365
transform 1 0 11760 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1693_
timestamp 1698431365
transform 1 0 16240 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1694_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1695_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1696_
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1697_
timestamp 1698431365
transform 1 0 20160 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1698_
timestamp 1698431365
transform 1 0 29904 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1699_
timestamp 1698431365
transform -1 0 31472 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1701_
timestamp 1698431365
transform 1 0 7952 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1702_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1703_
timestamp 1698431365
transform 1 0 7280 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1704_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 1 47040
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1705_
timestamp 1698431365
transform -1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1706_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5936 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1707_
timestamp 1698431365
transform 1 0 6272 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1708_
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1709_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1710_
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1711_
timestamp 1698431365
transform 1 0 14224 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1712_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1713_
timestamp 1698431365
transform -1 0 18816 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1714_
timestamp 1698431365
transform -1 0 20048 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1715_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1716_
timestamp 1698431365
transform 1 0 29456 0 1 58016
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1717_
timestamp 1698431365
transform 1 0 32704 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1718_
timestamp 1698431365
transform 1 0 30912 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1719_
timestamp 1698431365
transform 1 0 38976 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1720_
timestamp 1698431365
transform -1 0 42000 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1721_
timestamp 1698431365
transform 1 0 32928 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1722_
timestamp 1698431365
transform -1 0 39424 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1723_
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1724_
timestamp 1698431365
transform 1 0 38304 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1725_
timestamp 1698431365
transform 1 0 39424 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1726_
timestamp 1698431365
transform -1 0 40320 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1727_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40544 0 -1 61152
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1728_
timestamp 1698431365
transform -1 0 39424 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1729_
timestamp 1698431365
transform 1 0 37632 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1730_
timestamp 1698431365
transform -1 0 38304 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1731_
timestamp 1698431365
transform -1 0 38864 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1732_
timestamp 1698431365
transform 1 0 36960 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1733_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37632 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1734_
timestamp 1698431365
transform 1 0 36960 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1735_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39200 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1736_
timestamp 1698431365
transform -1 0 36624 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1737_
timestamp 1698431365
transform 1 0 37296 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1738_
timestamp 1698431365
transform 1 0 37744 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1739_
timestamp 1698431365
transform -1 0 39088 0 1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1698431365
transform -1 0 37856 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1741_
timestamp 1698431365
transform 1 0 38640 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1742_
timestamp 1698431365
transform -1 0 30576 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1743_
timestamp 1698431365
transform 1 0 19152 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1744_
timestamp 1698431365
transform 1 0 17360 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1745_
timestamp 1698431365
transform 1 0 17584 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1746_
timestamp 1698431365
transform 1 0 18368 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1747_
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1748_
timestamp 1698431365
transform 1 0 7392 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1749_
timestamp 1698431365
transform -1 0 6272 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1750_
timestamp 1698431365
transform 1 0 5936 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1751_
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1752_
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1753_
timestamp 1698431365
transform -1 0 12656 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1754_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1755_
timestamp 1698431365
transform -1 0 15344 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1756_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1757_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1758_
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1759_
timestamp 1698431365
transform 1 0 39536 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1760_
timestamp 1698431365
transform 1 0 39984 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1761_
timestamp 1698431365
transform 1 0 39424 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1762_
timestamp 1698431365
transform 1 0 40320 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1763_
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1764_
timestamp 1698431365
transform 1 0 32480 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform -1 0 41328 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1766_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10864 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1767_
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1768_
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1769_
timestamp 1698431365
transform 1 0 18704 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1770_
timestamp 1698431365
transform -1 0 38864 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1771_
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1773_
timestamp 1698431365
transform 1 0 39760 0 1 56448
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1774_
timestamp 1698431365
transform -1 0 42784 0 1 61152
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1775_
timestamp 1698431365
transform -1 0 41776 0 1 64288
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1776_
timestamp 1698431365
transform -1 0 39872 0 -1 65856
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1777_
timestamp 1698431365
transform 1 0 34720 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1778_
timestamp 1698431365
transform 1 0 35504 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1779_
timestamp 1698431365
transform 1 0 36064 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1780_
timestamp 1698431365
transform 1 0 30912 0 1 58016
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1781_
timestamp 1698431365
transform 1 0 30800 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1782_
timestamp 1698431365
transform 1 0 34608 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1783_
timestamp 1698431365
transform 1 0 36624 0 -1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1784_
timestamp 1698431365
transform 1 0 36512 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1785_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39088 0 -1 65856
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1786_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37856 0 1 65856
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1787_
timestamp 1698431365
transform -1 0 39648 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1698431365
transform -1 0 26880 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1789_
timestamp 1698431365
transform 1 0 14336 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1790_
timestamp 1698431365
transform 1 0 14560 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1791_
timestamp 1698431365
transform 1 0 14896 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1792_
timestamp 1698431365
transform 1 0 13664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1793_
timestamp 1698431365
transform 1 0 13440 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1794_
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1795_
timestamp 1698431365
transform 1 0 11760 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1796_
timestamp 1698431365
transform 1 0 10528 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1797_
timestamp 1698431365
transform -1 0 6720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1798_
timestamp 1698431365
transform 1 0 7728 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1799_
timestamp 1698431365
transform -1 0 5824 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1800_
timestamp 1698431365
transform 1 0 5600 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1801_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6160 0 1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1802_
timestamp 1698431365
transform -1 0 12432 0 1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1803_
timestamp 1698431365
transform -1 0 9184 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1804_
timestamp 1698431365
transform -1 0 8624 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1805_
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1806_
timestamp 1698431365
transform 1 0 8288 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1807_
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1809_
timestamp 1698431365
transform 1 0 11536 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1810_
timestamp 1698431365
transform 1 0 15344 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1811_
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1812_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1813_
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _1814_
timestamp 1698431365
transform 1 0 21504 0 -1 34496
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1815_
timestamp 1698431365
transform -1 0 42336 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1816_
timestamp 1698431365
transform -1 0 43344 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1817_
timestamp 1698431365
transform 1 0 41440 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1818_
timestamp 1698431365
transform 1 0 41776 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1819_
timestamp 1698431365
transform 1 0 41216 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1820_
timestamp 1698431365
transform 1 0 42112 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1821_
timestamp 1698431365
transform 1 0 39536 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1822_
timestamp 1698431365
transform 1 0 39760 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1823_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41776 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1824_
timestamp 1698431365
transform 1 0 40432 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1825_
timestamp 1698431365
transform 1 0 39760 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1826_
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1827_
timestamp 1698431365
transform 1 0 12096 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1828_
timestamp 1698431365
transform 1 0 23296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1829_
timestamp 1698431365
transform 1 0 40320 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1830_
timestamp 1698431365
transform 1 0 40320 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1831_
timestamp 1698431365
transform 1 0 41104 0 1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1832_
timestamp 1698431365
transform 1 0 42336 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1833_
timestamp 1698431365
transform 1 0 42448 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1834_
timestamp 1698431365
transform -1 0 43680 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1835_
timestamp 1698431365
transform -1 0 43344 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1836_
timestamp 1698431365
transform -1 0 43120 0 -1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1837_
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1838_
timestamp 1698431365
transform -1 0 40544 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1839_
timestamp 1698431365
transform -1 0 41664 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1840_
timestamp 1698431365
transform -1 0 42336 0 -1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1841_
timestamp 1698431365
transform -1 0 40320 0 -1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1842_
timestamp 1698431365
transform -1 0 39648 0 1 68992
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1843_
timestamp 1698431365
transform 1 0 25648 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1844_
timestamp 1698431365
transform 1 0 38528 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1845_
timestamp 1698431365
transform 1 0 39312 0 1 67424
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1846_
timestamp 1698431365
transform 1 0 42112 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1847_
timestamp 1698431365
transform 1 0 43456 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1848_
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1849_
timestamp 1698431365
transform -1 0 24080 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1850_
timestamp 1698431365
transform 1 0 21728 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1851_
timestamp 1698431365
transform 1 0 16240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1852_
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1853_
timestamp 1698431365
transform 1 0 16016 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1854_
timestamp 1698431365
transform -1 0 18704 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1855_
timestamp 1698431365
transform -1 0 16800 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1856_
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1858_
timestamp 1698431365
transform 1 0 14672 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1859_
timestamp 1698431365
transform 1 0 15456 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 10640 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1861_
timestamp 1698431365
transform 1 0 11200 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1862_
timestamp 1698431365
transform 1 0 11984 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_
timestamp 1698431365
transform 1 0 12208 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1864_
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1865_
timestamp 1698431365
transform -1 0 10304 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1866_
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1867_
timestamp 1698431365
transform 1 0 6608 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1868_
timestamp 1698431365
transform 1 0 7168 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1869_
timestamp 1698431365
transform 1 0 9520 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1870_
timestamp 1698431365
transform 1 0 10528 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1871_
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1872_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1873_
timestamp 1698431365
transform 1 0 17248 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1874_
timestamp 1698431365
transform 1 0 17696 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1875_
timestamp 1698431365
transform 1 0 21504 0 1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1876_
timestamp 1698431365
transform 1 0 43120 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1877_
timestamp 1698431365
transform 1 0 42896 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1698431365
transform 1 0 43456 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1879_
timestamp 1698431365
transform 1 0 43792 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1880_
timestamp 1698431365
transform 1 0 41888 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1881_
timestamp 1698431365
transform 1 0 42112 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1882_
timestamp 1698431365
transform 1 0 42448 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1883_
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1884_
timestamp 1698431365
transform 1 0 41440 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1885_
timestamp 1698431365
transform 1 0 8064 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1886_
timestamp 1698431365
transform -1 0 10416 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1887_
timestamp 1698431365
transform 1 0 14448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1888_
timestamp 1698431365
transform 1 0 40880 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1889_
timestamp 1698431365
transform 1 0 41328 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1890_
timestamp 1698431365
transform 1 0 42224 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1891_
timestamp 1698431365
transform 1 0 43344 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1892_
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1893_
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1894_
timestamp 1698431365
transform 1 0 40208 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1895_
timestamp 1698431365
transform 1 0 42000 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1896_
timestamp 1698431365
transform 1 0 42224 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1897_
timestamp 1698431365
transform 1 0 43008 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1898_
timestamp 1698431365
transform 1 0 43120 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1899_
timestamp 1698431365
transform 1 0 44016 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1900_
timestamp 1698431365
transform -1 0 46032 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1901_
timestamp 1698431365
transform -1 0 43120 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1902_
timestamp 1698431365
transform 1 0 43680 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1903_
timestamp 1698431365
transform -1 0 44464 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1904_
timestamp 1698431365
transform -1 0 44128 0 -1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1905_
timestamp 1698431365
transform -1 0 43008 0 1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1906_
timestamp 1698431365
transform -1 0 27664 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1907_
timestamp 1698431365
transform -1 0 27664 0 1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1908_
timestamp 1698431365
transform -1 0 26880 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1909_
timestamp 1698431365
transform -1 0 28224 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1910_
timestamp 1698431365
transform 1 0 26432 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1911_
timestamp 1698431365
transform -1 0 45136 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1912_
timestamp 1698431365
transform 1 0 44576 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1913_
timestamp 1698431365
transform 1 0 44128 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1914_
timestamp 1698431365
transform 1 0 43120 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1915_
timestamp 1698431365
transform 1 0 42448 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1698431365
transform 1 0 43792 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1917_
timestamp 1698431365
transform 1 0 45360 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1918_
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform 1 0 45920 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1920_
timestamp 1698431365
transform 1 0 43680 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1921_
timestamp 1698431365
transform -1 0 43344 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1922_
timestamp 1698431365
transform 1 0 43344 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1923_
timestamp 1698431365
transform 1 0 37296 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1924_
timestamp 1698431365
transform 1 0 22624 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1925_
timestamp 1698431365
transform 1 0 21280 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1926_
timestamp 1698431365
transform -1 0 39312 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1927_
timestamp 1698431365
transform 1 0 22288 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1928_
timestamp 1698431365
transform 1 0 17136 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1929_
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1930_
timestamp 1698431365
transform -1 0 19488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1931_
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1932_
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1933_
timestamp 1698431365
transform -1 0 17024 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1934_
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1935_
timestamp 1698431365
transform 1 0 17808 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1936_
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1937_
timestamp 1698431365
transform 1 0 15792 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform 1 0 14672 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1939_
timestamp 1698431365
transform 1 0 14560 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698431365
transform 1 0 14448 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1941_
timestamp 1698431365
transform 1 0 13888 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1942_
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1943_
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1944_
timestamp 1698431365
transform 1 0 11312 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1945_
timestamp 1698431365
transform -1 0 12320 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1946_
timestamp 1698431365
transform -1 0 11312 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1947_
timestamp 1698431365
transform -1 0 12992 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1948_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1949_
timestamp 1698431365
transform 1 0 10864 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1950_
timestamp 1698431365
transform 1 0 12096 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1951_
timestamp 1698431365
transform 1 0 11536 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1952_
timestamp 1698431365
transform 1 0 16576 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1953_
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1954_
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1955_
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform 1 0 43904 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1957_
timestamp 1698431365
transform 1 0 44240 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1698431365
transform 1 0 44576 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1959_
timestamp 1698431365
transform 1 0 45584 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1960_
timestamp 1698431365
transform 1 0 42672 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1961_
timestamp 1698431365
transform -1 0 40432 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1962_
timestamp 1698431365
transform 1 0 40768 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1963_
timestamp 1698431365
transform -1 0 42896 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1964_
timestamp 1698431365
transform 1 0 42896 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1965_
timestamp 1698431365
transform -1 0 39648 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1966_
timestamp 1698431365
transform -1 0 40208 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1967_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40208 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1968_
timestamp 1698431365
transform 1 0 40992 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1969_
timestamp 1698431365
transform -1 0 41440 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1970_
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1971_
timestamp 1698431365
transform 1 0 43008 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1972_
timestamp 1698431365
transform 1 0 44688 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1973_
timestamp 1698431365
transform 1 0 38416 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1974_
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1975_
timestamp 1698431365
transform 1 0 41440 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1976_
timestamp 1698431365
transform 1 0 42224 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1977_
timestamp 1698431365
transform 1 0 43232 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1978_
timestamp 1698431365
transform -1 0 45808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1979_
timestamp 1698431365
transform -1 0 46368 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1980_
timestamp 1698431365
transform -1 0 46032 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1981_
timestamp 1698431365
transform 1 0 45696 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1982_
timestamp 1698431365
transform 1 0 44800 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1983_
timestamp 1698431365
transform 1 0 44576 0 -1 54880
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1984_
timestamp 1698431365
transform -1 0 46704 0 -1 64288
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1985_
timestamp 1698431365
transform -1 0 27104 0 -1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1986_
timestamp 1698431365
transform -1 0 26656 0 -1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1987_
timestamp 1698431365
transform -1 0 25984 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1988_
timestamp 1698431365
transform -1 0 27552 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1698431365
transform 1 0 26096 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1990_
timestamp 1698431365
transform 1 0 45248 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1991_
timestamp 1698431365
transform -1 0 47040 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1992_
timestamp 1698431365
transform 1 0 45584 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1993_
timestamp 1698431365
transform 1 0 45472 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1994_
timestamp 1698431365
transform 1 0 45472 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1995_
timestamp 1698431365
transform -1 0 47264 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1996_
timestamp 1698431365
transform -1 0 46816 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1997_
timestamp 1698431365
transform 1 0 45472 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1998_
timestamp 1698431365
transform 1 0 46144 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform 1 0 46816 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2000_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2001_
timestamp 1698431365
transform 1 0 41328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform 1 0 42896 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2003_
timestamp 1698431365
transform 1 0 39760 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2004_
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2005_
timestamp 1698431365
transform 1 0 42224 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2006_
timestamp 1698431365
transform 1 0 40544 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2007_
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2008_
timestamp 1698431365
transform -1 0 34720 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2009_
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2010_
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2011_
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2012_
timestamp 1698431365
transform -1 0 42112 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2013_
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2014_
timestamp 1698431365
transform 1 0 40880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2015_
timestamp 1698431365
transform 1 0 42112 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2016_
timestamp 1698431365
transform 1 0 42448 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2017_
timestamp 1698431365
transform 1 0 43120 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2018_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2019_
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2020_
timestamp 1698431365
transform 1 0 39200 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2021_
timestamp 1698431365
transform 1 0 42560 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2022_
timestamp 1698431365
transform -1 0 44352 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2023_
timestamp 1698431365
transform -1 0 43904 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _2024_
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2025_
timestamp 1698431365
transform -1 0 23856 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2026_
timestamp 1698431365
transform 1 0 21504 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2027_
timestamp 1698431365
transform 1 0 21056 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2028_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2029_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2030_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1698431365
transform -1 0 21728 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2032_
timestamp 1698431365
transform 1 0 18592 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2033_
timestamp 1698431365
transform -1 0 20160 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2034_
timestamp 1698431365
transform 1 0 15344 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2035_
timestamp 1698431365
transform 1 0 15344 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2036_
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2037_
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2038_
timestamp 1698431365
transform -1 0 20496 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2039_
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2040_
timestamp 1698431365
transform 1 0 9856 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2041_
timestamp 1698431365
transform -1 0 10752 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2042_
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2043_
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2044_
timestamp 1698431365
transform 1 0 11760 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2045_
timestamp 1698431365
transform -1 0 11648 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2046_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform -1 0 18144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2048_
timestamp 1698431365
transform 1 0 15344 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1698431365
transform 1 0 14560 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2050_
timestamp 1698431365
transform 1 0 14000 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2051_
timestamp 1698431365
transform 1 0 15008 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2052_
timestamp 1698431365
transform 1 0 10976 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2053_
timestamp 1698431365
transform -1 0 11984 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2054_
timestamp 1698431365
transform -1 0 12096 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2055_
timestamp 1698431365
transform 1 0 11984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2056_
timestamp 1698431365
transform 1 0 11536 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2057_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2058_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2059_
timestamp 1698431365
transform 1 0 18032 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2060_
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2061_
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2062_
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2063_
timestamp 1698431365
transform -1 0 38192 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2064_
timestamp 1698431365
transform -1 0 38752 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2065_
timestamp 1698431365
transform -1 0 38528 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2066_
timestamp 1698431365
transform -1 0 38192 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2067_
timestamp 1698431365
transform 1 0 35056 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2068_
timestamp 1698431365
transform 1 0 45472 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2069_
timestamp 1698431365
transform 1 0 45136 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2070_
timestamp 1698431365
transform 1 0 45472 0 -1 50176
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2071_
timestamp 1698431365
transform -1 0 47040 0 -1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2072_
timestamp 1698431365
transform -1 0 26880 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2073_
timestamp 1698431365
transform -1 0 26544 0 1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2074_
timestamp 1698431365
transform -1 0 10864 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2075_
timestamp 1698431365
transform -1 0 27776 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2076_
timestamp 1698431365
transform -1 0 26096 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2077_
timestamp 1698431365
transform -1 0 46816 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2078_
timestamp 1698431365
transform 1 0 46256 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2079_
timestamp 1698431365
transform 1 0 45360 0 1 50176
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2080_
timestamp 1698431365
transform 1 0 45248 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2081_
timestamp 1698431365
transform 1 0 45696 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2082_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45808 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2083_
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2084_
timestamp 1698431365
transform 1 0 42448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2085_
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2086_
timestamp 1698431365
transform 1 0 43792 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2087_
timestamp 1698431365
transform -1 0 45584 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2088_
timestamp 1698431365
transform 1 0 42896 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2089_
timestamp 1698431365
transform 1 0 44576 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2091_
timestamp 1698431365
transform -1 0 43120 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2092_
timestamp 1698431365
transform -1 0 42896 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2093_
timestamp 1698431365
transform 1 0 41888 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2094_
timestamp 1698431365
transform 1 0 39536 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2095_
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2096_
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2097_
timestamp 1698431365
transform -1 0 35280 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2098_
timestamp 1698431365
transform 1 0 39312 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2099_
timestamp 1698431365
transform -1 0 39088 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2100_
timestamp 1698431365
transform 1 0 39312 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2101_
timestamp 1698431365
transform 1 0 39984 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2102_
timestamp 1698431365
transform 1 0 42560 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2103_
timestamp 1698431365
transform 1 0 43008 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2104_
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2105_
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2106_
timestamp 1698431365
transform 1 0 37296 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2107_
timestamp 1698431365
transform -1 0 42784 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2108_
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2110_
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2111_
timestamp 1698431365
transform -1 0 26768 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2112_
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2113_
timestamp 1698431365
transform -1 0 20496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2114_
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2115_
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2116_
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2117_
timestamp 1698431365
transform 1 0 21728 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2118_
timestamp 1698431365
transform 1 0 22400 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2119_
timestamp 1698431365
transform 1 0 18368 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2120_
timestamp 1698431365
transform -1 0 20720 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2121_
timestamp 1698431365
transform -1 0 18032 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2122_
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2123_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2124_
timestamp 1698431365
transform -1 0 14672 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2125_
timestamp 1698431365
transform -1 0 13888 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2126_
timestamp 1698431365
transform -1 0 15120 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2127_
timestamp 1698431365
transform 1 0 11312 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2128_
timestamp 1698431365
transform 1 0 13216 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2129_
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2130_
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2131_
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2132_
timestamp 1698431365
transform 1 0 16016 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2133_
timestamp 1698431365
transform 1 0 16576 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2134_
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2135_
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2136_
timestamp 1698431365
transform -1 0 20496 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2137_
timestamp 1698431365
transform 1 0 18816 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2138_
timestamp 1698431365
transform 1 0 20272 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2139_
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2140_
timestamp 1698431365
transform 1 0 23744 0 1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2141_
timestamp 1698431365
transform 1 0 37296 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2142_
timestamp 1698431365
transform 1 0 36400 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2143_
timestamp 1698431365
transform 1 0 37968 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2144_
timestamp 1698431365
transform 1 0 39312 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2145_
timestamp 1698431365
transform 1 0 37968 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2146_
timestamp 1698431365
transform 1 0 41776 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2147_
timestamp 1698431365
transform 1 0 44576 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2148_
timestamp 1698431365
transform 1 0 46032 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2149_
timestamp 1698431365
transform -1 0 47936 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2150_
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2151_
timestamp 1698431365
transform -1 0 27440 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2152_
timestamp 1698431365
transform -1 0 10080 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2153_
timestamp 1698431365
transform 1 0 27440 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2154_
timestamp 1698431365
transform -1 0 28448 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2155_
timestamp 1698431365
transform 1 0 26880 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2156_
timestamp 1698431365
transform -1 0 47040 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2157_
timestamp 1698431365
transform -1 0 48160 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2158_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2159_
timestamp 1698431365
transform 1 0 45472 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2160_
timestamp 1698431365
transform -1 0 46816 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2161_
timestamp 1698431365
transform -1 0 46592 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2162_
timestamp 1698431365
transform 1 0 37856 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2163_
timestamp 1698431365
transform 1 0 40656 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2164_
timestamp 1698431365
transform 1 0 41776 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2165_
timestamp 1698431365
transform 1 0 41552 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2166_
timestamp 1698431365
transform 1 0 42896 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2167_
timestamp 1698431365
transform -1 0 43456 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2168_
timestamp 1698431365
transform 1 0 43680 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2169_
timestamp 1698431365
transform -1 0 45472 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41888 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2171_
timestamp 1698431365
transform -1 0 40768 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2172_
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2173_
timestamp 1698431365
transform 1 0 38976 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2174_
timestamp 1698431365
transform 1 0 38864 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2175_
timestamp 1698431365
transform 1 0 40544 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2176_
timestamp 1698431365
transform 1 0 41440 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2177_
timestamp 1698431365
transform 1 0 42448 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2178_
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2179_
timestamp 1698431365
transform 1 0 39536 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2180_
timestamp 1698431365
transform 1 0 39648 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2181_
timestamp 1698431365
transform -1 0 41328 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2182_
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2183_
timestamp 1698431365
transform 1 0 40096 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2184_
timestamp 1698431365
transform 1 0 23744 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2185_
timestamp 1698431365
transform -1 0 23744 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2186_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2187_
timestamp 1698431365
transform 1 0 21504 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2188_
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2189_
timestamp 1698431365
transform 1 0 21056 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2190_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2191_
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2192_
timestamp 1698431365
transform -1 0 20384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2193_
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2194_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2195_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2196_
timestamp 1698431365
transform 1 0 14112 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2197_
timestamp 1698431365
transform -1 0 16800 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2198_
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2199_
timestamp 1698431365
transform 1 0 14448 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2200_
timestamp 1698431365
transform 1 0 16128 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2201_
timestamp 1698431365
transform 1 0 11088 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2202_
timestamp 1698431365
transform 1 0 12208 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2203_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2204_
timestamp 1698431365
transform -1 0 19040 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2205_
timestamp 1698431365
transform 1 0 17808 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2206_
timestamp 1698431365
transform -1 0 20720 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2207_
timestamp 1698431365
transform 1 0 19264 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2208_
timestamp 1698431365
transform -1 0 19264 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2209_
timestamp 1698431365
transform 1 0 19264 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2210_
timestamp 1698431365
transform 1 0 18256 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2211_
timestamp 1698431365
transform 1 0 19824 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2212_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2213_
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2214_
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2215_
timestamp 1698431365
transform -1 0 36848 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2216_
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2217_
timestamp 1698431365
transform 1 0 36960 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2218_
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2219_
timestamp 1698431365
transform 1 0 40880 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2220_
timestamp 1698431365
transform 1 0 43232 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2221_
timestamp 1698431365
transform 1 0 44576 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2222_
timestamp 1698431365
transform -1 0 46704 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2223_
timestamp 1698431365
transform 1 0 26656 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2224_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2225_
timestamp 1698431365
transform -1 0 29456 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2226_
timestamp 1698431365
transform -1 0 28336 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2227_
timestamp 1698431365
transform -1 0 28896 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2228_
timestamp 1698431365
transform -1 0 27440 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2229_
timestamp 1698431365
transform 1 0 46704 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2230_
timestamp 1698431365
transform 1 0 45584 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2231_
timestamp 1698431365
transform 1 0 45136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2232_
timestamp 1698431365
transform -1 0 44240 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2233_
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2234_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2235_
timestamp 1698431365
transform -1 0 45360 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2236_
timestamp 1698431365
transform 1 0 45360 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2237_
timestamp 1698431365
transform 1 0 40880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2238_
timestamp 1698431365
transform 1 0 41328 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2239_
timestamp 1698431365
transform 1 0 42224 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2240_
timestamp 1698431365
transform 1 0 41776 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform 1 0 42896 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2242_
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2243_
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2244_
timestamp 1698431365
transform 1 0 38304 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2245_
timestamp 1698431365
transform -1 0 38416 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2246_
timestamp 1698431365
transform -1 0 38976 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2247_
timestamp 1698431365
transform 1 0 38864 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2248_
timestamp 1698431365
transform 1 0 23408 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2249_
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2250_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2251_
timestamp 1698431365
transform 1 0 20272 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2252_
timestamp 1698431365
transform -1 0 22064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2253_
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2254_
timestamp 1698431365
transform 1 0 17584 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2255_
timestamp 1698431365
transform -1 0 18816 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2256_
timestamp 1698431365
transform 1 0 14560 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2257_
timestamp 1698431365
transform -1 0 16800 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2258_
timestamp 1698431365
transform -1 0 15456 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2259_
timestamp 1698431365
transform 1 0 13888 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2260_
timestamp 1698431365
transform 1 0 15120 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2261_
timestamp 1698431365
transform 1 0 14672 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2262_
timestamp 1698431365
transform -1 0 16240 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2263_
timestamp 1698431365
transform -1 0 21728 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2264_
timestamp 1698431365
transform -1 0 21952 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1698431365
transform -1 0 20832 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2266_
timestamp 1698431365
transform -1 0 20496 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2267_
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2268_
timestamp 1698431365
transform -1 0 18928 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2269_
timestamp 1698431365
transform 1 0 18592 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2270_
timestamp 1698431365
transform 1 0 18592 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2271_
timestamp 1698431365
transform 1 0 19488 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2272_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform -1 0 28336 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2274_
timestamp 1698431365
transform -1 0 33824 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2275_
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2276_
timestamp 1698431365
transform 1 0 26768 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2277_
timestamp 1698431365
transform 1 0 26656 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2278_
timestamp 1698431365
transform 1 0 25648 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2279_
timestamp 1698431365
transform 1 0 38528 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2280_
timestamp 1698431365
transform 1 0 41552 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2281_
timestamp 1698431365
transform -1 0 37968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2282_
timestamp 1698431365
transform 1 0 38528 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2283_
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2284_
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2285_
timestamp 1698431365
transform -1 0 43344 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2286_
timestamp 1698431365
transform 1 0 41888 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2287_
timestamp 1698431365
transform 1 0 41776 0 1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2288_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2289_
timestamp 1698431365
transform -1 0 46032 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2290_
timestamp 1698431365
transform -1 0 27776 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2291_
timestamp 1698431365
transform -1 0 28000 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2292_
timestamp 1698431365
transform -1 0 6160 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2293_
timestamp 1698431365
transform -1 0 45696 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2294_
timestamp 1698431365
transform 1 0 44240 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2295_
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2296_
timestamp 1698431365
transform -1 0 43904 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2297_
timestamp 1698431365
transform -1 0 44352 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2298_
timestamp 1698431365
transform 1 0 42560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2299_
timestamp 1698431365
transform 1 0 21952 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2300_
timestamp 1698431365
transform -1 0 23968 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2301_
timestamp 1698431365
transform -1 0 21168 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2302_
timestamp 1698431365
transform -1 0 20608 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2303_
timestamp 1698431365
transform -1 0 23968 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2304_
timestamp 1698431365
transform 1 0 21840 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2305_
timestamp 1698431365
transform -1 0 16352 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2306_
timestamp 1698431365
transform -1 0 24640 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2307_
timestamp 1698431365
transform 1 0 21728 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2308_
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2309_
timestamp 1698431365
transform 1 0 22624 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2310_
timestamp 1698431365
transform -1 0 23856 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2311_
timestamp 1698431365
transform -1 0 17360 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2313_
timestamp 1698431365
transform 1 0 15568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2314_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14896 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2315_
timestamp 1698431365
transform 1 0 15568 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2316_
timestamp 1698431365
transform 1 0 22624 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2317_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2318_
timestamp 1698431365
transform 1 0 28000 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2319_
timestamp 1698431365
transform -1 0 28000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2320_
timestamp 1698431365
transform -1 0 28224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2321_
timestamp 1698431365
transform -1 0 41888 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2322_
timestamp 1698431365
transform -1 0 42336 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2323_
timestamp 1698431365
transform 1 0 37856 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2324_
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2325_
timestamp 1698431365
transform 1 0 37968 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2326_
timestamp 1698431365
transform -1 0 39872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2327_
timestamp 1698431365
transform -1 0 39312 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2328_
timestamp 1698431365
transform -1 0 39872 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2329_
timestamp 1698431365
transform 1 0 38528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2330_
timestamp 1698431365
transform 1 0 37184 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2331_
timestamp 1698431365
transform 1 0 40880 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2332_
timestamp 1698431365
transform 1 0 38864 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2333_
timestamp 1698431365
transform -1 0 42000 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2334_
timestamp 1698431365
transform -1 0 42000 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2335_
timestamp 1698431365
transform -1 0 28336 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2336_
timestamp 1698431365
transform -1 0 26320 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2337_
timestamp 1698431365
transform -1 0 28224 0 -1 20384
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2338_
timestamp 1698431365
transform 1 0 3696 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2339_
timestamp 1698431365
transform -1 0 26208 0 1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2340_
timestamp 1698431365
transform -1 0 16464 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2341_
timestamp 1698431365
transform -1 0 7056 0 -1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2342_
timestamp 1698431365
transform 1 0 5600 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2343_
timestamp 1698431365
transform -1 0 7728 0 1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2344_
timestamp 1698431365
transform -1 0 6272 0 -1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2345_
timestamp 1698431365
transform -1 0 4592 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2346_
timestamp 1698431365
transform -1 0 7056 0 1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2347_
timestamp 1698431365
transform -1 0 8064 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2348_
timestamp 1698431365
transform -1 0 6272 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2349_
timestamp 1698431365
transform -1 0 6384 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2350_
timestamp 1698431365
transform -1 0 3696 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2351_
timestamp 1698431365
transform 1 0 8400 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2352_
timestamp 1698431365
transform 1 0 6384 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2353_
timestamp 1698431365
transform -1 0 6944 0 1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2354_
timestamp 1698431365
transform -1 0 6720 0 -1 51744
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2355_
timestamp 1698431365
transform -1 0 2912 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2356_
timestamp 1698431365
transform -1 0 4592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2357_
timestamp 1698431365
transform 1 0 6384 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2358_
timestamp 1698431365
transform 1 0 4704 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2359_
timestamp 1698431365
transform 1 0 4816 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2360_
timestamp 1698431365
transform 1 0 3024 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2361_
timestamp 1698431365
transform 1 0 5600 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2362_
timestamp 1698431365
transform 1 0 5152 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2363_
timestamp 1698431365
transform 1 0 4704 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2364_
timestamp 1698431365
transform 1 0 4032 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2365_
timestamp 1698431365
transform -1 0 5152 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2366_
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2367_
timestamp 1698431365
transform -1 0 6160 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2368_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2369_
timestamp 1698431365
transform -1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2370_
timestamp 1698431365
transform 1 0 4592 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2371_
timestamp 1698431365
transform -1 0 7392 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2372_
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2373_
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2374_
timestamp 1698431365
transform 1 0 3920 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2375_
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2376_
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2377_
timestamp 1698431365
transform -1 0 7392 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2378_
timestamp 1698431365
transform -1 0 3136 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2379_
timestamp 1698431365
transform -1 0 6832 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2380_
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2381_
timestamp 1698431365
transform 1 0 5488 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2382_
timestamp 1698431365
transform -1 0 5264 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2383_
timestamp 1698431365
transform 1 0 3920 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2384_
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2385_
timestamp 1698431365
transform -1 0 6944 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2386_
timestamp 1698431365
transform 1 0 5040 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2387_
timestamp 1698431365
transform -1 0 5040 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2388_
timestamp 1698431365
transform -1 0 6496 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2389_
timestamp 1698431365
transform -1 0 6272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2390_
timestamp 1698431365
transform -1 0 7952 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2391_
timestamp 1698431365
transform -1 0 6944 0 1 64288
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2392_
timestamp 1698431365
transform -1 0 6160 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2393_
timestamp 1698431365
transform -1 0 35280 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2394_
timestamp 1698431365
transform -1 0 34272 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2395_
timestamp 1698431365
transform 1 0 33488 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2396_
timestamp 1698431365
transform 1 0 33600 0 1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2397_
timestamp 1698431365
transform -1 0 35056 0 1 64288
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2398_
timestamp 1698431365
transform -1 0 31920 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2399_
timestamp 1698431365
transform -1 0 34384 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2400_
timestamp 1698431365
transform 1 0 31808 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2401_
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2402_
timestamp 1698431365
transform -1 0 32704 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2403_
timestamp 1698431365
transform 1 0 33600 0 1 65856
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2404_
timestamp 1698431365
transform 1 0 35056 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2405_
timestamp 1698431365
transform 1 0 35392 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2406_
timestamp 1698431365
transform 1 0 35056 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2407_
timestamp 1698431365
transform 1 0 33264 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2408_
timestamp 1698431365
transform -1 0 33712 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2409_
timestamp 1698431365
transform 1 0 32032 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2410_
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2411_
timestamp 1698431365
transform 1 0 34944 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2412_
timestamp 1698431365
transform -1 0 36624 0 1 65856
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2413_
timestamp 1698431365
transform -1 0 35952 0 -1 67424
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2414_
timestamp 1698431365
transform 1 0 31920 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2415_
timestamp 1698431365
transform 1 0 31360 0 1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2416_
timestamp 1698431365
transform -1 0 33936 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2417_
timestamp 1698431365
transform -1 0 33824 0 1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2418_
timestamp 1698431365
transform -1 0 32816 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2419_
timestamp 1698431365
transform -1 0 31808 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2420_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2421_
timestamp 1698431365
transform 1 0 32480 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2422_
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2423_
timestamp 1698431365
transform 1 0 33488 0 -1 68992
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2424_
timestamp 1698431365
transform 1 0 32928 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2425_
timestamp 1698431365
transform -1 0 35392 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2426_
timestamp 1698431365
transform 1 0 35952 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2427_
timestamp 1698431365
transform 1 0 33264 0 1 67424
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2428_
timestamp 1698431365
transform 1 0 36288 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2429_
timestamp 1698431365
transform -1 0 37184 0 -1 65856
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2430_
timestamp 1698431365
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2431_
timestamp 1698431365
transform 1 0 35280 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2432_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2433_
timestamp 1698431365
transform -1 0 37072 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2434_
timestamp 1698431365
transform 1 0 33152 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2435_
timestamp 1698431365
transform 1 0 34048 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2436_
timestamp 1698431365
transform 1 0 33824 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2437_
timestamp 1698431365
transform -1 0 36288 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2438_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2439_
timestamp 1698431365
transform -1 0 33600 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2440_
timestamp 1698431365
transform 1 0 33600 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2441_
timestamp 1698431365
transform 1 0 34944 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2442_
timestamp 1698431365
transform 1 0 35504 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2443_
timestamp 1698431365
transform 1 0 35280 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2444_
timestamp 1698431365
transform -1 0 38640 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2445_
timestamp 1698431365
transform -1 0 34384 0 -1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2446_
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2447_
timestamp 1698431365
transform -1 0 33600 0 1 70560
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2448_
timestamp 1698431365
transform -1 0 34272 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2449_
timestamp 1698431365
transform -1 0 32480 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2450_
timestamp 1698431365
transform -1 0 36624 0 1 70560
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2451_
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2452_
timestamp 1698431365
transform 1 0 38640 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2453_
timestamp 1698431365
transform 1 0 37072 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2454_
timestamp 1698431365
transform 1 0 37072 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2455_
timestamp 1698431365
transform -1 0 36064 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2456_
timestamp 1698431365
transform -1 0 37408 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2457_
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2458_
timestamp 1698431365
transform 1 0 34160 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2459_
timestamp 1698431365
transform 1 0 34944 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2460_
timestamp 1698431365
transform 1 0 35728 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2461_
timestamp 1698431365
transform -1 0 34048 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2462_
timestamp 1698431365
transform -1 0 33264 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2463_
timestamp 1698431365
transform 1 0 33264 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2464_
timestamp 1698431365
transform -1 0 34720 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2465_
timestamp 1698431365
transform 1 0 34720 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2466_
timestamp 1698431365
transform 1 0 36736 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2467_
timestamp 1698431365
transform 1 0 31248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1698431365
transform 1 0 34160 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2469_
timestamp 1698431365
transform 1 0 34944 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2470_
timestamp 1698431365
transform -1 0 36960 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2471_
timestamp 1698431365
transform 1 0 36960 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2472_
timestamp 1698431365
transform -1 0 39424 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2473_
timestamp 1698431365
transform 1 0 37520 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2474_
timestamp 1698431365
transform 1 0 36960 0 1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2475_
timestamp 1698431365
transform -1 0 38864 0 1 70560
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2476_
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2477_
timestamp 1698431365
transform -1 0 31696 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2478_
timestamp 1698431365
transform -1 0 31136 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2479_
timestamp 1698431365
transform -1 0 31248 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2480_
timestamp 1698431365
transform -1 0 31584 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2481_
timestamp 1698431365
transform 1 0 30016 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2482_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38752 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2483_
timestamp 1698431365
transform 1 0 37520 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2484_
timestamp 1698431365
transform 1 0 37968 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2485_
timestamp 1698431365
transform -1 0 40432 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2486_
timestamp 1698431365
transform -1 0 33600 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2487_
timestamp 1698431365
transform -1 0 34272 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2488_
timestamp 1698431365
transform 1 0 35280 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2489_
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2490_
timestamp 1698431365
transform 1 0 37072 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2491_
timestamp 1698431365
transform -1 0 38416 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2492_
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2493_
timestamp 1698431365
transform 1 0 36736 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2494_
timestamp 1698431365
transform -1 0 38192 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2495_
timestamp 1698431365
transform 1 0 37072 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2496_
timestamp 1698431365
transform 1 0 34384 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2497_
timestamp 1698431365
transform 1 0 34608 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2498_
timestamp 1698431365
transform 1 0 31248 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2499_
timestamp 1698431365
transform 1 0 29568 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform 1 0 29680 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2501_
timestamp 1698431365
transform 1 0 30240 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2502_
timestamp 1698431365
transform 1 0 31248 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2503_
timestamp 1698431365
transform 1 0 34048 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2504_
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2505_
timestamp 1698431365
transform 1 0 34272 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2506_
timestamp 1698431365
transform 1 0 34272 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2507_
timestamp 1698431365
transform -1 0 36512 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2508_
timestamp 1698431365
transform 1 0 34608 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2509_
timestamp 1698431365
transform 1 0 35168 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2510_
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2511_
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2512_
timestamp 1698431365
transform 1 0 37408 0 1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2513_
timestamp 1698431365
transform 1 0 37408 0 -1 37632
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2514_
timestamp 1698431365
transform -1 0 35392 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2515_
timestamp 1698431365
transform -1 0 37072 0 -1 72128
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2516_
timestamp 1698431365
transform 1 0 27328 0 -1 67424
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2517_
timestamp 1698431365
transform -1 0 29680 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2518_
timestamp 1698431365
transform -1 0 28224 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2519_
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2520_
timestamp 1698431365
transform 1 0 29232 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2521_
timestamp 1698431365
transform 1 0 30016 0 -1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2522_
timestamp 1698431365
transform 1 0 29120 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2523_
timestamp 1698431365
transform -1 0 39536 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2524_
timestamp 1698431365
transform 1 0 39536 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2525_
timestamp 1698431365
transform -1 0 38976 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2526_
timestamp 1698431365
transform -1 0 40208 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2527_
timestamp 1698431365
transform -1 0 39536 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2528_
timestamp 1698431365
transform 1 0 37744 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2529_
timestamp 1698431365
transform -1 0 38976 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2530_
timestamp 1698431365
transform 1 0 35392 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2531_
timestamp 1698431365
transform -1 0 37072 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2532_
timestamp 1698431365
transform -1 0 36512 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2533_
timestamp 1698431365
transform 1 0 31696 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2534_
timestamp 1698431365
transform -1 0 31248 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2535_
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2536_
timestamp 1698431365
transform -1 0 31024 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2537_
timestamp 1698431365
transform -1 0 30912 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2538_
timestamp 1698431365
transform 1 0 27552 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2539_
timestamp 1698431365
transform 1 0 29008 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2540_
timestamp 1698431365
transform 1 0 30688 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2541_
timestamp 1698431365
transform 1 0 32144 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2542_
timestamp 1698431365
transform -1 0 33488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1698431365
transform 1 0 32256 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2544_
timestamp 1698431365
transform -1 0 34384 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2545_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2546_
timestamp 1698431365
transform 1 0 35056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2547_
timestamp 1698431365
transform 1 0 34832 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2548_
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2549_
timestamp 1698431365
transform -1 0 40544 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2550_
timestamp 1698431365
transform 1 0 35056 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2551_
timestamp 1698431365
transform -1 0 36848 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2552_
timestamp 1698431365
transform -1 0 36400 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2553_
timestamp 1698431365
transform -1 0 36512 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2554_
timestamp 1698431365
transform 1 0 33376 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2555_
timestamp 1698431365
transform -1 0 36736 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2556_
timestamp 1698431365
transform 1 0 35616 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2557_
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2558_
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2559_
timestamp 1698431365
transform -1 0 30352 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2560_
timestamp 1698431365
transform 1 0 28112 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2561_
timestamp 1698431365
transform -1 0 30464 0 1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2562_
timestamp 1698431365
transform 1 0 29120 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2563_
timestamp 1698431365
transform -1 0 31024 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2564_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2565_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34048 0 -1 36064
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2566_
timestamp 1698431365
transform -1 0 38192 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2567_
timestamp 1698431365
transform -1 0 39536 0 -1 31360
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2568_
timestamp 1698431365
transform 1 0 35056 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2569_
timestamp 1698431365
transform 1 0 35728 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2570_
timestamp 1698431365
transform -1 0 36400 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2571_
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2572_
timestamp 1698431365
transform -1 0 36288 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2573_
timestamp 1698431365
transform -1 0 31360 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2574_
timestamp 1698431365
transform -1 0 31696 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2575_
timestamp 1698431365
transform 1 0 31696 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2576_
timestamp 1698431365
transform 1 0 31472 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2577_
timestamp 1698431365
transform -1 0 29008 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2578_
timestamp 1698431365
transform 1 0 30240 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2579_
timestamp 1698431365
transform 1 0 29344 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2580_
timestamp 1698431365
transform 1 0 29232 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2581_
timestamp 1698431365
transform -1 0 30576 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2582_
timestamp 1698431365
transform -1 0 31920 0 -1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2583_
timestamp 1698431365
transform -1 0 34608 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2584_
timestamp 1698431365
transform -1 0 36400 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2585_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2586_
timestamp 1698431365
transform -1 0 34272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2587_
timestamp 1698431365
transform 1 0 30800 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2588_
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2589_
timestamp 1698431365
transform 1 0 32816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2590_
timestamp 1698431365
transform 1 0 33600 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2591_
timestamp 1698431365
transform 1 0 35392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2592_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2593_
timestamp 1698431365
transform 1 0 36064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2594_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2595_
timestamp 1698431365
transform 1 0 32704 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2596_
timestamp 1698431365
transform -1 0 36288 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2597_
timestamp 1698431365
transform -1 0 37408 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2598_
timestamp 1698431365
transform -1 0 35952 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2599_
timestamp 1698431365
transform 1 0 32256 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2600_
timestamp 1698431365
transform -1 0 36064 0 -1 20384
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2601_
timestamp 1698431365
transform -1 0 34384 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2602_
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2603_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _2604_
timestamp 1698431365
transform 1 0 28560 0 -1 62720
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2605_
timestamp 1698431365
transform 1 0 29904 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2606_
timestamp 1698431365
transform 1 0 31584 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2607_
timestamp 1698431365
transform -1 0 25760 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _2608_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31248 0 -1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2609_
timestamp 1698431365
transform 1 0 31584 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2610_
timestamp 1698431365
transform -1 0 29456 0 -1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2611_
timestamp 1698431365
transform 1 0 18704 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2612_
timestamp 1698431365
transform 1 0 31360 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2613_
timestamp 1698431365
transform -1 0 34272 0 1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2614_
timestamp 1698431365
transform -1 0 34272 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2615_
timestamp 1698431365
transform 1 0 33488 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2616_
timestamp 1698431365
transform 1 0 32480 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2617_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2618_
timestamp 1698431365
transform -1 0 34944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2619_
timestamp 1698431365
transform -1 0 34160 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2620_
timestamp 1698431365
transform -1 0 34048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2621_
timestamp 1698431365
transform 1 0 32144 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2622_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2623_
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2624_
timestamp 1698431365
transform 1 0 31136 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2625_
timestamp 1698431365
transform 1 0 29232 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2626_
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2627_
timestamp 1698431365
transform -1 0 32592 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2628_
timestamp 1698431365
transform 1 0 31136 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2629_
timestamp 1698431365
transform 1 0 31248 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2630_
timestamp 1698431365
transform -1 0 32368 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2631_
timestamp 1698431365
transform 1 0 30800 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2632_
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2633_
timestamp 1698431365
transform 1 0 31808 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2634_
timestamp 1698431365
transform -1 0 36176 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2635_
timestamp 1698431365
transform -1 0 35728 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2636_
timestamp 1698431365
transform 1 0 34608 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2637_
timestamp 1698431365
transform -1 0 35840 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2638_
timestamp 1698431365
transform -1 0 35056 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2639_
timestamp 1698431365
transform 1 0 32816 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2640_
timestamp 1698431365
transform -1 0 37408 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2641_
timestamp 1698431365
transform -1 0 36400 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2642_
timestamp 1698431365
transform -1 0 37296 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2643_
timestamp 1698431365
transform 1 0 33376 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2644_
timestamp 1698431365
transform -1 0 36512 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2645_
timestamp 1698431365
transform -1 0 34496 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2646_
timestamp 1698431365
transform -1 0 33376 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2647_
timestamp 1698431365
transform -1 0 30912 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2648_
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2649_
timestamp 1698431365
transform -1 0 28784 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2650_
timestamp 1698431365
transform -1 0 27776 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2651_
timestamp 1698431365
transform -1 0 28784 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2652_
timestamp 1698431365
transform -1 0 29568 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2653_
timestamp 1698431365
transform -1 0 28784 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2654_
timestamp 1698431365
transform -1 0 31360 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2655_
timestamp 1698431365
transform 1 0 31360 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2656_
timestamp 1698431365
transform -1 0 31808 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2657_
timestamp 1698431365
transform -1 0 32144 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2658_
timestamp 1698431365
transform -1 0 32592 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2659_
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2660_
timestamp 1698431365
transform -1 0 36176 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2661_
timestamp 1698431365
transform -1 0 35616 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2662_
timestamp 1698431365
transform -1 0 35728 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2663_
timestamp 1698431365
transform 1 0 34608 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2664_
timestamp 1698431365
transform -1 0 34944 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2665_
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2666_
timestamp 1698431365
transform -1 0 33488 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2667_
timestamp 1698431365
transform -1 0 33488 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2668_
timestamp 1698431365
transform -1 0 36288 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2669_
timestamp 1698431365
transform 1 0 35168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2670_
timestamp 1698431365
transform -1 0 32032 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2671_
timestamp 1698431365
transform -1 0 32144 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2672_
timestamp 1698431365
transform 1 0 25200 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2673_
timestamp 1698431365
transform 1 0 24304 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2674_
timestamp 1698431365
transform 1 0 25312 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2675_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2676_
timestamp 1698431365
transform 1 0 29792 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2677_
timestamp 1698431365
transform -1 0 32032 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2678_
timestamp 1698431365
transform -1 0 32032 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2679_
timestamp 1698431365
transform 1 0 30128 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2680_
timestamp 1698431365
transform -1 0 31136 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2681_
timestamp 1698431365
transform 1 0 30352 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2682_
timestamp 1698431365
transform -1 0 32032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2683_
timestamp 1698431365
transform 1 0 31024 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2684_
timestamp 1698431365
transform 1 0 31360 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2685_
timestamp 1698431365
transform -1 0 34272 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2686_
timestamp 1698431365
transform -1 0 30688 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2687_
timestamp 1698431365
transform -1 0 30352 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2688_
timestamp 1698431365
transform -1 0 26432 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2689_
timestamp 1698431365
transform -1 0 26096 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2690_
timestamp 1698431365
transform -1 0 19936 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2691_
timestamp 1698431365
transform 1 0 25088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2692_
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2693_
timestamp 1698431365
transform -1 0 30912 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2694_
timestamp 1698431365
transform -1 0 30464 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2695_
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2696_
timestamp 1698431365
transform -1 0 30800 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2697_
timestamp 1698431365
transform 1 0 34272 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2698_
timestamp 1698431365
transform 1 0 31136 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2699_
timestamp 1698431365
transform -1 0 33824 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2700_
timestamp 1698431365
transform 1 0 26096 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2701_
timestamp 1698431365
transform 1 0 25536 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2702_
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2703_
timestamp 1698431365
transform 1 0 26656 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2704_
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2705_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2706_
timestamp 1698431365
transform -1 0 32368 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2707_
timestamp 1698431365
transform 1 0 31024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2708_
timestamp 1698431365
transform -1 0 30800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2709_
timestamp 1698431365
transform -1 0 29792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2710_
timestamp 1698431365
transform 1 0 29792 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2711_
timestamp 1698431365
transform 1 0 29456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2712_
timestamp 1698431365
transform 1 0 29568 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2713_
timestamp 1698431365
transform 1 0 29120 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2714_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2715_
timestamp 1698431365
transform 1 0 28224 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2716_
timestamp 1698431365
transform -1 0 31584 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2717_
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2718_
timestamp 1698431365
transform -1 0 30240 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2719_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2720_
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2721_
timestamp 1698431365
transform 1 0 32032 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2722_
timestamp 1698431365
transform -1 0 33600 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2723_
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2724_
timestamp 1698431365
transform -1 0 19936 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2725_
timestamp 1698431365
transform 1 0 19488 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2726_
timestamp 1698431365
transform -1 0 3136 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2727_
timestamp 1698431365
transform 1 0 9408 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2728_
timestamp 1698431365
transform 1 0 10080 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2729_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2730_
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2731_
timestamp 1698431365
transform -1 0 3360 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2732_
timestamp 1698431365
transform 1 0 19936 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2733_
timestamp 1698431365
transform -1 0 20608 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2734_
timestamp 1698431365
transform -1 0 10752 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2735_
timestamp 1698431365
transform -1 0 8624 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2736_
timestamp 1698431365
transform 1 0 19712 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2737_
timestamp 1698431365
transform -1 0 19376 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2738_
timestamp 1698431365
transform 1 0 8624 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2739_
timestamp 1698431365
transform 1 0 14672 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2740_
timestamp 1698431365
transform 1 0 15344 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2741_
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2742_
timestamp 1698431365
transform -1 0 10304 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2743_
timestamp 1698431365
transform -1 0 9744 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2744_
timestamp 1698431365
transform 1 0 9184 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2745_
timestamp 1698431365
transform -1 0 2688 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2746_
timestamp 1698431365
transform -1 0 3808 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2747_
timestamp 1698431365
transform -1 0 2352 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2748_
timestamp 1698431365
transform 1 0 2016 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2749_
timestamp 1698431365
transform -1 0 10864 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2750_
timestamp 1698431365
transform 1 0 8624 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2751_
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2752_
timestamp 1698431365
transform 1 0 2016 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2753_
timestamp 1698431365
transform 1 0 10080 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2754_
timestamp 1698431365
transform -1 0 10080 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2755_
timestamp 1698431365
transform 1 0 2016 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2756_
timestamp 1698431365
transform 1 0 3808 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2757_
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2758_
timestamp 1698431365
transform -1 0 3360 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2759_
timestamp 1698431365
transform 1 0 2016 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2760_
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2761_
timestamp 1698431365
transform -1 0 10528 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2762_
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2763_
timestamp 1698431365
transform -1 0 19712 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2764_
timestamp 1698431365
transform -1 0 10416 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2765_
timestamp 1698431365
transform 1 0 10192 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2766_
timestamp 1698431365
transform 1 0 8624 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2767_
timestamp 1698431365
transform -1 0 18256 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2768_
timestamp 1698431365
transform -1 0 14000 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2769_
timestamp 1698431365
transform -1 0 14896 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2770_
timestamp 1698431365
transform -1 0 12096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2771_
timestamp 1698431365
transform -1 0 11872 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2772_
timestamp 1698431365
transform -1 0 11424 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2773_
timestamp 1698431365
transform -1 0 11648 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2774_
timestamp 1698431365
transform 1 0 16576 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2775_
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2776_
timestamp 1698431365
transform -1 0 18480 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2777_
timestamp 1698431365
transform -1 0 15904 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2778_
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2779_
timestamp 1698431365
transform -1 0 16576 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2780_
timestamp 1698431365
transform -1 0 16912 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2781_
timestamp 1698431365
transform 1 0 14896 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2782_
timestamp 1698431365
transform 1 0 15456 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2783_
timestamp 1698431365
transform -1 0 16352 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2784_
timestamp 1698431365
transform -1 0 13888 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2785_
timestamp 1698431365
transform -1 0 12992 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2786_
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2787_
timestamp 1698431365
transform 1 0 13664 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2788_
timestamp 1698431365
transform 1 0 13552 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2789_
timestamp 1698431365
transform -1 0 17472 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2790_
timestamp 1698431365
transform 1 0 15232 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2791_
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2792_
timestamp 1698431365
transform 1 0 16464 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2793_
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2794_
timestamp 1698431365
transform 1 0 16688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2795_
timestamp 1698431365
transform -1 0 18816 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2796_
timestamp 1698431365
transform -1 0 18256 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2797_
timestamp 1698431365
transform -1 0 14896 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2798_
timestamp 1698431365
transform 1 0 12544 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2799_
timestamp 1698431365
transform -1 0 18256 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2800_
timestamp 1698431365
transform -1 0 12320 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2801_
timestamp 1698431365
transform 1 0 11088 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2802_
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2803_
timestamp 1698431365
transform -1 0 12544 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2804_
timestamp 1698431365
transform -1 0 11536 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2805_
timestamp 1698431365
transform -1 0 16128 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2806_
timestamp 1698431365
transform 1 0 11088 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2807_
timestamp 1698431365
transform -1 0 12544 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2808_
timestamp 1698431365
transform 1 0 11536 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2809_
timestamp 1698431365
transform 1 0 11984 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2810_
timestamp 1698431365
transform -1 0 13104 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2811_
timestamp 1698431365
transform -1 0 11088 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2812_
timestamp 1698431365
transform 1 0 11088 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2813_
timestamp 1698431365
transform 1 0 17584 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2814_
timestamp 1698431365
transform -1 0 18480 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2815_
timestamp 1698431365
transform 1 0 16688 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2816_
timestamp 1698431365
transform -1 0 17808 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2817_
timestamp 1698431365
transform -1 0 17024 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2818_
timestamp 1698431365
transform 1 0 22512 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2819_
timestamp 1698431365
transform 1 0 19600 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2820_
timestamp 1698431365
transform -1 0 25760 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2821_
timestamp 1698431365
transform 1 0 21616 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2822_
timestamp 1698431365
transform 1 0 22512 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2823_
timestamp 1698431365
transform 1 0 19040 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2824_
timestamp 1698431365
transform 1 0 21616 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2825_
timestamp 1698431365
transform -1 0 20720 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2826_
timestamp 1698431365
transform 1 0 18480 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2827_
timestamp 1698431365
transform 1 0 19824 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2828_
timestamp 1698431365
transform 1 0 22064 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2829_
timestamp 1698431365
transform 1 0 23856 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2830_
timestamp 1698431365
transform -1 0 25872 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2831_
timestamp 1698431365
transform 1 0 21280 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2832_
timestamp 1698431365
transform 1 0 22848 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2833_
timestamp 1698431365
transform 1 0 23744 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2834_
timestamp 1698431365
transform 1 0 24640 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2835_
timestamp 1698431365
transform -1 0 27216 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2836_
timestamp 1698431365
transform 1 0 23968 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2837_
timestamp 1698431365
transform 1 0 24528 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2838_
timestamp 1698431365
transform 1 0 25760 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2839_
timestamp 1698431365
transform 1 0 24304 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2840_
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2841_
timestamp 1698431365
transform -1 0 27328 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2842_
timestamp 1698431365
transform 1 0 27328 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2843_
timestamp 1698431365
transform -1 0 23296 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2844_
timestamp 1698431365
transform 1 0 25536 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2845_
timestamp 1698431365
transform 1 0 23744 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2846_
timestamp 1698431365
transform 1 0 25536 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2847_
timestamp 1698431365
transform 1 0 22176 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2848_
timestamp 1698431365
transform -1 0 22176 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2849_
timestamp 1698431365
transform 1 0 25872 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2850_
timestamp 1698431365
transform -1 0 24864 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2851_
timestamp 1698431365
transform 1 0 22848 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2852_
timestamp 1698431365
transform 1 0 14000 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2853_
timestamp 1698431365
transform 1 0 23408 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2854_
timestamp 1698431365
transform 1 0 23968 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2855_
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2856_
timestamp 1698431365
transform 1 0 23408 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2857_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2858_
timestamp 1698431365
transform -1 0 25200 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2859_
timestamp 1698431365
transform 1 0 22288 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2860_
timestamp 1698431365
transform -1 0 24864 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2861_
timestamp 1698431365
transform -1 0 15904 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2862_
timestamp 1698431365
transform -1 0 19152 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2863_
timestamp 1698431365
transform -1 0 16128 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2864_
timestamp 1698431365
transform -1 0 15120 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2865_
timestamp 1698431365
transform -1 0 14336 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2866_
timestamp 1698431365
transform -1 0 14336 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2867_
timestamp 1698431365
transform 1 0 13664 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2868_
timestamp 1698431365
transform -1 0 15232 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2869_
timestamp 1698431365
transform 1 0 13776 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2870_
timestamp 1698431365
transform -1 0 15456 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2871_
timestamp 1698431365
transform 1 0 16128 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2872_
timestamp 1698431365
transform 1 0 14112 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2873_
timestamp 1698431365
transform -1 0 15456 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2874_
timestamp 1698431365
transform 1 0 16800 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2875_
timestamp 1698431365
transform -1 0 18704 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2876_
timestamp 1698431365
transform -1 0 18032 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2877_
timestamp 1698431365
transform -1 0 18592 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2878_
timestamp 1698431365
transform 1 0 19824 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2879_
timestamp 1698431365
transform -1 0 22288 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2880_
timestamp 1698431365
transform 1 0 19936 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2881_
timestamp 1698431365
transform -1 0 21168 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2882_
timestamp 1698431365
transform -1 0 19376 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2883_
timestamp 1698431365
transform -1 0 19936 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2884_
timestamp 1698431365
transform -1 0 22624 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2885_
timestamp 1698431365
transform 1 0 23184 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2886_
timestamp 1698431365
transform 1 0 24864 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2887_
timestamp 1698431365
transform -1 0 20608 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2888_
timestamp 1698431365
transform 1 0 19936 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2889_
timestamp 1698431365
transform 1 0 21952 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2890_
timestamp 1698431365
transform 1 0 22848 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2891_
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2892_
timestamp 1698431365
transform 1 0 25984 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2893_
timestamp 1698431365
transform 1 0 24080 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2894_
timestamp 1698431365
transform 1 0 23744 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2895_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2896_
timestamp 1698431365
transform 1 0 23072 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2897_
timestamp 1698431365
transform -1 0 26208 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2898_
timestamp 1698431365
transform 1 0 21616 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2899_
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2900_
timestamp 1698431365
transform 1 0 23744 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2901_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2902_
timestamp 1698431365
transform 1 0 24304 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2903_
timestamp 1698431365
transform 1 0 23856 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2904_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2905_
timestamp 1698431365
transform 1 0 22624 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2906_
timestamp 1698431365
transform -1 0 25872 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2907_
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2908_
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2909_
timestamp 1698431365
transform 1 0 23968 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2910_
timestamp 1698431365
transform -1 0 23408 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2911_
timestamp 1698431365
transform 1 0 21392 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2912_
timestamp 1698431365
transform -1 0 16912 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2913_
timestamp 1698431365
transform -1 0 22848 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2914_
timestamp 1698431365
transform 1 0 19040 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2915_
timestamp 1698431365
transform 1 0 15344 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2916_
timestamp 1698431365
transform -1 0 16576 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2917_
timestamp 1698431365
transform -1 0 18256 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2918_
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2919_
timestamp 1698431365
transform 1 0 14000 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2920_
timestamp 1698431365
transform 1 0 14560 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2921_
timestamp 1698431365
transform 1 0 16128 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2922_
timestamp 1698431365
transform 1 0 14000 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2923_
timestamp 1698431365
transform 1 0 15232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2924_
timestamp 1698431365
transform -1 0 16240 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2925_
timestamp 1698431365
transform -1 0 13776 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2926_
timestamp 1698431365
transform 1 0 14784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2927_
timestamp 1698431365
transform -1 0 16016 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2928_
timestamp 1698431365
transform 1 0 13664 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2929_
timestamp 1698431365
transform -1 0 14896 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2930_
timestamp 1698431365
transform 1 0 14112 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2931_
timestamp 1698431365
transform -1 0 14000 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2932_
timestamp 1698431365
transform -1 0 13888 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2933_
timestamp 1698431365
transform -1 0 12768 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2934_
timestamp 1698431365
transform 1 0 11312 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2935_
timestamp 1698431365
transform 1 0 11872 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2936_
timestamp 1698431365
transform -1 0 13888 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2937_
timestamp 1698431365
transform 1 0 11312 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2938_
timestamp 1698431365
transform 1 0 11648 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2939_
timestamp 1698431365
transform -1 0 13888 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2940_
timestamp 1698431365
transform 1 0 11760 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2941_
timestamp 1698431365
transform 1 0 12096 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2942_
timestamp 1698431365
transform -1 0 12544 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2943_
timestamp 1698431365
transform -1 0 11312 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2944_
timestamp 1698431365
transform 1 0 10528 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2945_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2946_
timestamp 1698431365
transform 1 0 1792 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2947_
timestamp 1698431365
transform 1 0 31696 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2948_
timestamp 1698431365
transform 1 0 29344 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2949_
timestamp 1698431365
transform 1 0 25760 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2950_
timestamp 1698431365
transform -1 0 32256 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2951_
timestamp 1698431365
transform 1 0 22960 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2952_
timestamp 1698431365
transform -1 0 23744 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2953_
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2954_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2955_
timestamp 1698431365
transform 1 0 13776 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2956_
timestamp 1698431365
transform -1 0 16576 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2957_
timestamp 1698431365
transform 1 0 10416 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2958_
timestamp 1698431365
transform 1 0 8960 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2959_
timestamp 1698431365
transform 1 0 7392 0 1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2960_
timestamp 1698431365
transform 1 0 5712 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2961_
timestamp 1698431365
transform 1 0 3920 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2962_
timestamp 1698431365
transform -1 0 5040 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2963_
timestamp 1698431365
transform -1 0 7392 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2964_
timestamp 1698431365
transform 1 0 4144 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2965_
timestamp 1698431365
transform 1 0 2016 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2966_
timestamp 1698431365
transform 1 0 1792 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2967_
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2968_
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2969_
timestamp 1698431365
transform 1 0 4144 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2970_
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2971_
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2972_
timestamp 1698431365
transform 1 0 5488 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2973_
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2974_
timestamp 1698431365
transform -1 0 10416 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2975_
timestamp 1698431365
transform -1 0 10976 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2976_
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2977_
timestamp 1698431365
transform -1 0 11536 0 1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2978_
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2979_
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2980_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2981_
timestamp 1698431365
transform 1 0 8736 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2982_
timestamp 1698431365
transform -1 0 9632 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2983_
timestamp 1698431365
transform 1 0 9520 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2984_
timestamp 1698431365
transform -1 0 12656 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2985_
timestamp 1698431365
transform -1 0 13216 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2986_
timestamp 1698431365
transform 1 0 11984 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2987_
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2988_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2989_
timestamp 1698431365
transform 1 0 14448 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2990_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2991_
timestamp 1698431365
transform 1 0 11088 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2992_
timestamp 1698431365
transform 1 0 9744 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2993_
timestamp 1698431365
transform 1 0 9744 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2994_
timestamp 1698431365
transform 1 0 9632 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2995_
timestamp 1698431365
transform 1 0 15232 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2996_
timestamp 1698431365
transform 1 0 21504 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2997_
timestamp 1698431365
transform 1 0 21616 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2998_
timestamp 1698431365
transform 1 0 18256 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2999_
timestamp 1698431365
transform 1 0 25536 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3000_
timestamp 1698431365
transform 1 0 26880 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3001_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3002_
timestamp 1698431365
transform 1 0 28336 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3003_
timestamp 1698431365
transform 1 0 27216 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3004_
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3005_
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3006_
timestamp 1698431365
transform 1 0 24976 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3007_
timestamp 1698431365
transform 1 0 12208 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3008_
timestamp 1698431365
transform 1 0 13552 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3009_
timestamp 1698431365
transform 1 0 14000 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3010_
timestamp 1698431365
transform 1 0 13552 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3011_
timestamp 1698431365
transform 1 0 16016 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3012_
timestamp 1698431365
transform 1 0 21504 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3013_
timestamp 1698431365
transform 1 0 21168 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3014_
timestamp 1698431365
transform 1 0 17696 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3015_
timestamp 1698431365
transform 1 0 27664 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3016_
timestamp 1698431365
transform 1 0 26544 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3017_
timestamp 1698431365
transform 1 0 26208 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3018_
timestamp 1698431365
transform 1 0 26320 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3019_
timestamp 1698431365
transform 1 0 26544 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3020_
timestamp 1698431365
transform 1 0 25648 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3021_
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3022_
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3023_
timestamp 1698431365
transform 1 0 13216 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3024_
timestamp 1698431365
transform 1 0 14672 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3025_
timestamp 1698431365
transform 1 0 13776 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3026_
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3027_
timestamp 1698431365
transform 1 0 10752 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3028_
timestamp 1698431365
transform 1 0 9856 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3029_
timestamp 1698431365
transform 1 0 10864 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3030_
timestamp 1698431365
transform 1 0 9632 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5488 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_2
timestamp 1698431365
transform -1 0 3472 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__A1
timestamp 1698431365
transform 1 0 20608 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__A2
timestamp 1698431365
transform 1 0 22400 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__A1
timestamp 1698431365
transform -1 0 21728 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__A2
timestamp 1698431365
transform 1 0 23072 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A1
timestamp 1698431365
transform 1 0 26656 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1698431365
transform 1 0 26208 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__A2
timestamp 1698431365
transform -1 0 24864 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A1
timestamp 1698431365
transform 1 0 16800 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A2
timestamp 1698431365
transform -1 0 18816 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A2
timestamp 1698431365
transform 1 0 20160 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A1
timestamp 1698431365
transform 1 0 17920 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1698431365
transform 1 0 20160 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A1
timestamp 1698431365
transform 1 0 9744 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__I
timestamp 1698431365
transform 1 0 8960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__A2
timestamp 1698431365
transform 1 0 24304 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__A2
timestamp 1698431365
transform 1 0 22736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__A2
timestamp 1698431365
transform 1 0 25312 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__A2
timestamp 1698431365
transform 1 0 25648 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A1
timestamp 1698431365
transform -1 0 17248 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A2
timestamp 1698431365
transform 1 0 21392 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A2
timestamp 1698431365
transform -1 0 18256 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A2
timestamp 1698431365
transform 1 0 19040 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A1
timestamp 1698431365
transform -1 0 7056 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A2
timestamp 1698431365
transform 1 0 7616 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__I
timestamp 1698431365
transform 1 0 7504 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__I
timestamp 1698431365
transform 1 0 7280 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__I
timestamp 1698431365
transform -1 0 5376 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__I
timestamp 1698431365
transform 1 0 7952 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A2
timestamp 1698431365
transform -1 0 9296 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__A2
timestamp 1698431365
transform 1 0 6608 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__I
timestamp 1698431365
transform 1 0 11872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__I
timestamp 1698431365
transform 1 0 21168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__I
timestamp 1698431365
transform 1 0 21728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__I
timestamp 1698431365
transform 1 0 38864 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__I
timestamp 1698431365
transform -1 0 39648 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1510__I
timestamp 1698431365
transform 1 0 21168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A1
timestamp 1698431365
transform -1 0 22288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1698431365
transform -1 0 26320 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1698431365
transform 1 0 21952 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 22400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A1
timestamp 1698431365
transform 1 0 28000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__B2
timestamp 1698431365
transform 1 0 23072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A1
timestamp 1698431365
transform 1 0 25536 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__I
timestamp 1698431365
transform 1 0 39536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__I
timestamp 1698431365
transform 1 0 38864 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A2
timestamp 1698431365
transform 1 0 29232 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A1
timestamp 1698431365
transform 1 0 29680 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__B2
timestamp 1698431365
transform 1 0 22624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A1
timestamp 1698431365
transform 1 0 26096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__B2
timestamp 1698431365
transform 1 0 29232 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__C2
timestamp 1698431365
transform -1 0 23520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__I
timestamp 1698431365
transform -1 0 10528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__I
timestamp 1698431365
transform 1 0 26432 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1698431365
transform 1 0 29792 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__B2
timestamp 1698431365
transform 1 0 30240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__C2
timestamp 1698431365
transform -1 0 23520 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__I
timestamp 1698431365
transform 1 0 15344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__I
timestamp 1698431365
transform 1 0 27104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__I
timestamp 1698431365
transform 1 0 15232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__I
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__I
timestamp 1698431365
transform -1 0 39648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A1
timestamp 1698431365
transform 1 0 27776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A2
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__B2
timestamp 1698431365
transform 1 0 23744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A1
timestamp 1698431365
transform 1 0 26096 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__I
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A1
timestamp 1698431365
transform 1 0 22176 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A2
timestamp 1698431365
transform -1 0 19712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A1
timestamp 1698431365
transform -1 0 19488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1698431365
transform -1 0 18256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__I
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__I
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A1
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1698431365
transform 1 0 22736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__B
timestamp 1698431365
transform 1 0 22288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A1
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A2
timestamp 1698431365
transform -1 0 27776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__B2
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__I
timestamp 1698431365
transform -1 0 36960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__I0
timestamp 1698431365
transform 1 0 27776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__I1
timestamp 1698431365
transform 1 0 28224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__I2
timestamp 1698431365
transform 1 0 28672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__I3
timestamp 1698431365
transform 1 0 22624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__S0
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__S1
timestamp 1698431365
transform -1 0 22400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__I
timestamp 1698431365
transform 1 0 47040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__I0
timestamp 1698431365
transform 1 0 26320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__I1
timestamp 1698431365
transform 1 0 26544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__I2
timestamp 1698431365
transform 1 0 25872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__I3
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__S0
timestamp 1698431365
transform -1 0 21504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__S1
timestamp 1698431365
transform 1 0 26768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__I
timestamp 1698431365
transform -1 0 47264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A1
timestamp 1698431365
transform -1 0 18592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A2
timestamp 1698431365
transform 1 0 20608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A1
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A2
timestamp 1698431365
transform -1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__I0
timestamp 1698431365
transform 1 0 15120 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__I1
timestamp 1698431365
transform -1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__I3
timestamp 1698431365
transform 1 0 15680 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__S0
timestamp 1698431365
transform -1 0 20832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__S1
timestamp 1698431365
transform 1 0 19712 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__I
timestamp 1698431365
transform -1 0 47264 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__I
timestamp 1698431365
transform -1 0 19040 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A1
timestamp 1698431365
transform -1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A2
timestamp 1698431365
transform 1 0 18368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A1
timestamp 1698431365
transform -1 0 17696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A1
timestamp 1698431365
transform 1 0 18032 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A2
timestamp 1698431365
transform 1 0 19376 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A1
timestamp 1698431365
transform 1 0 17584 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1698431365
transform -1 0 18704 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A1
timestamp 1698431365
transform -1 0 17808 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A1
timestamp 1698431365
transform 1 0 22176 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__B2
timestamp 1698431365
transform 1 0 25312 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__B2
timestamp 1698431365
transform 1 0 26992 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__B2
timestamp 1698431365
transform -1 0 23968 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__I
timestamp 1698431365
transform -1 0 17248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1698431365
transform 1 0 8176 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A1
timestamp 1698431365
transform 1 0 5376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A3
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A4
timestamp 1698431365
transform 1 0 11088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A2
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A3
timestamp 1698431365
transform -1 0 6384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A3
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A4
timestamp 1698431365
transform 1 0 8960 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A2
timestamp 1698431365
transform 1 0 8512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A3
timestamp 1698431365
transform 1 0 8064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A2
timestamp 1698431365
transform 1 0 4480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A3
timestamp 1698431365
transform 1 0 4928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A1
timestamp 1698431365
transform -1 0 5600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A1
timestamp 1698431365
transform 1 0 6048 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform -1 0 5600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A3
timestamp 1698431365
transform 1 0 10080 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A4
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__I
timestamp 1698431365
transform 1 0 6160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform 1 0 8736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698431365
transform 1 0 31696 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A2
timestamp 1698431365
transform 1 0 30576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1698431365
transform 1 0 9968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A1
timestamp 1698431365
transform 1 0 31248 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A2
timestamp 1698431365
transform 1 0 30128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__I
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A2
timestamp 1698431365
transform 1 0 7392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A3
timestamp 1698431365
transform 1 0 9744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A2
timestamp 1698431365
transform 1 0 8624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A3
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1698431365
transform 1 0 18032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A2
timestamp 1698431365
transform 1 0 28560 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__I
timestamp 1698431365
transform 1 0 30688 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A2
timestamp 1698431365
transform 1 0 41664 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__I
timestamp 1698431365
transform -1 0 32928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A1
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A2
timestamp 1698431365
transform 1 0 39648 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__I
timestamp 1698431365
transform 1 0 38080 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A1
timestamp 1698431365
transform 1 0 40544 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A2
timestamp 1698431365
transform -1 0 41216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__I
timestamp 1698431365
transform 1 0 38976 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__I
timestamp 1698431365
transform 1 0 39088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__I
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A2
timestamp 1698431365
transform 1 0 37856 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__B1
timestamp 1698431365
transform 1 0 38528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__I
timestamp 1698431365
transform -1 0 35728 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A3
timestamp 1698431365
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A4
timestamp 1698431365
transform 1 0 39872 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1698431365
transform 1 0 29232 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A1
timestamp 1698431365
transform -1 0 19152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A2
timestamp 1698431365
transform 1 0 20272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__B2
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A2
timestamp 1698431365
transform 1 0 17360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1698431365
transform 1 0 9296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A3
timestamp 1698431365
transform 1 0 5712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A2
timestamp 1698431365
transform -1 0 4368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A3
timestamp 1698431365
transform 1 0 4592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A2
timestamp 1698431365
transform 1 0 5712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1698431365
transform 1 0 28784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__I
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__I
timestamp 1698431365
transform 1 0 37968 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A1
timestamp 1698431365
transform 1 0 42000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A2
timestamp 1698431365
transform 1 0 41552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1698431365
transform 1 0 37520 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__I
timestamp 1698431365
transform 1 0 30576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1698431365
transform -1 0 27328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1698431365
transform 1 0 14112 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A1
timestamp 1698431365
transform 1 0 15344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A1
timestamp 1698431365
transform 1 0 11984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A1
timestamp 1698431365
transform 1 0 5936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__B2
timestamp 1698431365
transform -1 0 8064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A2
timestamp 1698431365
transform -1 0 8624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A1
timestamp 1698431365
transform 1 0 8848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A1
timestamp 1698431365
transform 1 0 6720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A1
timestamp 1698431365
transform 1 0 12544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A1
timestamp 1698431365
transform -1 0 41216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__I
timestamp 1698431365
transform 1 0 39312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A2
timestamp 1698431365
transform -1 0 39760 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1698431365
transform 1 0 39872 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A2
timestamp 1698431365
transform -1 0 41328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A1
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A1
timestamp 1698431365
transform 1 0 41888 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A1
timestamp 1698431365
transform 1 0 40544 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A1
timestamp 1698431365
transform 1 0 24640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A1
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A1
timestamp 1698431365
transform 1 0 11760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A2
timestamp 1698431365
transform 1 0 7056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1698431365
transform 1 0 11424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A2
timestamp 1698431365
transform 1 0 43344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A1
timestamp 1698431365
transform 1 0 42000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A2
timestamp 1698431365
transform 1 0 41216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A1
timestamp 1698431365
transform 1 0 40992 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A2
timestamp 1698431365
transform 1 0 40656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A1
timestamp 1698431365
transform 1 0 39536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A2
timestamp 1698431365
transform 1 0 41552 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A1
timestamp 1698431365
transform 1 0 42448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__I
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A2
timestamp 1698431365
transform 1 0 42784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A1
timestamp 1698431365
transform 1 0 42224 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A1
timestamp 1698431365
transform 1 0 25424 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1698431365
transform 1 0 27104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__I
timestamp 1698431365
transform 1 0 42896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A2
timestamp 1698431365
transform -1 0 38416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__I
timestamp 1698431365
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A2
timestamp 1698431365
transform 1 0 9744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__I
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__A2
timestamp 1698431365
transform 1 0 41888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__I
timestamp 1698431365
transform 1 0 38864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A1
timestamp 1698431365
transform -1 0 41216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A2
timestamp 1698431365
transform 1 0 41552 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__A2
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__I
timestamp 1698431365
transform 1 0 41664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A1
timestamp 1698431365
transform 1 0 37968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A2
timestamp 1698431365
transform 1 0 38416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A1
timestamp 1698431365
transform 1 0 42224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1698431365
transform 1 0 42672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A2
timestamp 1698431365
transform 1 0 42224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__A2
timestamp 1698431365
transform 1 0 43680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A1
timestamp 1698431365
transform 1 0 25424 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A2
timestamp 1698431365
transform 1 0 27776 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1698431365
transform -1 0 28448 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1698431365
transform -1 0 28000 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__A2
timestamp 1698431365
transform -1 0 45472 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A2
timestamp 1698431365
transform 1 0 45248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A2
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__I
timestamp 1698431365
transform 1 0 34944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__I
timestamp 1698431365
transform 1 0 34496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A2
timestamp 1698431365
transform -1 0 42336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1698431365
transform 1 0 39984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A2
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A1
timestamp 1698431365
transform 1 0 38416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__B2
timestamp 1698431365
transform 1 0 22064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__A2
timestamp 1698431365
transform 1 0 21280 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1698431365
transform -1 0 11200 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A2
timestamp 1698431365
transform -1 0 9296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__B
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A2
timestamp 1698431365
transform -1 0 12992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A1
timestamp 1698431365
transform 1 0 16128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A1
timestamp 1698431365
transform -1 0 14000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A1
timestamp 1698431365
transform 1 0 37184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A2
timestamp 1698431365
transform 1 0 38416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1698431365
transform 1 0 37856 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A1
timestamp 1698431365
transform 1 0 25312 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A2
timestamp 1698431365
transform 1 0 28000 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__I
timestamp 1698431365
transform 1 0 11088 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__A1
timestamp 1698431365
transform 1 0 28448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__A2
timestamp 1698431365
transform 1 0 28000 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__A2
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__I
timestamp 1698431365
transform 1 0 39312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A2
timestamp 1698431365
transform 1 0 41216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__A2
timestamp 1698431365
transform 1 0 39088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__I
timestamp 1698431365
transform -1 0 38864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__A1
timestamp 1698431365
transform 1 0 40992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A2
timestamp 1698431365
transform -1 0 21616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A2
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A1
timestamp 1698431365
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A1
timestamp 1698431365
transform -1 0 14112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__A2
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__A2
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__I
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A1
timestamp 1698431365
transform 1 0 26992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A2
timestamp 1698431365
transform 1 0 29232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A3
timestamp 1698431365
transform -1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__A2
timestamp 1698431365
transform 1 0 27664 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__I
timestamp 1698431365
transform -1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A1
timestamp 1698431365
transform 1 0 29008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A2
timestamp 1698431365
transform 1 0 29456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A1
timestamp 1698431365
transform 1 0 27664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__A2
timestamp 1698431365
transform 1 0 26656 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A1
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A2
timestamp 1698431365
transform 1 0 47712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A1
timestamp 1698431365
transform 1 0 43680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__A2
timestamp 1698431365
transform 1 0 41552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__A1
timestamp 1698431365
transform 1 0 40096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__A2
timestamp 1698431365
transform -1 0 38864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1698431365
transform -1 0 22288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A2
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A1
timestamp 1698431365
transform 1 0 16240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A2
timestamp 1698431365
transform 1 0 15008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__A1
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__A2
timestamp 1698431365
transform -1 0 21168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A2
timestamp 1698431365
transform 1 0 20384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A2
timestamp 1698431365
transform 1 0 20048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2215__I
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A1
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A1
timestamp 1698431365
transform 1 0 26432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A2
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A3
timestamp 1698431365
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__A2
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__A2
timestamp 1698431365
transform -1 0 27216 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__A1
timestamp 1698431365
transform 1 0 29120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__A2
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__A1
timestamp 1698431365
transform -1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__A1
timestamp 1698431365
transform -1 0 46480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A1
timestamp 1698431365
transform -1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1698431365
transform 1 0 39088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__A1
timestamp 1698431365
transform 1 0 26544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__A2
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A1
timestamp 1698431365
transform -1 0 16016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A2
timestamp 1698431365
transform -1 0 20272 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2273__A1
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__I
timestamp 1698431365
transform -1 0 34272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1698431365
transform 1 0 27552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__A1
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A1
timestamp 1698431365
transform 1 0 39648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A2
timestamp 1698431365
transform 1 0 38304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A2
timestamp 1698431365
transform -1 0 28448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__I
timestamp 1698431365
transform -1 0 6608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2295__A1
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2295__A2
timestamp 1698431365
transform -1 0 26208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2306__A2
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A1
timestamp 1698431365
transform 1 0 37408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A2
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2324__A1
timestamp 1698431365
transform 1 0 28112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A1
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A2
timestamp 1698431365
transform -1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2337__A2
timestamp 1698431365
transform -1 0 29120 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__I
timestamp 1698431365
transform -1 0 4816 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A1
timestamp 1698431365
transform 1 0 24192 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__A1
timestamp 1698431365
transform 1 0 7728 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__A3
timestamp 1698431365
transform 1 0 6608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2342__A2
timestamp 1698431365
transform -1 0 6384 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A1
timestamp 1698431365
transform -1 0 6272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A1
timestamp 1698431365
transform 1 0 6832 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A3
timestamp 1698431365
transform 1 0 5936 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A3
timestamp 1698431365
transform 1 0 9632 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__A1
timestamp 1698431365
transform -1 0 6608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A1
timestamp 1698431365
transform -1 0 7952 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A1
timestamp 1698431365
transform 1 0 6160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A1
timestamp 1698431365
transform 1 0 6720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__I
timestamp 1698431365
transform 1 0 4816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2358__A1
timestamp 1698431365
transform -1 0 3696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A2
timestamp 1698431365
transform 1 0 5712 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A1
timestamp 1698431365
transform 1 0 5488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__A1
timestamp 1698431365
transform -1 0 3920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__A1
timestamp 1698431365
transform 1 0 3808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__A3
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A1
timestamp 1698431365
transform -1 0 7616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1698431365
transform -1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A1
timestamp 1698431365
transform -1 0 5488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__A1
timestamp 1698431365
transform -1 0 6944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__A2
timestamp 1698431365
transform 1 0 8624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1698431365
transform 1 0 7168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__A2
timestamp 1698431365
transform -1 0 34720 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2394__A2
timestamp 1698431365
transform 1 0 33488 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A2
timestamp 1698431365
transform 1 0 34272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1698431365
transform -1 0 31360 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__A2
timestamp 1698431365
transform -1 0 34608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A2
timestamp 1698431365
transform 1 0 36288 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__A2
timestamp 1698431365
transform 1 0 33936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2414__A1
timestamp 1698431365
transform 1 0 31696 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2417__A1
timestamp 1698431365
transform 1 0 34048 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A1
timestamp 1698431365
transform 1 0 34160 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__I
timestamp 1698431365
transform -1 0 35840 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__A2
timestamp 1698431365
transform 1 0 38976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A2
timestamp 1698431365
transform 1 0 36512 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A2
timestamp 1698431365
transform 1 0 33712 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A2
timestamp 1698431365
transform 1 0 33600 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A1
timestamp 1698431365
transform 1 0 35168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1698431365
transform 1 0 39536 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A2
timestamp 1698431365
transform -1 0 34944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A2
timestamp 1698431365
transform 1 0 32368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2468__A2
timestamp 1698431365
transform 1 0 33936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform -1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__A2
timestamp 1698431365
transform 1 0 39088 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__A1
timestamp 1698431365
transform -1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A1
timestamp 1698431365
transform 1 0 29792 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A2
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1698431365
transform -1 0 31360 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A2
timestamp 1698431365
transform 1 0 29344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A2
timestamp 1698431365
transform -1 0 29680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A2
timestamp 1698431365
transform 1 0 34384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A2
timestamp 1698431365
transform 1 0 34048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1698431365
transform 1 0 34608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A2
timestamp 1698431365
transform 1 0 35168 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__A2
timestamp 1698431365
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__A2
timestamp 1698431365
transform 1 0 35616 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1698431365
transform -1 0 28000 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A2
timestamp 1698431365
transform -1 0 31920 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A3
timestamp 1698431365
transform 1 0 31024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A1
timestamp 1698431365
transform 1 0 30576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A2
timestamp 1698431365
transform 1 0 31024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1698431365
transform -1 0 30800 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1698431365
transform 1 0 29792 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A2
timestamp 1698431365
transform 1 0 30240 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2524__A1
timestamp 1698431365
transform -1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__A1
timestamp 1698431365
transform 1 0 39200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A2
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A2
timestamp 1698431365
transform -1 0 32144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__A2
timestamp 1698431365
transform -1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__A2
timestamp 1698431365
transform -1 0 36624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__A1
timestamp 1698431365
transform -1 0 29008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__A3
timestamp 1698431365
transform -1 0 32032 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A1
timestamp 1698431365
transform 1 0 28896 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A1
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A2
timestamp 1698431365
transform 1 0 38416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A3
timestamp 1698431365
transform 1 0 40320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__A2
timestamp 1698431365
transform 1 0 26096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__B
timestamp 1698431365
transform -1 0 30240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__A2
timestamp 1698431365
transform -1 0 31024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A2
timestamp 1698431365
transform -1 0 35056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A2
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A2
timestamp 1698431365
transform -1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__A2
timestamp 1698431365
transform 1 0 36064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__A1
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__B
timestamp 1698431365
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__A3
timestamp 1698431365
transform -1 0 31248 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__A1
timestamp 1698431365
transform -1 0 31584 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__I
timestamp 1698431365
transform -1 0 26096 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__A1
timestamp 1698431365
transform -1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__B
timestamp 1698431365
transform -1 0 30016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__I
timestamp 1698431365
transform 1 0 18480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__A1
timestamp 1698431365
transform 1 0 34384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__A1
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__B
timestamp 1698431365
transform 1 0 30912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__A1
timestamp 1698431365
transform 1 0 31136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__A2
timestamp 1698431365
transform 1 0 30128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__A1
timestamp 1698431365
transform -1 0 32592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A2
timestamp 1698431365
transform 1 0 32368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A3
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__A2
timestamp 1698431365
transform -1 0 36624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__A1
timestamp 1698431365
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A2
timestamp 1698431365
transform 1 0 36736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A1
timestamp 1698431365
transform 1 0 27216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__I
timestamp 1698431365
transform 1 0 28448 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__A1
timestamp 1698431365
transform -1 0 27104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A1
timestamp 1698431365
transform -1 0 34272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A1
timestamp 1698431365
transform 1 0 34160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__B
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__A1
timestamp 1698431365
transform 1 0 25984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__A1
timestamp 1698431365
transform -1 0 25088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__A1
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__A2
timestamp 1698431365
transform 1 0 29904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__A1
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__I
timestamp 1698431365
transform -1 0 20832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__A1
timestamp 1698431365
transform 1 0 26880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A1
timestamp 1698431365
transform 1 0 30240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A2
timestamp 1698431365
transform 1 0 29792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__A1
timestamp 1698431365
transform 1 0 29344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__B
timestamp 1698431365
transform -1 0 30688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__I0
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__I1
timestamp 1698431365
transform 1 0 32032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__A1
timestamp 1698431365
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__A2
timestamp 1698431365
transform -1 0 19040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__I
timestamp 1698431365
transform -1 0 19040 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__A1
timestamp 1698431365
transform 1 0 20944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A1
timestamp 1698431365
transform 1 0 2912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A2
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__I
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__A1
timestamp 1698431365
transform -1 0 2016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__A2
timestamp 1698431365
transform 1 0 4704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__C
timestamp 1698431365
transform -1 0 3584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__A1
timestamp 1698431365
transform 1 0 3360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__A2
timestamp 1698431365
transform -1 0 2016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__A1
timestamp 1698431365
transform 1 0 3808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__A2
timestamp 1698431365
transform 1 0 3808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__C
timestamp 1698431365
transform 1 0 4256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__A1
timestamp 1698431365
transform 1 0 21392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__A2
timestamp 1698431365
transform 1 0 19264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__I
timestamp 1698431365
transform -1 0 10976 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A1
timestamp 1698431365
transform 1 0 11424 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A1
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__A1
timestamp 1698431365
transform 1 0 19600 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2738__A1
timestamp 1698431365
transform 1 0 7280 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2738__A2
timestamp 1698431365
transform -1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__I
timestamp 1698431365
transform -1 0 15344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__B
timestamp 1698431365
transform 1 0 10528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__A1
timestamp 1698431365
transform 1 0 10528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A1
timestamp 1698431365
transform 1 0 10528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A2
timestamp 1698431365
transform 1 0 10976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__B
timestamp 1698431365
transform 1 0 10304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__I
timestamp 1698431365
transform 1 0 3584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__I
timestamp 1698431365
transform 1 0 4704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__A1
timestamp 1698431365
transform 1 0 2352 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2748__C
timestamp 1698431365
transform -1 0 2016 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__A1
timestamp 1698431365
transform 1 0 8400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2750__A1
timestamp 1698431365
transform 1 0 7504 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2750__A2
timestamp 1698431365
transform -1 0 8176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__B
timestamp 1698431365
transform 1 0 10304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2752__A1
timestamp 1698431365
transform 1 0 2912 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2753__I
timestamp 1698431365
transform -1 0 9408 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__I
timestamp 1698431365
transform 1 0 11648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__A1
timestamp 1698431365
transform -1 0 3808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2758__A1
timestamp 1698431365
transform -1 0 2016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A1
timestamp 1698431365
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A2
timestamp 1698431365
transform -1 0 10304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__A1
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2762__A1
timestamp 1698431365
transform 1 0 19712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__A1
timestamp 1698431365
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__A2
timestamp 1698431365
transform -1 0 10640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__I
timestamp 1698431365
transform 1 0 11088 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__A2
timestamp 1698431365
transform 1 0 9744 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__C
timestamp 1698431365
transform -1 0 10192 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2770__A1
timestamp 1698431365
transform 1 0 11200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__A1
timestamp 1698431365
transform 1 0 11872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__C
timestamp 1698431365
transform -1 0 11424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2772__A1
timestamp 1698431365
transform 1 0 12320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__A1
timestamp 1698431365
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__C
timestamp 1698431365
transform -1 0 11872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2775__A1
timestamp 1698431365
transform -1 0 19040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__A1
timestamp 1698431365
transform -1 0 15344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2778__B
timestamp 1698431365
transform 1 0 17136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__A1
timestamp 1698431365
transform -1 0 16016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2780__A1
timestamp 1698431365
transform -1 0 15456 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2782__I
timestamp 1698431365
transform 1 0 15232 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2783__B
timestamp 1698431365
transform 1 0 16352 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2784__A1
timestamp 1698431365
transform 1 0 14560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A1
timestamp 1698431365
transform 1 0 13216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__C
timestamp 1698431365
transform 1 0 12320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2786__A1
timestamp 1698431365
transform 1 0 14112 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2787__I
timestamp 1698431365
transform 1 0 13440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__A1
timestamp 1698431365
transform -1 0 15344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__C
timestamp 1698431365
transform -1 0 15120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2789__A1
timestamp 1698431365
transform -1 0 17920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__A1
timestamp 1698431365
transform 1 0 15008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__B
timestamp 1698431365
transform 1 0 17808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2792__A1
timestamp 1698431365
transform -1 0 16464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2793__A1
timestamp 1698431365
transform 1 0 16016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2794__B
timestamp 1698431365
transform 1 0 17472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2795__A1
timestamp 1698431365
transform -1 0 18256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2797__I
timestamp 1698431365
transform 1 0 14784 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A1
timestamp 1698431365
transform 1 0 13104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2801__A1
timestamp 1698431365
transform 1 0 10864 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2802__B
timestamp 1698431365
transform -1 0 14336 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2803__A1
timestamp 1698431365
transform 1 0 12544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2804__A1
timestamp 1698431365
transform 1 0 10304 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2805__I
timestamp 1698431365
transform -1 0 14784 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2807__A1
timestamp 1698431365
transform -1 0 11984 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2808__A1
timestamp 1698431365
transform 1 0 10752 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2810__A1
timestamp 1698431365
transform 1 0 12992 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2811__A1
timestamp 1698431365
transform 1 0 10864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2813__I
timestamp 1698431365
transform 1 0 17584 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2816__A1
timestamp 1698431365
transform -1 0 16912 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2818__A1
timestamp 1698431365
transform 1 0 23296 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2819__A1
timestamp 1698431365
transform 1 0 19376 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2820__I
timestamp 1698431365
transform 1 0 24864 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2823__A1
timestamp 1698431365
transform 1 0 18816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2826__A1
timestamp 1698431365
transform 1 0 18256 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__A1
timestamp 1698431365
transform 1 0 23072 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2836__A1
timestamp 1698431365
transform 1 0 23520 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2837__I
timestamp 1698431365
transform 1 0 24528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2839__A1
timestamp 1698431365
transform -1 0 23296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2840__A1
timestamp 1698431365
transform 1 0 23184 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2842__A1
timestamp 1698431365
transform 1 0 28112 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2843__A1
timestamp 1698431365
transform 1 0 21392 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2846__A1
timestamp 1698431365
transform -1 0 25536 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2848__A1
timestamp 1698431365
transform 1 0 21392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2850__A1
timestamp 1698431365
transform -1 0 24304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2851__A1
timestamp 1698431365
transform 1 0 22176 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2855__A1
timestamp 1698431365
transform 1 0 26768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__A1
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2858__A1
timestamp 1698431365
transform -1 0 25648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2859__A1
timestamp 1698431365
transform -1 0 22400 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2861__I
timestamp 1698431365
transform 1 0 15456 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2865__A1
timestamp 1698431365
transform 1 0 13440 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2866__C
timestamp 1698431365
transform -1 0 13776 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2867__A1
timestamp 1698431365
transform -1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2868__A1
timestamp 1698431365
transform 1 0 15904 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2868__C
timestamp 1698431365
transform 1 0 15232 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2869__A1
timestamp 1698431365
transform 1 0 14560 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__C
timestamp 1698431365
transform 1 0 13888 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2871__A1
timestamp 1698431365
transform 1 0 15904 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2872__I
timestamp 1698431365
transform -1 0 14112 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2873__A1
timestamp 1698431365
transform 1 0 15456 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2876__A1
timestamp 1698431365
transform -1 0 16464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2878__A1
timestamp 1698431365
transform -1 0 19824 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2880__A1
timestamp 1698431365
transform -1 0 19936 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__A1
timestamp 1698431365
transform -1 0 17360 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__C
timestamp 1698431365
transform -1 0 18704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2886__A1
timestamp 1698431365
transform 1 0 25648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2890__A1
timestamp 1698431365
transform 1 0 22624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2892__A1
timestamp 1698431365
transform 1 0 26544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A1
timestamp 1698431365
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2896__A1
timestamp 1698431365
transform 1 0 22848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2897__C
timestamp 1698431365
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__A1
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2903__A1
timestamp 1698431365
transform -1 0 23856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2905__A1
timestamp 1698431365
transform 1 0 21728 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__A1
timestamp 1698431365
transform -1 0 26320 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__C
timestamp 1698431365
transform -1 0 24752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2907__A1
timestamp 1698431365
transform -1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2908__A1
timestamp 1698431365
transform 1 0 22848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2910__A1
timestamp 1698431365
transform 1 0 23184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2911__A1
timestamp 1698431365
transform -1 0 21392 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2913__B
timestamp 1698431365
transform -1 0 21952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2919__A1
timestamp 1698431365
transform 1 0 14224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2920__B
timestamp 1698431365
transform -1 0 14896 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2922__A1
timestamp 1698431365
transform 1 0 13776 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2923__B
timestamp 1698431365
transform -1 0 16352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2925__A1
timestamp 1698431365
transform 1 0 12992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__B
timestamp 1698431365
transform -1 0 16800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2928__A1
timestamp 1698431365
transform 1 0 13440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2934__A1
timestamp 1698431365
transform 1 0 11088 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2937__A1
timestamp 1698431365
transform 1 0 12096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2940__A1
timestamp 1698431365
transform 1 0 12544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2943__A1
timestamp 1698431365
transform 1 0 10528 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2944__B
timestamp 1698431365
transform 1 0 11648 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2945__CLK
timestamp 1698431365
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2946__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2947__CLK
timestamp 1698431365
transform 1 0 31472 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2948__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2949__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2950__CLK
timestamp 1698431365
transform 1 0 29232 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2951__CLK
timestamp 1698431365
transform 1 0 22288 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2952__CLK
timestamp 1698431365
transform 1 0 23968 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2953__CLK
timestamp 1698431365
transform 1 0 20496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2954__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2955__CLK
timestamp 1698431365
transform 1 0 17024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2956__CLK
timestamp 1698431365
transform 1 0 16800 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2957__CLK
timestamp 1698431365
transform 1 0 13664 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2958__CLK
timestamp 1698431365
transform 1 0 12432 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2959__CLK
timestamp 1698431365
transform 1 0 10864 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2960__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2960__D
timestamp 1698431365
transform -1 0 9184 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2961__CLK
timestamp 1698431365
transform 1 0 7392 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2962__CLK
timestamp 1698431365
transform 1 0 5712 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2963__CLK
timestamp 1698431365
transform 1 0 7392 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2964__CLK
timestamp 1698431365
transform -1 0 8400 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2965__CLK
timestamp 1698431365
transform 1 0 4592 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2966__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2967__CLK
timestamp 1698431365
transform 1 0 5040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2968__CLK
timestamp 1698431365
transform 1 0 7952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2969__CLK
timestamp 1698431365
transform 1 0 7616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2970__CLK
timestamp 1698431365
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2971__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2972__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2973__CLK
timestamp 1698431365
transform 1 0 8288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3006__CLK
timestamp 1698431365
transform -1 0 24528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3006__D
timestamp 1698431365
transform -1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3021__CLK
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3021__D
timestamp 1698431365
transform 1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3022__CLK
timestamp 1698431365
transform 1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3022__D
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform -1 0 23856 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_clk_I
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_clk_I
timestamp 1698431365
transform 1 0 23184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout73_I
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout78_I
timestamp 1698431365
transform -1 0 3808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout79_I
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout82_I
timestamp 1698431365
transform 1 0 2464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout83_I
timestamp 1698431365
transform 1 0 3808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout84_I
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout85_I
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout95_I
timestamp 1698431365
transform -1 0 3248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout96_I
timestamp 1698431365
transform 1 0 4032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 2800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 14896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 3584 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 1792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 1792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 1792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 2016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 1792 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 1792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 1792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 1792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 1792 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 1792 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 1792 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 1792 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 1792 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 1792 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 2464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 2464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 31024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 10864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 18928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 46480 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 44688 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 42896 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 41440 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 39088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 37520 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 36064 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 33376 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1698431365
transform 1 0 45248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1698431365
transform 1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1698431365
transform 1 0 45920 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1698431365
transform 1 0 46592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1698431365
transform -1 0 46816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1698431365
transform 1 0 46592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output45_I
timestamp 1698431365
transform 1 0 46592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output46_I
timestamp 1698431365
transform -1 0 46816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1698431365
transform -1 0 46816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1698431365
transform -1 0 46928 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1698431365
transform -1 0 46816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698431365
transform -1 0 46816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1698431365
transform -1 0 46816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698431365
transform -1 0 46816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1698431365
transform -1 0 46816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1698431365
transform -1 0 46816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output72_I
timestamp 1698431365
transform -1 0 22176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_rebuffer6_I
timestamp 1698431365
transform 1 0 32144 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23856 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698431365
transform -1 0 13104 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698431365
transform -1 0 22960 0 -1 64288
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout73
timestamp 1698431365
transform 1 0 2016 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout74
timestamp 1698431365
transform -1 0 3136 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout75
timestamp 1698431365
transform -1 0 3360 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout76
timestamp 1698431365
transform 1 0 16016 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout77
timestamp 1698431365
transform 1 0 15344 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout78
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout79
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout80
timestamp 1698431365
transform 1 0 11088 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout81
timestamp 1698431365
transform -1 0 10976 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout82
timestamp 1698431365
transform -1 0 2240 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout83
timestamp 1698431365
transform 1 0 3136 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout84
timestamp 1698431365
transform -1 0 27104 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout85
timestamp 1698431365
transform 1 0 27440 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout86
timestamp 1698431365
transform -1 0 4032 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout87
timestamp 1698431365
transform 1 0 9968 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout88
timestamp 1698431365
transform 1 0 9856 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout89
timestamp 1698431365
transform -1 0 7280 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout90
timestamp 1698431365
transform -1 0 8624 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout91
timestamp 1698431365
transform -1 0 16800 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout92
timestamp 1698431365
transform 1 0 14784 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout93
timestamp 1698431365
transform 1 0 18144 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout94
timestamp 1698431365
transform 1 0 8176 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout95
timestamp 1698431365
transform 1 0 2352 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout96
timestamp 1698431365
transform -1 0 3136 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_10 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_19
timestamp 1698431365
transform 1 0 3472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_27 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_31 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698431365
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_44
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_46
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_55
timestamp 1698431365
transform 1 0 7504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_63
timestamp 1698431365
transform 1 0 8400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_78
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_82
timestamp 1698431365
transform 1 0 10528 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_91
timestamp 1698431365
transform 1 0 11536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_112
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_116
timestamp 1698431365
transform 1 0 14336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_118
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_127
timestamp 1698431365
transform 1 0 15568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_154
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_163
timestamp 1698431365
transform 1 0 19600 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_190
timestamp 1698431365
transform 1 0 22624 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_199
timestamp 1698431365
transform 1 0 23632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_222
timestamp 1698431365
transform 1 0 26208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_226
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_260
timestamp 1698431365
transform 1 0 30464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_262
timestamp 1698431365
transform 1 0 30688 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_324
timestamp 1698431365
transform 1 0 37632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_332
timestamp 1698431365
transform 1 0 38528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_336
timestamp 1698431365
transform 1 0 38976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_350
timestamp 1698431365
transform 1 0 40544 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_366
timestamp 1698431365
transform 1 0 42336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_370
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_384
timestamp 1698431365
transform 1 0 44352 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_404
timestamp 1698431365
transform 1 0 46592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_104
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_106
timestamp 1698431365
transform 1 0 13216 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_121
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_137
timestamp 1698431365
transform 1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_182
timestamp 1698431365
transform 1 0 21728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_192
timestamp 1698431365
transform 1 0 22848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_235
timestamp 1698431365
transform 1 0 27664 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_251
timestamp 1698431365
transform 1 0 29456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_253
timestamp 1698431365
transform 1 0 29680 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_263
timestamp 1698431365
transform 1 0 30800 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_298
timestamp 1698431365
transform 1 0 34720 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_312
timestamp 1698431365
transform 1 0 36288 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_328
timestamp 1698431365
transform 1 0 38080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_344
timestamp 1698431365
transform 1 0 39872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_384
timestamp 1698431365
transform 1 0 44352 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_400
timestamp 1698431365
transform 1 0 46144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_124
timestamp 1698431365
transform 1 0 15232 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_126
timestamp 1698431365
transform 1 0 15456 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_150
timestamp 1698431365
transform 1 0 18144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_214
timestamp 1698431365
transform 1 0 25312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_216
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_240
timestamp 1698431365
transform 1 0 28224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_277
timestamp 1698431365
transform 1 0 32368 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_293
timestamp 1698431365
transform 1 0 34160 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_297
timestamp 1698431365
transform 1 0 34608 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_321
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_331
timestamp 1698431365
transform 1 0 38416 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_355
timestamp 1698431365
transform 1 0 41104 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_371
timestamp 1698431365
transform 1 0 42896 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_379
timestamp 1698431365
transform 1 0 43792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_403
timestamp 1698431365
transform 1 0 46480 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_416
timestamp 1698431365
transform 1 0 47936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_104
timestamp 1698431365
transform 1 0 12992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_121
timestamp 1698431365
transform 1 0 14896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_164
timestamp 1698431365
transform 1 0 19712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_166
timestamp 1698431365
transform 1 0 19936 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_177
timestamp 1698431365
transform 1 0 21168 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_181
timestamp 1698431365
transform 1 0 21616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_224
timestamp 1698431365
transform 1 0 26432 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_263
timestamp 1698431365
transform 1 0 30800 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_267
timestamp 1698431365
transform 1 0 31248 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_344
timestamp 1698431365
transform 1 0 39872 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_356
timestamp 1698431365
transform 1 0 41216 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_374
timestamp 1698431365
transform 1 0 43232 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_406
timestamp 1698431365
transform 1 0 46816 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_414
timestamp 1698431365
transform 1 0 47712 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1698431365
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_135
timestamp 1698431365
transform 1 0 16464 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_143
timestamp 1698431365
transform 1 0 17360 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_147
timestamp 1698431365
transform 1 0 17808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_157
timestamp 1698431365
transform 1 0 18928 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_173
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_193
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_207
timestamp 1698431365
transform 1 0 24528 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_223
timestamp 1698431365
transform 1 0 26320 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_227
timestamp 1698431365
transform 1 0 26768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_229
timestamp 1698431365
transform 1 0 26992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_238
timestamp 1698431365
transform 1 0 28000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_242
timestamp 1698431365
transform 1 0 28448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_259
timestamp 1698431365
transform 1 0 30352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_263
timestamp 1698431365
transform 1 0 30800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_300
timestamp 1698431365
transform 1 0 34944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_310
timestamp 1698431365
transform 1 0 36064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_312
timestamp 1698431365
transform 1 0 36288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_375
timestamp 1698431365
transform 1 0 43344 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_383
timestamp 1698431365
transform 1 0 44240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_403
timestamp 1698431365
transform 1 0 46480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_156
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_164
timestamp 1698431365
transform 1 0 19712 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_185
timestamp 1698431365
transform 1 0 22064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_193
timestamp 1698431365
transform 1 0 22960 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_225
timestamp 1698431365
transform 1 0 26544 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_246
timestamp 1698431365
transform 1 0 28896 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_262
timestamp 1698431365
transform 1 0 30688 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_270
timestamp 1698431365
transform 1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_290
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_322
timestamp 1698431365
transform 1 0 37408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_338
timestamp 1698431365
transform 1 0 39200 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_356
timestamp 1698431365
transform 1 0 41216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_366
timestamp 1698431365
transform 1 0 42336 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_398
timestamp 1698431365
transform 1 0 45920 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_414
timestamp 1698431365
transform 1 0 47712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_115
timestamp 1698431365
transform 1 0 14224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_130
timestamp 1698431365
transform 1 0 15904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_164
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_205
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_229
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_231
timestamp 1698431365
transform 1 0 27216 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_277
timestamp 1698431365
transform 1 0 32368 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_285
timestamp 1698431365
transform 1 0 33264 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_289
timestamp 1698431365
transform 1 0 33712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_291
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_306
timestamp 1698431365
transform 1 0 35616 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_333
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_337
timestamp 1698431365
transform 1 0 39088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_339
timestamp 1698431365
transform 1 0 39312 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_363
timestamp 1698431365
transform 1 0 42000 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_379
timestamp 1698431365
transform 1 0 43792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698431365
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_104
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_134
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_244
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_260
timestamp 1698431365
transform 1 0 30464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_264
timestamp 1698431365
transform 1 0 30912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_273
timestamp 1698431365
transform 1 0 31920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_294
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_296
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_303
timestamp 1698431365
transform 1 0 35280 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_311
timestamp 1698431365
transform 1 0 36176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_315
timestamp 1698431365
transform 1 0 36624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_317
timestamp 1698431365
transform 1 0 36848 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_336
timestamp 1698431365
transform 1 0 38976 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_344
timestamp 1698431365
transform 1 0 39872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_348
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_384
timestamp 1698431365
transform 1 0 44352 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_131
timestamp 1698431365
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_143
timestamp 1698431365
transform 1 0 17360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_147
timestamp 1698431365
transform 1 0 17808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_157
timestamp 1698431365
transform 1 0 18928 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_161
timestamp 1698431365
transform 1 0 19376 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_179
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_188
timestamp 1698431365
transform 1 0 22400 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_204
timestamp 1698431365
transform 1 0 24192 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_208
timestamp 1698431365
transform 1 0 24640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_212
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_216
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_226
timestamp 1698431365
transform 1 0 26656 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_232
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_236
timestamp 1698431365
transform 1 0 27776 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_274
timestamp 1698431365
transform 1 0 32032 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_290
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_292
timestamp 1698431365
transform 1 0 34048 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_307
timestamp 1698431365
transform 1 0 35728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_324
timestamp 1698431365
transform 1 0 37632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_331
timestamp 1698431365
transform 1 0 38416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_358
timestamp 1698431365
transform 1 0 41440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_360
timestamp 1698431365
transform 1 0 41664 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_403
timestamp 1698431365
transform 1 0 46480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_112
timestamp 1698431365
transform 1 0 13888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_202
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_204
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_234
timestamp 1698431365
transform 1 0 27552 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_260
timestamp 1698431365
transform 1 0 30464 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_268
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_272
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_274
timestamp 1698431365
transform 1 0 32032 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_287
timestamp 1698431365
transform 1 0 33488 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_318
timestamp 1698431365
transform 1 0 36960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_344
timestamp 1698431365
transform 1 0 39872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_348
timestamp 1698431365
transform 1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_368
timestamp 1698431365
transform 1 0 42560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_386
timestamp 1698431365
transform 1 0 44576 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_418
timestamp 1698431365
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_85
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_128
timestamp 1698431365
transform 1 0 15680 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_144
timestamp 1698431365
transform 1 0 17472 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_152
timestamp 1698431365
transform 1 0 18368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_162
timestamp 1698431365
transform 1 0 19488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_213
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_215
timestamp 1698431365
transform 1 0 25424 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_252
timestamp 1698431365
transform 1 0 29568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_256
timestamp 1698431365
transform 1 0 30016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_260
timestamp 1698431365
transform 1 0 30464 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_268
timestamp 1698431365
transform 1 0 31360 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_296
timestamp 1698431365
transform 1 0 34496 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_304
timestamp 1698431365
transform 1 0 35392 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_308
timestamp 1698431365
transform 1 0 35840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_327
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_359
timestamp 1698431365
transform 1 0 41552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_369
timestamp 1698431365
transform 1 0 42672 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_96
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_111
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_134
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_168
timestamp 1698431365
transform 1 0 20160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_172
timestamp 1698431365
transform 1 0 20608 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_226
timestamp 1698431365
transform 1 0 26656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_237
timestamp 1698431365
transform 1 0 27888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_241
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_257
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_265
timestamp 1698431365
transform 1 0 31024 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_274
timestamp 1698431365
transform 1 0 32032 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_287
timestamp 1698431365
transform 1 0 33488 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_303
timestamp 1698431365
transform 1 0 35280 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_311
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_315
timestamp 1698431365
transform 1 0 36624 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_383
timestamp 1698431365
transform 1 0 44240 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_399
timestamp 1698431365
transform 1 0 46032 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_403
timestamp 1698431365
transform 1 0 46480 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_93
timestamp 1698431365
transform 1 0 11760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_95
timestamp 1698431365
transform 1 0 11984 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_112
timestamp 1698431365
transform 1 0 13888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_127
timestamp 1698431365
transform 1 0 15568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_143
timestamp 1698431365
transform 1 0 17360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_151
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_165
timestamp 1698431365
transform 1 0 19824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_169
timestamp 1698431365
transform 1 0 20272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_197
timestamp 1698431365
transform 1 0 23408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_199
timestamp 1698431365
transform 1 0 23632 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_218
timestamp 1698431365
transform 1 0 25760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_222
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_283
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_291
timestamp 1698431365
transform 1 0 33936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_295
timestamp 1698431365
transform 1 0 34384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_305
timestamp 1698431365
transform 1 0 35504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_307
timestamp 1698431365
transform 1 0 35728 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_337
timestamp 1698431365
transform 1 0 39088 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_341
timestamp 1698431365
transform 1 0 39536 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_350
timestamp 1698431365
transform 1 0 40544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_376
timestamp 1698431365
transform 1 0 43456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_419
timestamp 1698431365
transform 1 0 48272 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_88
timestamp 1698431365
transform 1 0 11200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_90
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698431365
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_184
timestamp 1698431365
transform 1 0 21952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_193
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_239
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_247
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_263
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_265
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_274
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_296
timestamp 1698431365
transform 1 0 34496 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_309
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_332
timestamp 1698431365
transform 1 0 38528 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_368
timestamp 1698431365
transform 1 0 42560 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_372
timestamp 1698431365
transform 1 0 43008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_397
timestamp 1698431365
transform 1 0 45808 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_413
timestamp 1698431365
transform 1 0 47600 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_69
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_85
timestamp 1698431365
transform 1 0 10864 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_138
timestamp 1698431365
transform 1 0 16800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_140
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_149
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_165
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698431365
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_201
timestamp 1698431365
transform 1 0 23856 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_217
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_221
timestamp 1698431365
transform 1 0 26096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_223
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_230
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_264
timestamp 1698431365
transform 1 0 30912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_268
timestamp 1698431365
transform 1 0 31360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_272
timestamp 1698431365
transform 1 0 31808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_322
timestamp 1698431365
transform 1 0 37408 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_363
timestamp 1698431365
transform 1 0 42000 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_371
timestamp 1698431365
transform 1 0 42896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_375
timestamp 1698431365
transform 1 0 43344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_403
timestamp 1698431365
transform 1 0 46480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_108
timestamp 1698431365
transform 1 0 13440 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_124
timestamp 1698431365
transform 1 0 15232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_132
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_135
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_154
timestamp 1698431365
transform 1 0 18592 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_170
timestamp 1698431365
transform 1 0 20384 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_174
timestamp 1698431365
transform 1 0 20832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_182
timestamp 1698431365
transform 1 0 21728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_195
timestamp 1698431365
transform 1 0 23184 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_225
timestamp 1698431365
transform 1 0 26544 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_257
timestamp 1698431365
transform 1 0 30128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_259
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_262
timestamp 1698431365
transform 1 0 30688 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_300
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_312
timestamp 1698431365
transform 1 0 36288 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_319
timestamp 1698431365
transform 1 0 37072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_326
timestamp 1698431365
transform 1 0 37856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_79
timestamp 1698431365
transform 1 0 10192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_122
timestamp 1698431365
transform 1 0 15008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_126
timestamp 1698431365
transform 1 0 15456 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_158
timestamp 1698431365
transform 1 0 19040 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_192
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_202
timestamp 1698431365
transform 1 0 23968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_204
timestamp 1698431365
transform 1 0 24192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_207
timestamp 1698431365
transform 1 0 24528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_249
timestamp 1698431365
transform 1 0 29232 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_275
timestamp 1698431365
transform 1 0 32144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_279
timestamp 1698431365
transform 1 0 32592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_283
timestamp 1698431365
transform 1 0 33040 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_307
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_353
timestamp 1698431365
transform 1 0 40880 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_367
timestamp 1698431365
transform 1 0 42448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_369
timestamp 1698431365
transform 1 0 42672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_376
timestamp 1698431365
transform 1 0 43456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1698431365
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_399
timestamp 1698431365
transform 1 0 46032 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_407
timestamp 1698431365
transform 1 0 46928 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_416
timestamp 1698431365
transform 1 0 47936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698431365
transform 1 0 10304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698431365
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_91
timestamp 1698431365
transform 1 0 11536 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_107
timestamp 1698431365
transform 1 0 13328 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_148
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_161
timestamp 1698431365
transform 1 0 19376 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_169
timestamp 1698431365
transform 1 0 20272 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_173
timestamp 1698431365
transform 1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_175
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_183
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_187
timestamp 1698431365
transform 1 0 22288 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_203
timestamp 1698431365
transform 1 0 24080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_236
timestamp 1698431365
transform 1 0 27776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_240
timestamp 1698431365
transform 1 0 28224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_242
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_245
timestamp 1698431365
transform 1 0 28784 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_249
timestamp 1698431365
transform 1 0 29232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_294
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_310
timestamp 1698431365
transform 1 0 36064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_312
timestamp 1698431365
transform 1 0 36288 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_315
timestamp 1698431365
transform 1 0 36624 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_331
timestamp 1698431365
transform 1 0 38416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_335
timestamp 1698431365
transform 1 0 38864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_343
timestamp 1698431365
transform 1 0 39760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_347
timestamp 1698431365
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_366
timestamp 1698431365
transform 1 0 42336 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_380
timestamp 1698431365
transform 1 0 43904 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_384
timestamp 1698431365
transform 1 0 44352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_398
timestamp 1698431365
transform 1 0 45920 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_88
timestamp 1698431365
transform 1 0 11200 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_151
timestamp 1698431365
transform 1 0 18256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_160
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_164
timestamp 1698431365
transform 1 0 19712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_209
timestamp 1698431365
transform 1 0 24752 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_211
timestamp 1698431365
transform 1 0 24976 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_269
timestamp 1698431365
transform 1 0 31472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_273
timestamp 1698431365
transform 1 0 31920 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_279
timestamp 1698431365
transform 1 0 32592 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_295
timestamp 1698431365
transform 1 0 34384 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_306
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_321
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_328
timestamp 1698431365
transform 1 0 38080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_332
timestamp 1698431365
transform 1 0 38528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_334
timestamp 1698431365
transform 1 0 38752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_340
timestamp 1698431365
transform 1 0 39424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_344
timestamp 1698431365
transform 1 0 39872 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_348
timestamp 1698431365
transform 1 0 40320 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_356
timestamp 1698431365
transform 1 0 41216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_377
timestamp 1698431365
transform 1 0 43568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_419
timestamp 1698431365
transform 1 0 48272 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_74
timestamp 1698431365
transform 1 0 9632 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_126
timestamp 1698431365
transform 1 0 15456 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_161
timestamp 1698431365
transform 1 0 19376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_163
timestamp 1698431365
transform 1 0 19600 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_177
timestamp 1698431365
transform 1 0 21168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_240
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_249
timestamp 1698431365
transform 1 0 29232 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_253
timestamp 1698431365
transform 1 0 29680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_257
timestamp 1698431365
transform 1 0 30128 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_265
timestamp 1698431365
transform 1 0 31024 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_284
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_293
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_297
timestamp 1698431365
transform 1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_301
timestamp 1698431365
transform 1 0 35056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_303
timestamp 1698431365
transform 1 0 35280 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_317
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_337
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_114
timestamp 1698431365
transform 1 0 14112 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_124
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_156
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_204
timestamp 1698431365
transform 1 0 24192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_218
timestamp 1698431365
transform 1 0 25760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_222
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_281
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_283
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_300
timestamp 1698431365
transform 1 0 34944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_363
timestamp 1698431365
transform 1 0 42000 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_379
timestamp 1698431365
transform 1 0 43792 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_399
timestamp 1698431365
transform 1 0 46032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_403
timestamp 1698431365
transform 1 0 46480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_405
timestamp 1698431365
transform 1 0 46704 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_74
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_114
timestamp 1698431365
transform 1 0 14112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_116
timestamp 1698431365
transform 1 0 14336 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_125
timestamp 1698431365
transform 1 0 15344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698431365
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_160
timestamp 1698431365
transform 1 0 19264 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_174
timestamp 1698431365
transform 1 0 20832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_197
timestamp 1698431365
transform 1 0 23408 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_201
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_203
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_240
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_244
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_248
timestamp 1698431365
transform 1 0 29120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_252
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_358
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_377
timestamp 1698431365
transform 1 0 43568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_381
timestamp 1698431365
transform 1 0 44016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_396
timestamp 1698431365
transform 1 0 45696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_404
timestamp 1698431365
transform 1 0 46592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_22
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_30
timestamp 1698431365
transform 1 0 4704 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_44
timestamp 1698431365
transform 1 0 6272 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_84
timestamp 1698431365
transform 1 0 10752 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_133
timestamp 1698431365
transform 1 0 16240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_135
timestamp 1698431365
transform 1 0 16464 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_149
timestamp 1698431365
transform 1 0 18032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_191
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_207
timestamp 1698431365
transform 1 0 24528 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_286
timestamp 1698431365
transform 1 0 33376 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_302
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_327
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_331
timestamp 1698431365
transform 1 0 38416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_335
timestamp 1698431365
transform 1 0 38864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_339
timestamp 1698431365
transform 1 0 39312 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_347
timestamp 1698431365
transform 1 0 40208 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_351
timestamp 1698431365
transform 1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_368
timestamp 1698431365
transform 1 0 42560 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_399
timestamp 1698431365
transform 1 0 46032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_403
timestamp 1698431365
transform 1 0 46480 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_406
timestamp 1698431365
transform 1 0 46816 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_414
timestamp 1698431365
transform 1 0 47712 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_418
timestamp 1698431365
transform 1 0 48160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_26
timestamp 1698431365
transform 1 0 4256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_30
timestamp 1698431365
transform 1 0 4704 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_60
timestamp 1698431365
transform 1 0 8064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_81
timestamp 1698431365
transform 1 0 10416 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_92
timestamp 1698431365
transform 1 0 11648 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_114
timestamp 1698431365
transform 1 0 14112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_118
timestamp 1698431365
transform 1 0 14560 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_149
timestamp 1698431365
transform 1 0 18032 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_155
timestamp 1698431365
transform 1 0 18704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_163
timestamp 1698431365
transform 1 0 19600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_238
timestamp 1698431365
transform 1 0 28000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_242
timestamp 1698431365
transform 1 0 28448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_263
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_390
timestamp 1698431365
transform 1 0 45024 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_399
timestamp 1698431365
transform 1 0 46032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_403
timestamp 1698431365
transform 1 0 46480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_405
timestamp 1698431365
transform 1 0 46704 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_49
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_58
timestamp 1698431365
transform 1 0 7840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_85
timestamp 1698431365
transform 1 0 10864 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_98
timestamp 1698431365
transform 1 0 12320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_133
timestamp 1698431365
transform 1 0 16240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_135
timestamp 1698431365
transform 1 0 16464 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_147
timestamp 1698431365
transform 1 0 17808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_194
timestamp 1698431365
transform 1 0 23072 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_210
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_228
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_251
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_335
timestamp 1698431365
transform 1 0 38864 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_352
timestamp 1698431365
transform 1 0 40768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_356
timestamp 1698431365
transform 1 0 41216 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_360
timestamp 1698431365
transform 1 0 41664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_371
timestamp 1698431365
transform 1 0 42896 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_379
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_391
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_411
timestamp 1698431365
transform 1 0 47376 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_419
timestamp 1698431365
transform 1 0 48272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_22
timestamp 1698431365
transform 1 0 3808 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_46
timestamp 1698431365
transform 1 0 6496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_85
timestamp 1698431365
transform 1 0 10864 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_122
timestamp 1698431365
transform 1 0 15008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_124
timestamp 1698431365
transform 1 0 15232 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_130
timestamp 1698431365
transform 1 0 15904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_134
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_194
timestamp 1698431365
transform 1 0 23072 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_198
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_246
timestamp 1698431365
transform 1 0 28896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_250
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_332
timestamp 1698431365
transform 1 0 38528 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_357
timestamp 1698431365
transform 1 0 41328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_361
timestamp 1698431365
transform 1 0 41776 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_393
timestamp 1698431365
transform 1 0 45360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_400
timestamp 1698431365
transform 1 0 46144 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_10
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_50
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_66
timestamp 1698431365
transform 1 0 8736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_70
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_72
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_98
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_113
timestamp 1698431365
transform 1 0 14000 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_145
timestamp 1698431365
transform 1 0 17584 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_161
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_189
timestamp 1698431365
transform 1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_227
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_259
timestamp 1698431365
transform 1 0 30352 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_285
timestamp 1698431365
transform 1 0 33264 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_345
timestamp 1698431365
transform 1 0 39984 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_375
timestamp 1698431365
transform 1 0 43344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_377
timestamp 1698431365
transform 1 0 43568 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_380
timestamp 1698431365
transform 1 0 43904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_403
timestamp 1698431365
transform 1 0 46480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_26
timestamp 1698431365
transform 1 0 4256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_38
timestamp 1698431365
transform 1 0 5600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_45
timestamp 1698431365
transform 1 0 6384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_82
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_89
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_97
timestamp 1698431365
transform 1 0 12208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_123
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_153
timestamp 1698431365
transform 1 0 18480 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_176
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_180
timestamp 1698431365
transform 1 0 21504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_188
timestamp 1698431365
transform 1 0 22400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_190
timestamp 1698431365
transform 1 0 22624 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_201
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_224
timestamp 1698431365
transform 1 0 26432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_249
timestamp 1698431365
transform 1 0 29232 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_253
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_257
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_261
timestamp 1698431365
transform 1 0 30576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_297
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_310
timestamp 1698431365
transform 1 0 36064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_329
timestamp 1698431365
transform 1 0 38192 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_333
timestamp 1698431365
transform 1 0 38640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_394
timestamp 1698431365
transform 1 0 45472 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_410
timestamp 1698431365
transform 1 0 47264 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_80
timestamp 1698431365
transform 1 0 10304 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_88
timestamp 1698431365
transform 1 0 11200 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_144
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_146
timestamp 1698431365
transform 1 0 17696 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_160
timestamp 1698431365
transform 1 0 19264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_182
timestamp 1698431365
transform 1 0 21728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_190
timestamp 1698431365
transform 1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_192
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_199
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_207
timestamp 1698431365
transform 1 0 24528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_211
timestamp 1698431365
transform 1 0 24976 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_220
timestamp 1698431365
transform 1 0 25984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_226
timestamp 1698431365
transform 1 0 26656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_230
timestamp 1698431365
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_267
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_281
timestamp 1698431365
transform 1 0 32816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_289
timestamp 1698431365
transform 1 0 33712 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_294
timestamp 1698431365
transform 1 0 34272 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_319
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_322
timestamp 1698431365
transform 1 0 37408 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_338
timestamp 1698431365
transform 1 0 39200 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_342
timestamp 1698431365
transform 1 0 39648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_344
timestamp 1698431365
transform 1 0 39872 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_404
timestamp 1698431365
transform 1 0 46592 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_33
timestamp 1698431365
transform 1 0 5040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_103
timestamp 1698431365
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_179
timestamp 1698431365
transform 1 0 21392 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_183
timestamp 1698431365
transform 1 0 21840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_228
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_251
timestamp 1698431365
transform 1 0 29456 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_259
timestamp 1698431365
transform 1 0 30352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_261
timestamp 1698431365
transform 1 0 30576 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698431365
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698431365
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_326
timestamp 1698431365
transform 1 0 37856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_328
timestamp 1698431365
transform 1 0 38080 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_331
timestamp 1698431365
transform 1 0 38416 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_347
timestamp 1698431365
transform 1 0 40208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_368
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_384
timestamp 1698431365
transform 1 0 44352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_415
timestamp 1698431365
transform 1 0 47824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_22
timestamp 1698431365
transform 1 0 3808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_47
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_50
timestamp 1698431365
transform 1 0 6944 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_54
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_65
timestamp 1698431365
transform 1 0 8624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_73
timestamp 1698431365
transform 1 0 9520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_75
timestamp 1698431365
transform 1 0 9744 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_88
timestamp 1698431365
transform 1 0 11200 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_92
timestamp 1698431365
transform 1 0 11648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_119
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_127
timestamp 1698431365
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_155
timestamp 1698431365
transform 1 0 18704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_159
timestamp 1698431365
transform 1 0 19152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_163
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_179
timestamp 1698431365
transform 1 0 21392 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_218
timestamp 1698431365
transform 1 0 25760 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_234
timestamp 1698431365
transform 1 0 27552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_295
timestamp 1698431365
transform 1 0 34384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_297
timestamp 1698431365
transform 1 0 34608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_358
timestamp 1698431365
transform 1 0 41440 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_374
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_393
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_415
timestamp 1698431365
transform 1 0 47824 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_16
timestamp 1698431365
transform 1 0 3136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_20
timestamp 1698431365
transform 1 0 3584 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_52
timestamp 1698431365
transform 1 0 7168 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_60
timestamp 1698431365
transform 1 0 8064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_62
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_105
timestamp 1698431365
transform 1 0 13104 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_113
timestamp 1698431365
transform 1 0 14000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_115
timestamp 1698431365
transform 1 0 14224 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_122
timestamp 1698431365
transform 1 0 15008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_124
timestamp 1698431365
transform 1 0 15232 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_174
timestamp 1698431365
transform 1 0 20832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_232
timestamp 1698431365
transform 1 0 27328 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_245
timestamp 1698431365
transform 1 0 28784 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_249
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_251
timestamp 1698431365
transform 1 0 29456 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_264
timestamp 1698431365
transform 1 0 30912 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_384
timestamp 1698431365
transform 1 0 44352 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_400
timestamp 1698431365
transform 1 0 46144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_406
timestamp 1698431365
transform 1 0 46816 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_414
timestamp 1698431365
transform 1 0 47712 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1698431365
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_31
timestamp 1698431365
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_43
timestamp 1698431365
transform 1 0 6160 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_59
timestamp 1698431365
transform 1 0 7952 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_67
timestamp 1698431365
transform 1 0 8848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_80
timestamp 1698431365
transform 1 0 10304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_93
timestamp 1698431365
transform 1 0 11760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_97
timestamp 1698431365
transform 1 0 12208 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_122
timestamp 1698431365
transform 1 0 15008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_130
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_132
timestamp 1698431365
transform 1 0 16128 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_138
timestamp 1698431365
transform 1 0 16800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_142
timestamp 1698431365
transform 1 0 17248 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_150
timestamp 1698431365
transform 1 0 18144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_221
timestamp 1698431365
transform 1 0 26096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_225
timestamp 1698431365
transform 1 0 26544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_227
timestamp 1698431365
transform 1 0 26768 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_263
timestamp 1698431365
transform 1 0 30800 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_271
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_275
timestamp 1698431365
transform 1 0 32144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_277
timestamp 1698431365
transform 1 0 32368 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_300
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_319
timestamp 1698431365
transform 1 0 37072 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_343
timestamp 1698431365
transform 1 0 39760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_345
timestamp 1698431365
transform 1 0 39984 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_354
timestamp 1698431365
transform 1 0 40992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_358
timestamp 1698431365
transform 1 0 41440 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_374
timestamp 1698431365
transform 1 0 43232 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_395
timestamp 1698431365
transform 1 0 45584 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_412
timestamp 1698431365
transform 1 0 47488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_10
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_26
timestamp 1698431365
transform 1 0 4256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_30
timestamp 1698431365
transform 1 0 4704 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_33
timestamp 1698431365
transform 1 0 5040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_42
timestamp 1698431365
transform 1 0 6048 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_50
timestamp 1698431365
transform 1 0 6944 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_56
timestamp 1698431365
transform 1 0 7616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_91
timestamp 1698431365
transform 1 0 11536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_98
timestamp 1698431365
transform 1 0 12320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_102
timestamp 1698431365
transform 1 0 12768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_123
timestamp 1698431365
transform 1 0 15120 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_127
timestamp 1698431365
transform 1 0 15568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_135
timestamp 1698431365
transform 1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_152
timestamp 1698431365
transform 1 0 18368 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_159
timestamp 1698431365
transform 1 0 19152 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_167
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_171
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_174
timestamp 1698431365
transform 1 0 20832 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_178
timestamp 1698431365
transform 1 0 21280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_180
timestamp 1698431365
transform 1 0 21504 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_187
timestamp 1698431365
transform 1 0 22288 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_203
timestamp 1698431365
transform 1 0 24080 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_207
timestamp 1698431365
transform 1 0 24528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_259
timestamp 1698431365
transform 1 0 30352 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_267
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_298
timestamp 1698431365
transform 1 0 34720 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_339
timestamp 1698431365
transform 1 0 39312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_343
timestamp 1698431365
transform 1 0 39760 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_347
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_361
timestamp 1698431365
transform 1 0 41776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_365
timestamp 1698431365
transform 1 0 42224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_417
timestamp 1698431365
transform 1 0 48048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_6
timestamp 1698431365
transform 1 0 2016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_16
timestamp 1698431365
transform 1 0 3136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_113
timestamp 1698431365
transform 1 0 14000 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_139
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_200
timestamp 1698431365
transform 1 0 23744 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_216
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_224
timestamp 1698431365
transform 1 0 26432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_228
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_230
timestamp 1698431365
transform 1 0 27104 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_252
timestamp 1698431365
transform 1 0 29568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_256
timestamp 1698431365
transform 1 0 30016 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_264
timestamp 1698431365
transform 1 0 30912 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_268
timestamp 1698431365
transform 1 0 31360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_294
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_302
timestamp 1698431365
transform 1 0 35168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_333
timestamp 1698431365
transform 1 0 38640 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_341
timestamp 1698431365
transform 1 0 39536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_370
timestamp 1698431365
transform 1 0 42784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_378
timestamp 1698431365
transform 1 0 43680 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_54
timestamp 1698431365
transform 1 0 7392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_56
timestamp 1698431365
transform 1 0 7616 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_90
timestamp 1698431365
transform 1 0 11424 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_127
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_155
timestamp 1698431365
transform 1 0 18704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_159
timestamp 1698431365
transform 1 0 19152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_161
timestamp 1698431365
transform 1 0 19376 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_181
timestamp 1698431365
transform 1 0 21616 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_189
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_201
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_220
timestamp 1698431365
transform 1 0 25984 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_341
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_370
timestamp 1698431365
transform 1 0 42784 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_402
timestamp 1698431365
transform 1 0 46368 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_24
timestamp 1698431365
transform 1 0 4032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_62
timestamp 1698431365
transform 1 0 8288 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_66
timestamp 1698431365
transform 1 0 8736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_68
timestamp 1698431365
transform 1 0 8960 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_75
timestamp 1698431365
transform 1 0 9744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_79
timestamp 1698431365
transform 1 0 10192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_81
timestamp 1698431365
transform 1 0 10416 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_99
timestamp 1698431365
transform 1 0 12432 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_154
timestamp 1698431365
transform 1 0 18592 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_170
timestamp 1698431365
transform 1 0 20384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_179
timestamp 1698431365
transform 1 0 21392 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_203
timestamp 1698431365
transform 1 0 24080 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_235
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_276
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_280
timestamp 1698431365
transform 1 0 32704 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_287
timestamp 1698431365
transform 1 0 33488 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_291
timestamp 1698431365
transform 1 0 33936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_293
timestamp 1698431365
transform 1 0 34160 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_333
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_362
timestamp 1698431365
transform 1 0 41888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_366
timestamp 1698431365
transform 1 0 42336 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_371
timestamp 1698431365
transform 1 0 42896 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_379
timestamp 1698431365
transform 1 0 43792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_403
timestamp 1698431365
transform 1 0 46480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_411
timestamp 1698431365
transform 1 0 47376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_415
timestamp 1698431365
transform 1 0 47824 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_18
timestamp 1698431365
transform 1 0 3360 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_24
timestamp 1698431365
transform 1 0 4032 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_28
timestamp 1698431365
transform 1 0 4480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_63
timestamp 1698431365
transform 1 0 8400 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_78
timestamp 1698431365
transform 1 0 10080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_82
timestamp 1698431365
transform 1 0 10528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_84
timestamp 1698431365
transform 1 0 10752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_101
timestamp 1698431365
transform 1 0 12656 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_109
timestamp 1698431365
transform 1 0 13552 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_118
timestamp 1698431365
transform 1 0 14560 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_126
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_148
timestamp 1698431365
transform 1 0 17920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_152
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_159
timestamp 1698431365
transform 1 0 19152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_161
timestamp 1698431365
transform 1 0 19376 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_173
timestamp 1698431365
transform 1 0 20720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_177
timestamp 1698431365
transform 1 0 21168 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_181
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_196
timestamp 1698431365
transform 1 0 23296 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_204
timestamp 1698431365
transform 1 0 24192 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_243
timestamp 1698431365
transform 1 0 28560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_247
timestamp 1698431365
transform 1 0 29008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_249
timestamp 1698431365
transform 1 0 29232 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_267
timestamp 1698431365
transform 1 0 31248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_269
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_305
timestamp 1698431365
transform 1 0 35504 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_313
timestamp 1698431365
transform 1 0 36400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_317
timestamp 1698431365
transform 1 0 36848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_325
timestamp 1698431365
transform 1 0 37744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_327
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_336
timestamp 1698431365
transform 1 0 38976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_358
timestamp 1698431365
transform 1 0 41440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_362
timestamp 1698431365
transform 1 0 41888 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_394
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_416
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_16
timestamp 1698431365
transform 1 0 3136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_20
timestamp 1698431365
transform 1 0 3584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_24
timestamp 1698431365
transform 1 0 4032 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_56
timestamp 1698431365
transform 1 0 7616 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_64
timestamp 1698431365
transform 1 0 8512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_68
timestamp 1698431365
transform 1 0 8960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_86
timestamp 1698431365
transform 1 0 10976 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_94
timestamp 1698431365
transform 1 0 11872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_96
timestamp 1698431365
transform 1 0 12096 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_125
timestamp 1698431365
transform 1 0 15344 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_129
timestamp 1698431365
transform 1 0 15792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_144
timestamp 1698431365
transform 1 0 17472 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_148
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_157
timestamp 1698431365
transform 1 0 18928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_159
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_168
timestamp 1698431365
transform 1 0 20160 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_186
timestamp 1698431365
transform 1 0 22176 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_202
timestamp 1698431365
transform 1 0 23968 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_235
timestamp 1698431365
transform 1 0 27664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_261
timestamp 1698431365
transform 1 0 30576 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_305
timestamp 1698431365
transform 1 0 35504 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_341
timestamp 1698431365
transform 1 0 39536 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_348
timestamp 1698431365
transform 1 0 40320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_359
timestamp 1698431365
transform 1 0 41552 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_363
timestamp 1698431365
transform 1 0 42000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_391
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_393
timestamp 1698431365
transform 1 0 45360 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_418
timestamp 1698431365
transform 1 0 48160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_16
timestamp 1698431365
transform 1 0 3136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_20
timestamp 1698431365
transform 1 0 3584 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_24
timestamp 1698431365
transform 1 0 4032 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_27
timestamp 1698431365
transform 1 0 4368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_92
timestamp 1698431365
transform 1 0 11648 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_101
timestamp 1698431365
transform 1 0 12656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_103
timestamp 1698431365
transform 1 0 12880 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_148
timestamp 1698431365
transform 1 0 17920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_152
timestamp 1698431365
transform 1 0 18368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_162
timestamp 1698431365
transform 1 0 19488 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_222
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_224
timestamp 1698431365
transform 1 0 26432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_227
timestamp 1698431365
transform 1 0 26768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_231
timestamp 1698431365
transform 1 0 27216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_245
timestamp 1698431365
transform 1 0 28784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_249
timestamp 1698431365
transform 1 0 29232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_253
timestamp 1698431365
transform 1 0 29680 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_333
timestamp 1698431365
transform 1 0 38640 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_341
timestamp 1698431365
transform 1 0 39536 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_344
timestamp 1698431365
transform 1 0 39872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_367
timestamp 1698431365
transform 1 0 42448 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_379
timestamp 1698431365
transform 1 0 43792 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_383
timestamp 1698431365
transform 1 0 44240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_385
timestamp 1698431365
transform 1 0 44464 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_399
timestamp 1698431365
transform 1 0 46032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_401
timestamp 1698431365
transform 1 0 46256 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_412
timestamp 1698431365
transform 1 0 47488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_20
timestamp 1698431365
transform 1 0 3584 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_31
timestamp 1698431365
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_69
timestamp 1698431365
transform 1 0 9072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_73
timestamp 1698431365
transform 1 0 9520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_77
timestamp 1698431365
transform 1 0 9968 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_85
timestamp 1698431365
transform 1 0 10864 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_89
timestamp 1698431365
transform 1 0 11312 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_96
timestamp 1698431365
transform 1 0 12096 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_123
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_139
timestamp 1698431365
transform 1 0 16912 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_161
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_182
timestamp 1698431365
transform 1 0 21728 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_221
timestamp 1698431365
transform 1 0 26096 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_259
timestamp 1698431365
transform 1 0 30352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_261
timestamp 1698431365
transform 1 0 30576 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_268
timestamp 1698431365
transform 1 0 31360 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_292
timestamp 1698431365
transform 1 0 34048 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_296
timestamp 1698431365
transform 1 0 34496 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_321
timestamp 1698431365
transform 1 0 37296 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_346
timestamp 1698431365
transform 1 0 40096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_350
timestamp 1698431365
transform 1 0 40544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_377
timestamp 1698431365
transform 1 0 43568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_399
timestamp 1698431365
transform 1 0 46032 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_415
timestamp 1698431365
transform 1 0 47824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_419
timestamp 1698431365
transform 1 0 48272 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_54
timestamp 1698431365
transform 1 0 7392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_56
timestamp 1698431365
transform 1 0 7616 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_84
timestamp 1698431365
transform 1 0 10752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_86
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_93
timestamp 1698431365
transform 1 0 11760 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_133
timestamp 1698431365
transform 1 0 16240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_167
timestamp 1698431365
transform 1 0 20048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_204
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_218
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_221
timestamp 1698431365
transform 1 0 26096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_225
timestamp 1698431365
transform 1 0 26544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_229
timestamp 1698431365
transform 1 0 26992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_231
timestamp 1698431365
transform 1 0 27216 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_234
timestamp 1698431365
transform 1 0 27552 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_238
timestamp 1698431365
transform 1 0 28000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_242
timestamp 1698431365
transform 1 0 28448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_246
timestamp 1698431365
transform 1 0 28896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_248
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_273
timestamp 1698431365
transform 1 0 31920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_377
timestamp 1698431365
transform 1 0 43568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_385
timestamp 1698431365
transform 1 0 44464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_389
timestamp 1698431365
transform 1 0 44912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_391
timestamp 1698431365
transform 1 0 45136 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_408
timestamp 1698431365
transform 1 0 47040 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_10
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_18
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_24
timestamp 1698431365
transform 1 0 4032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_64
timestamp 1698431365
transform 1 0 8512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_68
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_72
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_102
timestamp 1698431365
transform 1 0 12768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_111
timestamp 1698431365
transform 1 0 13776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_121
timestamp 1698431365
transform 1 0 14896 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_137
timestamp 1698431365
transform 1 0 16688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_139
timestamp 1698431365
transform 1 0 16912 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_150
timestamp 1698431365
transform 1 0 18144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_154
timestamp 1698431365
transform 1 0 18592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_156
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_159
timestamp 1698431365
transform 1 0 19152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_161
timestamp 1698431365
transform 1 0 19376 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_167
timestamp 1698431365
transform 1 0 20048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_188
timestamp 1698431365
transform 1 0 22400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_192
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_285
timestamp 1698431365
transform 1 0 33264 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_301
timestamp 1698431365
transform 1 0 35056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_347
timestamp 1698431365
transform 1 0 40208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_349
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_358
timestamp 1698431365
transform 1 0 41440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_362
timestamp 1698431365
transform 1 0 41888 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_378
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698431365
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698431365
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_409
timestamp 1698431365
transform 1 0 47152 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_413
timestamp 1698431365
transform 1 0 47600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_415
timestamp 1698431365
transform 1 0 47824 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_6
timestamp 1698431365
transform 1 0 2016 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_22
timestamp 1698431365
transform 1 0 3808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_24
timestamp 1698431365
transform 1 0 4032 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_54
timestamp 1698431365
transform 1 0 7392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_58
timestamp 1698431365
transform 1 0 7840 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_88
timestamp 1698431365
transform 1 0 11200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_119
timestamp 1698431365
transform 1 0 14672 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_123
timestamp 1698431365
transform 1 0 15120 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_135
timestamp 1698431365
transform 1 0 16464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_146
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_148
timestamp 1698431365
transform 1 0 17920 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_156
timestamp 1698431365
transform 1 0 18816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_158
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_192
timestamp 1698431365
transform 1 0 22848 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_220
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_228
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_232
timestamp 1698431365
transform 1 0 27328 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_259
timestamp 1698431365
transform 1 0 30352 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_302
timestamp 1698431365
transform 1 0 35168 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_318
timestamp 1698431365
transform 1 0 36960 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_365
timestamp 1698431365
transform 1 0 42224 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_369
timestamp 1698431365
transform 1 0 42672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_371
timestamp 1698431365
transform 1 0 42896 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_385
timestamp 1698431365
transform 1 0 44464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_389
timestamp 1698431365
transform 1 0 44912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_6
timestamp 1698431365
transform 1 0 2016 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_14
timestamp 1698431365
transform 1 0 2912 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_18
timestamp 1698431365
transform 1 0 3360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_24
timestamp 1698431365
transform 1 0 4032 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_65
timestamp 1698431365
transform 1 0 8624 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_115
timestamp 1698431365
transform 1 0 14224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_193
timestamp 1698431365
transform 1 0 22960 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_201
timestamp 1698431365
transform 1 0 23856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_205
timestamp 1698431365
transform 1 0 24304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_207
timestamp 1698431365
transform 1 0 24528 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_213
timestamp 1698431365
transform 1 0 25200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_217
timestamp 1698431365
transform 1 0 25648 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_225
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_249
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_258
timestamp 1698431365
transform 1 0 30240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_265
timestamp 1698431365
transform 1 0 31024 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_281
timestamp 1698431365
transform 1 0 32816 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_297
timestamp 1698431365
transform 1 0 34608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_309
timestamp 1698431365
transform 1 0 35952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_336
timestamp 1698431365
transform 1 0 38976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_340
timestamp 1698431365
transform 1 0 39424 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_347
timestamp 1698431365
transform 1 0 40208 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_379
timestamp 1698431365
transform 1 0 43792 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_419
timestamp 1698431365
transform 1 0 48272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_16
timestamp 1698431365
transform 1 0 3136 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_25
timestamp 1698431365
transform 1 0 4144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_33
timestamp 1698431365
transform 1 0 5040 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_35
timestamp 1698431365
transform 1 0 5264 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_101
timestamp 1698431365
transform 1 0 12656 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_117
timestamp 1698431365
transform 1 0 14448 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_137
timestamp 1698431365
transform 1 0 16688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698431365
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_174
timestamp 1698431365
transform 1 0 20832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_176
timestamp 1698431365
transform 1 0 21056 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_179
timestamp 1698431365
transform 1 0 21392 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_181
timestamp 1698431365
transform 1 0 21616 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_184
timestamp 1698431365
transform 1 0 21952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_188
timestamp 1698431365
transform 1 0 22400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_192
timestamp 1698431365
transform 1 0 22848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_194
timestamp 1698431365
transform 1 0 23072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_225
timestamp 1698431365
transform 1 0 26544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_229
timestamp 1698431365
transform 1 0 26992 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_247
timestamp 1698431365
transform 1 0 29008 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_261
timestamp 1698431365
transform 1 0 30576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_265
timestamp 1698431365
transform 1 0 31024 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_273
timestamp 1698431365
transform 1 0 31920 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_277
timestamp 1698431365
transform 1 0 32368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_295
timestamp 1698431365
transform 1 0 34384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_299
timestamp 1698431365
transform 1 0 34832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_301
timestamp 1698431365
transform 1 0 35056 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_304
timestamp 1698431365
transform 1 0 35392 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_344
timestamp 1698431365
transform 1 0 39872 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_348
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_363
timestamp 1698431365
transform 1 0 42000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_367
timestamp 1698431365
transform 1 0 42448 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_380
timestamp 1698431365
transform 1 0 43904 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_412
timestamp 1698431365
transform 1 0 47488 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_43
timestamp 1698431365
transform 1 0 6160 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_85
timestamp 1698431365
transform 1 0 10864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_89
timestamp 1698431365
transform 1 0 11312 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_93
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_96
timestamp 1698431365
transform 1 0 12096 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_136
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_138
timestamp 1698431365
transform 1 0 16800 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_144
timestamp 1698431365
transform 1 0 17472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_148
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_164
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_168
timestamp 1698431365
transform 1 0 20160 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_185
timestamp 1698431365
transform 1 0 22064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_271
timestamp 1698431365
transform 1 0 31696 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_295
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_329
timestamp 1698431365
transform 1 0 38192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_337
timestamp 1698431365
transform 1 0 39088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_349
timestamp 1698431365
transform 1 0 40432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_351
timestamp 1698431365
transform 1 0 40656 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_363
timestamp 1698431365
transform 1 0 42000 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_411
timestamp 1698431365
transform 1 0 47376 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_419
timestamp 1698431365
transform 1 0 48272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_33
timestamp 1698431365
transform 1 0 5040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_35
timestamp 1698431365
transform 1 0 5264 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_80
timestamp 1698431365
transform 1 0 10304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_94
timestamp 1698431365
transform 1 0 11872 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_124
timestamp 1698431365
transform 1 0 15232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_132
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_171
timestamp 1698431365
transform 1 0 20496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_177
timestamp 1698431365
transform 1 0 21168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_202
timestamp 1698431365
transform 1 0 23968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_246
timestamp 1698431365
transform 1 0 28896 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_254
timestamp 1698431365
transform 1 0 29792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_256
timestamp 1698431365
transform 1 0 30016 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_265
timestamp 1698431365
transform 1 0 31024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_275
timestamp 1698431365
transform 1 0 32144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_287
timestamp 1698431365
transform 1 0 33488 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_291
timestamp 1698431365
transform 1 0 33936 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_316
timestamp 1698431365
transform 1 0 36736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_318
timestamp 1698431365
transform 1 0 36960 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_329
timestamp 1698431365
transform 1 0 38192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_342
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_356
timestamp 1698431365
transform 1 0 41216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_363
timestamp 1698431365
transform 1 0 42000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_367
timestamp 1698431365
transform 1 0 42448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_371
timestamp 1698431365
transform 1 0 42896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_373
timestamp 1698431365
transform 1 0 43120 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_400
timestamp 1698431365
transform 1 0 46144 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_18
timestamp 1698431365
transform 1 0 3360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_22
timestamp 1698431365
transform 1 0 3808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_45
timestamp 1698431365
transform 1 0 6384 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_54
timestamp 1698431365
transform 1 0 7392 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_58
timestamp 1698431365
transform 1 0 7840 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_64
timestamp 1698431365
transform 1 0 8512 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_96
timestamp 1698431365
transform 1 0 12096 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_115
timestamp 1698431365
transform 1 0 14224 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_119
timestamp 1698431365
transform 1 0 14672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_121
timestamp 1698431365
transform 1 0 14896 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_145
timestamp 1698431365
transform 1 0 17584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_149
timestamp 1698431365
transform 1 0 18032 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_157
timestamp 1698431365
transform 1 0 18928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_159
timestamp 1698431365
transform 1 0 19152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_181
timestamp 1698431365
transform 1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_183
timestamp 1698431365
transform 1 0 21840 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_186
timestamp 1698431365
transform 1 0 22176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_190
timestamp 1698431365
transform 1 0 22624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_194
timestamp 1698431365
transform 1 0 23072 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_202
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_204
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_210
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_275
timestamp 1698431365
transform 1 0 32144 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_299
timestamp 1698431365
transform 1 0 34832 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_335
timestamp 1698431365
transform 1 0 38864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_357
timestamp 1698431365
transform 1 0 41328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_361
timestamp 1698431365
transform 1 0 41776 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_377
timestamp 1698431365
transform 1 0 43568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_402
timestamp 1698431365
transform 1 0 46368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_28
timestamp 1698431365
transform 1 0 4480 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_35
timestamp 1698431365
transform 1 0 5264 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_39
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_45
timestamp 1698431365
transform 1 0 6384 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_61
timestamp 1698431365
transform 1 0 8176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_67
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_76
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_80
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_86
timestamp 1698431365
transform 1 0 10976 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_90
timestamp 1698431365
transform 1 0 11424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_94
timestamp 1698431365
transform 1 0 11872 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_126
timestamp 1698431365
transform 1 0 15456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_130
timestamp 1698431365
transform 1 0 15904 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_146
timestamp 1698431365
transform 1 0 17696 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_154
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_182
timestamp 1698431365
transform 1 0 21728 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_189
timestamp 1698431365
transform 1 0 22512 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_220
timestamp 1698431365
transform 1 0 25984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_224
timestamp 1698431365
transform 1 0 26432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_254
timestamp 1698431365
transform 1 0 29792 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_262
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_298
timestamp 1698431365
transform 1 0 34720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_312
timestamp 1698431365
transform 1 0 36288 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_330
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_338
timestamp 1698431365
transform 1 0 39200 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_347
timestamp 1698431365
transform 1 0 40208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698431365
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_358
timestamp 1698431365
transform 1 0 41440 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_390
timestamp 1698431365
transform 1 0 45024 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_399
timestamp 1698431365
transform 1 0 46032 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_415
timestamp 1698431365
transform 1 0 47824 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_10
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_43
timestamp 1698431365
transform 1 0 6160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_92
timestamp 1698431365
transform 1 0 11648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_96
timestamp 1698431365
transform 1 0 12096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_100
timestamp 1698431365
transform 1 0 12544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_113
timestamp 1698431365
transform 1 0 14000 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_123
timestamp 1698431365
transform 1 0 15120 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_131
timestamp 1698431365
transform 1 0 16016 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_133
timestamp 1698431365
transform 1 0 16240 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_136
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_152
timestamp 1698431365
transform 1 0 18368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_160
timestamp 1698431365
transform 1 0 19264 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_166
timestamp 1698431365
transform 1 0 19936 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_232
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_236
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_240
timestamp 1698431365
transform 1 0 28224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_287
timestamp 1698431365
transform 1 0 33488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_293
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_297
timestamp 1698431365
transform 1 0 34608 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_305
timestamp 1698431365
transform 1 0 35504 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_309
timestamp 1698431365
transform 1 0 35952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_334
timestamp 1698431365
transform 1 0 38752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_338
timestamp 1698431365
transform 1 0 39200 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_346
timestamp 1698431365
transform 1 0 40096 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_350
timestamp 1698431365
transform 1 0 40544 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_353
timestamp 1698431365
transform 1 0 40880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_355
timestamp 1698431365
transform 1 0 41104 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_358
timestamp 1698431365
transform 1 0 41440 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_379
timestamp 1698431365
transform 1 0 43792 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_395
timestamp 1698431365
transform 1 0 45584 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_408
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_416
timestamp 1698431365
transform 1 0 47936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_16
timestamp 1698431365
transform 1 0 3136 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_22
timestamp 1698431365
transform 1 0 3808 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_104
timestamp 1698431365
transform 1 0 12992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_108
timestamp 1698431365
transform 1 0 13440 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_119
timestamp 1698431365
transform 1 0 14672 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_123
timestamp 1698431365
transform 1 0 15120 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_146
timestamp 1698431365
transform 1 0 17696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_148
timestamp 1698431365
transform 1 0 17920 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_187
timestamp 1698431365
transform 1 0 22288 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_195
timestamp 1698431365
transform 1 0 23184 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_220
timestamp 1698431365
transform 1 0 25984 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_222
timestamp 1698431365
transform 1 0 26208 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_252
timestamp 1698431365
transform 1 0 29568 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_268
timestamp 1698431365
transform 1 0 31360 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_314
timestamp 1698431365
transform 1 0 36512 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_322
timestamp 1698431365
transform 1 0 37408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_324
timestamp 1698431365
transform 1 0 37632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_333
timestamp 1698431365
transform 1 0 38640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_337
timestamp 1698431365
transform 1 0 39088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_341
timestamp 1698431365
transform 1 0 39536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_356
timestamp 1698431365
transform 1 0 41216 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_377
timestamp 1698431365
transform 1 0 43568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_385
timestamp 1698431365
transform 1 0 44464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_389
timestamp 1698431365
transform 1 0 44912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_391
timestamp 1698431365
transform 1 0 45136 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_414
timestamp 1698431365
transform 1 0 47712 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_418
timestamp 1698431365
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_28
timestamp 1698431365
transform 1 0 4480 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_41
timestamp 1698431365
transform 1 0 5936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_54
timestamp 1698431365
transform 1 0 7392 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_121
timestamp 1698431365
transform 1 0 14896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_125
timestamp 1698431365
transform 1 0 15344 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_151
timestamp 1698431365
transform 1 0 18256 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_159
timestamp 1698431365
transform 1 0 19152 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_163
timestamp 1698431365
transform 1 0 19600 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_165
timestamp 1698431365
transform 1 0 19824 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_196
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_205
timestamp 1698431365
transform 1 0 24304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_219
timestamp 1698431365
transform 1 0 25872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_223
timestamp 1698431365
transform 1 0 26320 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_239
timestamp 1698431365
transform 1 0 28112 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_249
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_279
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_287
timestamp 1698431365
transform 1 0 33488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_289
timestamp 1698431365
transform 1 0 33712 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_298
timestamp 1698431365
transform 1 0 34720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_302
timestamp 1698431365
transform 1 0 35168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_310
timestamp 1698431365
transform 1 0 36064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_363
timestamp 1698431365
transform 1 0 42000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_378
timestamp 1698431365
transform 1 0 43680 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_382
timestamp 1698431365
transform 1 0 44128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_395
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_397
timestamp 1698431365
transform 1 0 45808 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_416
timestamp 1698431365
transform 1 0 47936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_18
timestamp 1698431365
transform 1 0 3360 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_22
timestamp 1698431365
transform 1 0 3808 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_64
timestamp 1698431365
transform 1 0 8512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_112
timestamp 1698431365
transform 1 0 13888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_116
timestamp 1698431365
transform 1 0 14336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_120
timestamp 1698431365
transform 1 0 14784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_122
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_130
timestamp 1698431365
transform 1 0 15904 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698431365
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_159
timestamp 1698431365
transform 1 0 19152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_161
timestamp 1698431365
transform 1 0 19376 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_180
timestamp 1698431365
transform 1 0 21504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_184
timestamp 1698431365
transform 1 0 21952 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_188
timestamp 1698431365
transform 1 0 22400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_192
timestamp 1698431365
transform 1 0 22848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_194
timestamp 1698431365
transform 1 0 23072 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_201
timestamp 1698431365
transform 1 0 23856 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_205
timestamp 1698431365
transform 1 0 24304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_207
timestamp 1698431365
transform 1 0 24528 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_251
timestamp 1698431365
transform 1 0 29456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_277
timestamp 1698431365
transform 1 0 32368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_279
timestamp 1698431365
transform 1 0 32592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_290
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_319
timestamp 1698431365
transform 1 0 37072 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_335
timestamp 1698431365
transform 1 0 38864 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_339
timestamp 1698431365
transform 1 0 39312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_361
timestamp 1698431365
transform 1 0 41776 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_365
timestamp 1698431365
transform 1 0 42224 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_381
timestamp 1698431365
transform 1 0 44016 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_385
timestamp 1698431365
transform 1 0 44464 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_391
timestamp 1698431365
transform 1 0 45136 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_399
timestamp 1698431365
transform 1 0 46032 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_415
timestamp 1698431365
transform 1 0 47824 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698431365
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_66
timestamp 1698431365
transform 1 0 8736 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_96
timestamp 1698431365
transform 1 0 12096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_100
timestamp 1698431365
transform 1 0 12544 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_111
timestamp 1698431365
transform 1 0 13776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_139
timestamp 1698431365
transform 1 0 16912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_161
timestamp 1698431365
transform 1 0 19376 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_165
timestamp 1698431365
transform 1 0 19824 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_190
timestamp 1698431365
transform 1 0 22624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_208
timestamp 1698431365
transform 1 0 24640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_212
timestamp 1698431365
transform 1 0 25088 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_220
timestamp 1698431365
transform 1 0 25984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_230
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_238
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_242
timestamp 1698431365
transform 1 0 28448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_253
timestamp 1698431365
transform 1 0 29680 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_260
timestamp 1698431365
transform 1 0 30464 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_276
timestamp 1698431365
transform 1 0 32256 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_308
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_314
timestamp 1698431365
transform 1 0 36512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_333
timestamp 1698431365
transform 1 0 38640 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_341
timestamp 1698431365
transform 1 0 39536 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_343
timestamp 1698431365
transform 1 0 39760 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_346
timestamp 1698431365
transform 1 0 40096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_353
timestamp 1698431365
transform 1 0 40880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_357
timestamp 1698431365
transform 1 0 41328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_361
timestamp 1698431365
transform 1 0 41776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_363
timestamp 1698431365
transform 1 0 42000 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_372
timestamp 1698431365
transform 1 0 43008 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_376
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_411
timestamp 1698431365
transform 1 0 47376 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_419
timestamp 1698431365
transform 1 0 48272 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_10
timestamp 1698431365
transform 1 0 2464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_14
timestamp 1698431365
transform 1 0 2912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_44
timestamp 1698431365
transform 1 0 6272 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_52
timestamp 1698431365
transform 1 0 7168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_54
timestamp 1698431365
transform 1 0 7392 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_57
timestamp 1698431365
transform 1 0 7728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_84
timestamp 1698431365
transform 1 0 10752 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_90
timestamp 1698431365
transform 1 0 11424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_94
timestamp 1698431365
transform 1 0 11872 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_102
timestamp 1698431365
transform 1 0 12768 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_106
timestamp 1698431365
transform 1 0 13216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_116
timestamp 1698431365
transform 1 0 14336 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_132
timestamp 1698431365
transform 1 0 16128 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_147
timestamp 1698431365
transform 1 0 17808 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_158
timestamp 1698431365
transform 1 0 19040 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_166
timestamp 1698431365
transform 1 0 19936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_170
timestamp 1698431365
transform 1 0 20384 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_175
timestamp 1698431365
transform 1 0 20944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_179
timestamp 1698431365
transform 1 0 21392 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_183
timestamp 1698431365
transform 1 0 21840 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_185
timestamp 1698431365
transform 1 0 22064 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_188
timestamp 1698431365
transform 1 0 22400 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_254
timestamp 1698431365
transform 1 0 29792 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_258
timestamp 1698431365
transform 1 0 30240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_264
timestamp 1698431365
transform 1 0 30912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_268
timestamp 1698431365
transform 1 0 31360 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_286
timestamp 1698431365
transform 1 0 33376 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_292
timestamp 1698431365
transform 1 0 34048 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_294
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_302
timestamp 1698431365
transform 1 0 35168 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_318
timestamp 1698431365
transform 1 0 36960 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_326
timestamp 1698431365
transform 1 0 37856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_330
timestamp 1698431365
transform 1 0 38304 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_348
timestamp 1698431365
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_360
timestamp 1698431365
transform 1 0 41664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_370
timestamp 1698431365
transform 1 0 42784 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_374
timestamp 1698431365
transform 1 0 43232 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_387
timestamp 1698431365
transform 1 0 44688 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_403
timestamp 1698431365
transform 1 0 46480 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_12
timestamp 1698431365
transform 1 0 2688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_16
timestamp 1698431365
transform 1 0 3136 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_20
timestamp 1698431365
transform 1 0 3584 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_89
timestamp 1698431365
transform 1 0 11312 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_127
timestamp 1698431365
transform 1 0 15568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_159
timestamp 1698431365
transform 1 0 19152 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_163
timestamp 1698431365
transform 1 0 19600 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_166
timestamp 1698431365
transform 1 0 19936 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_172
timestamp 1698431365
transform 1 0 20608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_174
timestamp 1698431365
transform 1 0 20832 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_191
timestamp 1698431365
transform 1 0 22736 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_197
timestamp 1698431365
transform 1 0 23408 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_201
timestamp 1698431365
transform 1 0 23856 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_215
timestamp 1698431365
transform 1 0 25424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_219
timestamp 1698431365
transform 1 0 25872 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_223
timestamp 1698431365
transform 1 0 26320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_227
timestamp 1698431365
transform 1 0 26768 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_243
timestamp 1698431365
transform 1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_279
timestamp 1698431365
transform 1 0 32592 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_305
timestamp 1698431365
transform 1 0 35504 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_313
timestamp 1698431365
transform 1 0 36400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_327
timestamp 1698431365
transform 1 0 37968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_329
timestamp 1698431365
transform 1 0 38192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_336
timestamp 1698431365
transform 1 0 38976 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_340
timestamp 1698431365
transform 1 0 39424 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_353
timestamp 1698431365
transform 1 0 40880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_379
timestamp 1698431365
transform 1 0 43792 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_383
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_419
timestamp 1698431365
transform 1 0 48272 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_22
timestamp 1698431365
transform 1 0 3808 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_24
timestamp 1698431365
transform 1 0 4032 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_29
timestamp 1698431365
transform 1 0 4592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_33
timestamp 1698431365
transform 1 0 5040 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_41
timestamp 1698431365
transform 1 0 5936 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_62
timestamp 1698431365
transform 1 0 8288 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_80
timestamp 1698431365
transform 1 0 10304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_90
timestamp 1698431365
transform 1 0 11424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_94
timestamp 1698431365
transform 1 0 11872 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_102
timestamp 1698431365
transform 1 0 12768 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_135
timestamp 1698431365
transform 1 0 16464 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1698431365
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_144
timestamp 1698431365
transform 1 0 17472 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_201
timestamp 1698431365
transform 1 0 23856 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_220
timestamp 1698431365
transform 1 0 25984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_222
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_255
timestamp 1698431365
transform 1 0 29904 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_263
timestamp 1698431365
transform 1 0 30800 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_267
timestamp 1698431365
transform 1 0 31248 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_274
timestamp 1698431365
transform 1 0 32032 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_278
timestamp 1698431365
transform 1 0 32480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_290
timestamp 1698431365
transform 1 0 33824 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_292
timestamp 1698431365
transform 1 0 34048 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_310
timestamp 1698431365
transform 1 0 36064 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_314
timestamp 1698431365
transform 1 0 36512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_348
timestamp 1698431365
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_357
timestamp 1698431365
transform 1 0 41328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_365
timestamp 1698431365
transform 1 0 42224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_375
timestamp 1698431365
transform 1 0 43344 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_388
timestamp 1698431365
transform 1 0 44800 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_402
timestamp 1698431365
transform 1 0 46368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_406
timestamp 1698431365
transform 1 0 46816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_33
timestamp 1698431365
transform 1 0 5040 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_45
timestamp 1698431365
transform 1 0 6384 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_70
timestamp 1698431365
transform 1 0 9184 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_103
timestamp 1698431365
transform 1 0 12880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_126
timestamp 1698431365
transform 1 0 15456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_164
timestamp 1698431365
transform 1 0 19712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_166
timestamp 1698431365
transform 1 0 19936 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_193
timestamp 1698431365
transform 1 0 22960 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_234
timestamp 1698431365
transform 1 0 27552 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_238
timestamp 1698431365
transform 1 0 28000 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_242
timestamp 1698431365
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_290
timestamp 1698431365
transform 1 0 33824 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_321
timestamp 1698431365
transform 1 0 37296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_323
timestamp 1698431365
transform 1 0 37520 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_329
timestamp 1698431365
transform 1 0 38192 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_333
timestamp 1698431365
transform 1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_361
timestamp 1698431365
transform 1 0 41776 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_369
timestamp 1698431365
transform 1 0 42672 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_391
timestamp 1698431365
transform 1 0 45136 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_416
timestamp 1698431365
transform 1 0 47936 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_24
timestamp 1698431365
transform 1 0 4032 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_30
timestamp 1698431365
transform 1 0 4704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_34
timestamp 1698431365
transform 1 0 5152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_80
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_89
timestamp 1698431365
transform 1 0 11312 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_93
timestamp 1698431365
transform 1 0 11760 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_100
timestamp 1698431365
transform 1 0 12544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_104
timestamp 1698431365
transform 1 0 12992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_106
timestamp 1698431365
transform 1 0 13216 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_113
timestamp 1698431365
transform 1 0 14000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_117
timestamp 1698431365
transform 1 0 14448 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_121
timestamp 1698431365
transform 1 0 14896 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_144
timestamp 1698431365
transform 1 0 17472 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_151
timestamp 1698431365
transform 1 0 18256 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_165
timestamp 1698431365
transform 1 0 19824 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_175
timestamp 1698431365
transform 1 0 20944 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_179
timestamp 1698431365
transform 1 0 21392 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_198
timestamp 1698431365
transform 1 0 23520 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_202
timestamp 1698431365
transform 1 0 23968 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_228
timestamp 1698431365
transform 1 0 26880 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_232
timestamp 1698431365
transform 1 0 27328 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_234
timestamp 1698431365
transform 1 0 27552 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_264
timestamp 1698431365
transform 1 0 30912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_266
timestamp 1698431365
transform 1 0 31136 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_275
timestamp 1698431365
transform 1 0 32144 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698431365
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_287
timestamp 1698431365
transform 1 0 33488 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_291
timestamp 1698431365
transform 1 0 33936 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_301
timestamp 1698431365
transform 1 0 35056 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_305
timestamp 1698431365
transform 1 0 35504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_312
timestamp 1698431365
transform 1 0 36288 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_316
timestamp 1698431365
transform 1 0 36736 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_332
timestamp 1698431365
transform 1 0 38528 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_340
timestamp 1698431365
transform 1 0 39424 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_357
timestamp 1698431365
transform 1 0 41328 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_361
timestamp 1698431365
transform 1 0 41776 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_369
timestamp 1698431365
transform 1 0 42672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_371
timestamp 1698431365
transform 1 0 42896 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_384
timestamp 1698431365
transform 1 0 44352 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_392
timestamp 1698431365
transform 1 0 45248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_418
timestamp 1698431365
transform 1 0 48160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_51
timestamp 1698431365
transform 1 0 7056 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_53
timestamp 1698431365
transform 1 0 7280 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_91
timestamp 1698431365
transform 1 0 11536 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_99
timestamp 1698431365
transform 1 0 12432 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_103
timestamp 1698431365
transform 1 0 12880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_123
timestamp 1698431365
transform 1 0 15120 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_126
timestamp 1698431365
transform 1 0 15456 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_142
timestamp 1698431365
transform 1 0 17248 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_170
timestamp 1698431365
transform 1 0 20384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698431365
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_183
timestamp 1698431365
transform 1 0 21840 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_187
timestamp 1698431365
transform 1 0 22288 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_195
timestamp 1698431365
transform 1 0 23184 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_252
timestamp 1698431365
transform 1 0 29568 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_256
timestamp 1698431365
transform 1 0 30016 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_260
timestamp 1698431365
transform 1 0 30464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_270
timestamp 1698431365
transform 1 0 31584 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_274
timestamp 1698431365
transform 1 0 32032 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_282
timestamp 1698431365
transform 1 0 32928 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_313
timestamp 1698431365
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_321
timestamp 1698431365
transform 1 0 37296 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_323
timestamp 1698431365
transform 1 0 37520 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_332
timestamp 1698431365
transform 1 0 38528 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_364
timestamp 1698431365
transform 1 0 42112 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_368
timestamp 1698431365
transform 1 0 42560 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_391
timestamp 1698431365
transform 1 0 45136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_6
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_8
timestamp 1698431365
transform 1 0 2240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_11
timestamp 1698431365
transform 1 0 2576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_17
timestamp 1698431365
transform 1 0 3248 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_21
timestamp 1698431365
transform 1 0 3696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_23
timestamp 1698431365
transform 1 0 3920 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_48
timestamp 1698431365
transform 1 0 6720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_50
timestamp 1698431365
transform 1 0 6944 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_82
timestamp 1698431365
transform 1 0 10528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_84
timestamp 1698431365
transform 1 0 10752 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_114
timestamp 1698431365
transform 1 0 14112 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_130
timestamp 1698431365
transform 1 0 15904 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_138
timestamp 1698431365
transform 1 0 16800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_150
timestamp 1698431365
transform 1 0 18144 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_154
timestamp 1698431365
transform 1 0 18592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_158
timestamp 1698431365
transform 1 0 19040 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_166
timestamp 1698431365
transform 1 0 19936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_175
timestamp 1698431365
transform 1 0 20944 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_183
timestamp 1698431365
transform 1 0 21840 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_255
timestamp 1698431365
transform 1 0 29904 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_264
timestamp 1698431365
transform 1 0 30912 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_290
timestamp 1698431365
transform 1 0 33824 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_298
timestamp 1698431365
transform 1 0 34720 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_302
timestamp 1698431365
transform 1 0 35168 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_308
timestamp 1698431365
transform 1 0 35840 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_314
timestamp 1698431365
transform 1 0 36512 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_330
timestamp 1698431365
transform 1 0 38304 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_340
timestamp 1698431365
transform 1 0 39424 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_348
timestamp 1698431365
transform 1 0 40320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_358
timestamp 1698431365
transform 1 0 41440 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_362
timestamp 1698431365
transform 1 0 41888 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_364
timestamp 1698431365
transform 1 0 42112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_384
timestamp 1698431365
transform 1 0 44352 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_400
timestamp 1698431365
transform 1 0 46144 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_6
timestamp 1698431365
transform 1 0 2016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_14
timestamp 1698431365
transform 1 0 2912 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_18
timestamp 1698431365
transform 1 0 3360 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_27
timestamp 1698431365
transform 1 0 4368 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_29
timestamp 1698431365
transform 1 0 4592 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_94
timestamp 1698431365
transform 1 0 11872 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1698431365
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_112
timestamp 1698431365
transform 1 0 13888 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_116
timestamp 1698431365
transform 1 0 14336 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_118
timestamp 1698431365
transform 1 0 14560 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_148
timestamp 1698431365
transform 1 0 17920 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_152
timestamp 1698431365
transform 1 0 18368 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_172
timestamp 1698431365
transform 1 0 20608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_194
timestamp 1698431365
transform 1 0 23072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_251
timestamp 1698431365
transform 1 0 29456 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_267
timestamp 1698431365
transform 1 0 31248 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_269
timestamp 1698431365
transform 1 0 31472 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_284
timestamp 1698431365
transform 1 0 33152 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_292
timestamp 1698431365
transform 1 0 34048 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_303
timestamp 1698431365
transform 1 0 35280 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_312
timestamp 1698431365
transform 1 0 36288 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_319
timestamp 1698431365
transform 1 0 37072 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_334
timestamp 1698431365
transform 1 0 38752 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_368
timestamp 1698431365
transform 1 0 42560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_372
timestamp 1698431365
transform 1 0 43008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_380
timestamp 1698431365
transform 1 0 43904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_419
timestamp 1698431365
transform 1 0 48272 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_46
timestamp 1698431365
transform 1 0 6496 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_50
timestamp 1698431365
transform 1 0 6944 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_54
timestamp 1698431365
transform 1 0 7392 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_57
timestamp 1698431365
transform 1 0 7728 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_61
timestamp 1698431365
transform 1 0 8176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_85
timestamp 1698431365
transform 1 0 10864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_98
timestamp 1698431365
transform 1 0 12320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_102
timestamp 1698431365
transform 1 0 12768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_110
timestamp 1698431365
transform 1 0 13664 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_118
timestamp 1698431365
transform 1 0 14560 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_122
timestamp 1698431365
transform 1 0 15008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_137
timestamp 1698431365
transform 1 0 16688 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698431365
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_162
timestamp 1698431365
transform 1 0 19488 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_170
timestamp 1698431365
transform 1 0 20384 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_176
timestamp 1698431365
transform 1 0 21056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_178
timestamp 1698431365
transform 1 0 21280 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_192
timestamp 1698431365
transform 1 0 22848 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_204
timestamp 1698431365
transform 1 0 24192 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_260
timestamp 1698431365
transform 1 0 30464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_270
timestamp 1698431365
transform 1 0 31584 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698431365
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_286
timestamp 1698431365
transform 1 0 33376 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_292
timestamp 1698431365
transform 1 0 34048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_296
timestamp 1698431365
transform 1 0 34496 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_304
timestamp 1698431365
transform 1 0 35392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_306
timestamp 1698431365
transform 1 0 35616 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_325
timestamp 1698431365
transform 1 0 37744 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_341
timestamp 1698431365
transform 1 0 39536 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_358
timestamp 1698431365
transform 1 0 41440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_365
timestamp 1698431365
transform 1 0 42224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_369
timestamp 1698431365
transform 1 0 42672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_373
timestamp 1698431365
transform 1 0 43120 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_377
timestamp 1698431365
transform 1 0 43568 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_393
timestamp 1698431365
transform 1 0 45360 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_401
timestamp 1698431365
transform 1 0 46256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_403
timestamp 1698431365
transform 1 0 46480 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_406
timestamp 1698431365
transform 1 0 46816 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_414
timestamp 1698431365
transform 1 0 47712 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698431365
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_31
timestamp 1698431365
transform 1 0 4816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_51
timestamp 1698431365
transform 1 0 7056 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_59
timestamp 1698431365
transform 1 0 7952 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_91
timestamp 1698431365
transform 1 0 11536 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_99
timestamp 1698431365
transform 1 0 12432 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_103
timestamp 1698431365
transform 1 0 12880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_115
timestamp 1698431365
transform 1 0 14224 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_119
timestamp 1698431365
transform 1 0 14672 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_128
timestamp 1698431365
transform 1 0 15680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_134
timestamp 1698431365
transform 1 0 16352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_138
timestamp 1698431365
transform 1 0 16800 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_146
timestamp 1698431365
transform 1 0 17696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_150
timestamp 1698431365
transform 1 0 18144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_157
timestamp 1698431365
transform 1 0 18928 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_173
timestamp 1698431365
transform 1 0 20720 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_218
timestamp 1698431365
transform 1 0 25760 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_227
timestamp 1698431365
transform 1 0 26768 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_231
timestamp 1698431365
transform 1 0 27216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_239
timestamp 1698431365
transform 1 0 28112 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_243
timestamp 1698431365
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_276
timestamp 1698431365
transform 1 0 32256 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_289
timestamp 1698431365
transform 1 0 33712 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_293
timestamp 1698431365
transform 1 0 34160 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_309
timestamp 1698431365
transform 1 0 35952 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_313
timestamp 1698431365
transform 1 0 36400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_335
timestamp 1698431365
transform 1 0 38864 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_351
timestamp 1698431365
transform 1 0 40656 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_353
timestamp 1698431365
transform 1 0 40880 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_366
timestamp 1698431365
transform 1 0 42336 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_391
timestamp 1698431365
transform 1 0 45136 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_8
timestamp 1698431365
transform 1 0 2240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_12
timestamp 1698431365
transform 1 0 2688 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_28
timestamp 1698431365
transform 1 0 4480 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_36
timestamp 1698431365
transform 1 0 5376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_58
timestamp 1698431365
transform 1 0 7840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_62
timestamp 1698431365
transform 1 0 8288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_82
timestamp 1698431365
transform 1 0 10528 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_90
timestamp 1698431365
transform 1 0 11424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_100
timestamp 1698431365
transform 1 0 12544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_151
timestamp 1698431365
transform 1 0 18256 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_198
timestamp 1698431365
transform 1 0 23520 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_200
timestamp 1698431365
transform 1 0 23744 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_207
timestamp 1698431365
transform 1 0 24528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698431365
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_237
timestamp 1698431365
transform 1 0 27888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_270
timestamp 1698431365
transform 1 0 31584 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_274
timestamp 1698431365
transform 1 0 32032 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_278
timestamp 1698431365
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_284
timestamp 1698431365
transform 1 0 33152 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_298
timestamp 1698431365
transform 1 0 34720 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_314
timestamp 1698431365
transform 1 0 36512 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_322
timestamp 1698431365
transform 1 0 37408 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_357
timestamp 1698431365
transform 1 0 41328 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_361
timestamp 1698431365
transform 1 0 41776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_363
timestamp 1698431365
transform 1 0 42000 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_384
timestamp 1698431365
transform 1 0 44352 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_410
timestamp 1698431365
transform 1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_418
timestamp 1698431365
transform 1 0 48160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_63
timestamp 1698431365
transform 1 0 8400 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_71
timestamp 1698431365
transform 1 0 9296 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_75
timestamp 1698431365
transform 1 0 9744 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_112
timestamp 1698431365
transform 1 0 13888 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_133
timestamp 1698431365
transform 1 0 16240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_236
timestamp 1698431365
transform 1 0 27776 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_240
timestamp 1698431365
transform 1 0 28224 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_279
timestamp 1698431365
transform 1 0 32592 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_283
timestamp 1698431365
transform 1 0 33040 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_300
timestamp 1698431365
transform 1 0 34944 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_304
timestamp 1698431365
transform 1 0 35392 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_310
timestamp 1698431365
transform 1 0 36064 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_341
timestamp 1698431365
transform 1 0 39536 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_357
timestamp 1698431365
transform 1 0 41328 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_373
timestamp 1698431365
transform 1 0 43120 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_377
timestamp 1698431365
transform 1 0 43568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_391
timestamp 1698431365
transform 1 0 45136 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_393
timestamp 1698431365
transform 1 0 45360 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_410
timestamp 1698431365
transform 1 0 47264 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_418
timestamp 1698431365
transform 1 0 48160 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_8
timestamp 1698431365
transform 1 0 2240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_12
timestamp 1698431365
transform 1 0 2688 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_28
timestamp 1698431365
transform 1 0 4480 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_32
timestamp 1698431365
transform 1 0 4928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_35
timestamp 1698431365
transform 1 0 5264 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_53
timestamp 1698431365
transform 1 0 7280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_55
timestamp 1698431365
transform 1 0 7504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_76
timestamp 1698431365
transform 1 0 9856 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_86
timestamp 1698431365
transform 1 0 10976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_88
timestamp 1698431365
transform 1 0 11200 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_94
timestamp 1698431365
transform 1 0 11872 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_98
timestamp 1698431365
transform 1 0 12320 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_106
timestamp 1698431365
transform 1 0 13216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_115
timestamp 1698431365
transform 1 0 14224 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_131
timestamp 1698431365
transform 1 0 16016 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_135
timestamp 1698431365
transform 1 0 16464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_137
timestamp 1698431365
transform 1 0 16688 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_147
timestamp 1698431365
transform 1 0 17808 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_151
timestamp 1698431365
transform 1 0 18256 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_217
timestamp 1698431365
transform 1 0 25648 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_255
timestamp 1698431365
transform 1 0 29904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_259
timestamp 1698431365
transform 1 0 30352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_263
timestamp 1698431365
transform 1 0 30800 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_279
timestamp 1698431365
transform 1 0 32592 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_322
timestamp 1698431365
transform 1 0 37408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_335
timestamp 1698431365
transform 1 0 38864 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_343
timestamp 1698431365
transform 1 0 39760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_347
timestamp 1698431365
transform 1 0 40208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_349
timestamp 1698431365
transform 1 0 40432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_357
timestamp 1698431365
transform 1 0 41328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_361
timestamp 1698431365
transform 1 0 41776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_365
timestamp 1698431365
transform 1 0 42224 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_397
timestamp 1698431365
transform 1 0 45808 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_401
timestamp 1698431365
transform 1 0 46256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_403
timestamp 1698431365
transform 1 0 46480 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_33
timestamp 1698431365
transform 1 0 5040 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_50
timestamp 1698431365
transform 1 0 6944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_52
timestamp 1698431365
transform 1 0 7168 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_66
timestamp 1698431365
transform 1 0 8736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_78
timestamp 1698431365
transform 1 0 10080 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_82
timestamp 1698431365
transform 1 0 10528 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_86
timestamp 1698431365
transform 1 0 10976 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_102
timestamp 1698431365
transform 1 0 12768 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_104
timestamp 1698431365
transform 1 0 12992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_112
timestamp 1698431365
transform 1 0 13888 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_120
timestamp 1698431365
transform 1 0 14784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_122
timestamp 1698431365
transform 1 0 15008 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_125
timestamp 1698431365
transform 1 0 15344 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_131
timestamp 1698431365
transform 1 0 16016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_193
timestamp 1698431365
transform 1 0 22960 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_242
timestamp 1698431365
transform 1 0 28448 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_244
timestamp 1698431365
transform 1 0 28672 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_251
timestamp 1698431365
transform 1 0 29456 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_265
timestamp 1698431365
transform 1 0 31024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_269
timestamp 1698431365
transform 1 0 31472 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_273
timestamp 1698431365
transform 1 0 31920 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_277
timestamp 1698431365
transform 1 0 32368 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_279
timestamp 1698431365
transform 1 0 32592 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_288
timestamp 1698431365
transform 1 0 33600 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_296
timestamp 1698431365
transform 1 0 34496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_300
timestamp 1698431365
transform 1 0 34944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_302
timestamp 1698431365
transform 1 0 35168 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_322
timestamp 1698431365
transform 1 0 37408 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_330
timestamp 1698431365
transform 1 0 38304 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_334
timestamp 1698431365
transform 1 0 38752 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_337
timestamp 1698431365
transform 1 0 39088 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_341
timestamp 1698431365
transform 1 0 39536 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_367
timestamp 1698431365
transform 1 0 42448 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_381
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_392
timestamp 1698431365
transform 1 0 45248 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_408
timestamp 1698431365
transform 1 0 47040 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_416
timestamp 1698431365
transform 1 0 47936 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_10
timestamp 1698431365
transform 1 0 2464 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_14
timestamp 1698431365
transform 1 0 2912 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_21
timestamp 1698431365
transform 1 0 3696 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_53
timestamp 1698431365
transform 1 0 7280 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_69
timestamp 1698431365
transform 1 0 9072 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_80
timestamp 1698431365
transform 1 0 10304 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_113
timestamp 1698431365
transform 1 0 14000 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_122
timestamp 1698431365
transform 1 0 15008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_124
timestamp 1698431365
transform 1 0 15232 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_131
timestamp 1698431365
transform 1 0 16016 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_159
timestamp 1698431365
transform 1 0 19152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_163
timestamp 1698431365
transform 1 0 19600 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_269
timestamp 1698431365
transform 1 0 31472 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_277
timestamp 1698431365
transform 1 0 32368 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_279
timestamp 1698431365
transform 1 0 32592 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_286
timestamp 1698431365
transform 1 0 33376 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_294
timestamp 1698431365
transform 1 0 34272 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_326
timestamp 1698431365
transform 1 0 37856 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_328
timestamp 1698431365
transform 1 0 38080 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_340
timestamp 1698431365
transform 1 0 39424 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_344
timestamp 1698431365
transform 1 0 39872 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_348
timestamp 1698431365
transform 1 0 40320 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_360
timestamp 1698431365
transform 1 0 41664 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_364
timestamp 1698431365
transform 1 0 42112 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_378
timestamp 1698431365
transform 1 0 43680 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_380
timestamp 1698431365
transform 1 0 43904 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_403
timestamp 1698431365
transform 1 0 46480 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_407
timestamp 1698431365
transform 1 0 46928 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_415
timestamp 1698431365
transform 1 0 47824 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_419
timestamp 1698431365
transform 1 0 48272 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_8
timestamp 1698431365
transform 1 0 2240 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_12
timestamp 1698431365
transform 1 0 2688 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_28
timestamp 1698431365
transform 1 0 4480 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_32
timestamp 1698431365
transform 1 0 4928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_51
timestamp 1698431365
transform 1 0 7056 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_59
timestamp 1698431365
transform 1 0 7952 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_80
timestamp 1698431365
transform 1 0 10304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_84
timestamp 1698431365
transform 1 0 10752 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_88
timestamp 1698431365
transform 1 0 11200 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_92
timestamp 1698431365
transform 1 0 11648 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_100
timestamp 1698431365
transform 1 0 12544 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_104
timestamp 1698431365
transform 1 0 12992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_136
timestamp 1698431365
transform 1 0 16576 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_144
timestamp 1698431365
transform 1 0 17472 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_147
timestamp 1698431365
transform 1 0 17808 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_151
timestamp 1698431365
transform 1 0 18256 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_161
timestamp 1698431365
transform 1 0 19376 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_169
timestamp 1698431365
transform 1 0 20272 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_173
timestamp 1698431365
transform 1 0 20720 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_185
timestamp 1698431365
transform 1 0 22064 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_188
timestamp 1698431365
transform 1 0 22400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_192
timestamp 1698431365
transform 1 0 22848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_196
timestamp 1698431365
transform 1 0 23296 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_213
timestamp 1698431365
transform 1 0 25200 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_215
timestamp 1698431365
transform 1 0 25424 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_231
timestamp 1698431365
transform 1 0 27216 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_239
timestamp 1698431365
transform 1 0 28112 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_277
timestamp 1698431365
transform 1 0 32368 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_309
timestamp 1698431365
transform 1 0 35952 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_313
timestamp 1698431365
transform 1 0 36400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_325
timestamp 1698431365
transform 1 0 37744 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_328
timestamp 1698431365
transform 1 0 38080 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_332
timestamp 1698431365
transform 1 0 38528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_340
timestamp 1698431365
transform 1 0 39424 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_342
timestamp 1698431365
transform 1 0 39648 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_348
timestamp 1698431365
transform 1 0 40320 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_352
timestamp 1698431365
transform 1 0 40768 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_356
timestamp 1698431365
transform 1 0 41216 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_364
timestamp 1698431365
transform 1 0 42112 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_366
timestamp 1698431365
transform 1 0 42336 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_384
timestamp 1698431365
transform 1 0 44352 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_399
timestamp 1698431365
transform 1 0 46032 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_34
timestamp 1698431365
transform 1 0 5152 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_38
timestamp 1698431365
transform 1 0 5600 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_40
timestamp 1698431365
transform 1 0 5824 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_43
timestamp 1698431365
transform 1 0 6160 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_47
timestamp 1698431365
transform 1 0 6608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_51
timestamp 1698431365
transform 1 0 7056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_55
timestamp 1698431365
transform 1 0 7504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_65
timestamp 1698431365
transform 1 0 8624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_67
timestamp 1698431365
transform 1 0 8848 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_80
timestamp 1698431365
transform 1 0 10304 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_84
timestamp 1698431365
transform 1 0 10752 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_116
timestamp 1698431365
transform 1 0 14336 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_132
timestamp 1698431365
transform 1 0 16128 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_144
timestamp 1698431365
transform 1 0 17472 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_187
timestamp 1698431365
transform 1 0 22288 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_191
timestamp 1698431365
transform 1 0 22736 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_193
timestamp 1698431365
transform 1 0 22960 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_196
timestamp 1698431365
transform 1 0 23296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_205
timestamp 1698431365
transform 1 0 24304 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_209
timestamp 1698431365
transform 1 0 24752 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_219
timestamp 1698431365
transform 1 0 25872 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_223
timestamp 1698431365
transform 1 0 26320 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_227
timestamp 1698431365
transform 1 0 26768 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_257
timestamp 1698431365
transform 1 0 30128 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_269
timestamp 1698431365
transform 1 0 31472 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_277
timestamp 1698431365
transform 1 0 32368 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_279
timestamp 1698431365
transform 1 0 32592 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_290
timestamp 1698431365
transform 1 0 33824 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_294
timestamp 1698431365
transform 1 0 34272 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_302
timestamp 1698431365
transform 1 0 35168 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_304
timestamp 1698431365
transform 1 0 35392 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_330
timestamp 1698431365
transform 1 0 38304 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_334
timestamp 1698431365
transform 1 0 38752 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_338
timestamp 1698431365
transform 1 0 39200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_342
timestamp 1698431365
transform 1 0 39648 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_346
timestamp 1698431365
transform 1 0 40096 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_384
timestamp 1698431365
transform 1 0 44352 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_392
timestamp 1698431365
transform 1 0 45248 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_408
timestamp 1698431365
transform 1 0 47040 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_6
timestamp 1698431365
transform 1 0 2016 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_22
timestamp 1698431365
transform 1 0 3808 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_30
timestamp 1698431365
transform 1 0 4704 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_41
timestamp 1698431365
transform 1 0 5936 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_86
timestamp 1698431365
transform 1 0 10976 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_102
timestamp 1698431365
transform 1 0 12768 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_104
timestamp 1698431365
transform 1 0 12992 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_123
timestamp 1698431365
transform 1 0 15120 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_131
timestamp 1698431365
transform 1 0 16016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_135
timestamp 1698431365
transform 1 0 16464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_143
timestamp 1698431365
transform 1 0 17360 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_147
timestamp 1698431365
transform 1 0 17808 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_153
timestamp 1698431365
transform 1 0 18480 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_161
timestamp 1698431365
transform 1 0 19376 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_173
timestamp 1698431365
transform 1 0 20720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_194
timestamp 1698431365
transform 1 0 23072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_198
timestamp 1698431365
transform 1 0 23520 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_206
timestamp 1698431365
transform 1 0 24416 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_263
timestamp 1698431365
transform 1 0 30800 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_265
timestamp 1698431365
transform 1 0 31024 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_295
timestamp 1698431365
transform 1 0 34384 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_297
timestamp 1698431365
transform 1 0 34608 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_304
timestamp 1698431365
transform 1 0 35392 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_314
timestamp 1698431365
transform 1 0 36512 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_337
timestamp 1698431365
transform 1 0 39088 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_339
timestamp 1698431365
transform 1 0 39312 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_356
timestamp 1698431365
transform 1 0 41216 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_372
timestamp 1698431365
transform 1 0 43008 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_380
timestamp 1698431365
transform 1 0 43904 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_384
timestamp 1698431365
transform 1 0 44352 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_419
timestamp 1698431365
transform 1 0 48272 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_10
timestamp 1698431365
transform 1 0 2464 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_18
timestamp 1698431365
transform 1 0 3360 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_22
timestamp 1698431365
transform 1 0 3808 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_29
timestamp 1698431365
transform 1 0 4592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_33
timestamp 1698431365
transform 1 0 5040 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_60
timestamp 1698431365
transform 1 0 8064 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_67
timestamp 1698431365
transform 1 0 8848 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_69
timestamp 1698431365
transform 1 0 9072 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_76
timestamp 1698431365
transform 1 0 9856 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_84
timestamp 1698431365
transform 1 0 10752 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_86
timestamp 1698431365
transform 1 0 10976 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_116
timestamp 1698431365
transform 1 0 14336 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_122
timestamp 1698431365
transform 1 0 15008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_144
timestamp 1698431365
transform 1 0 17472 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_209
timestamp 1698431365
transform 1 0 24752 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_218
timestamp 1698431365
transform 1 0 25760 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_234
timestamp 1698431365
transform 1 0 27552 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_242
timestamp 1698431365
transform 1 0 28448 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_256
timestamp 1698431365
transform 1 0 30016 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_264
timestamp 1698431365
transform 1 0 30912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_293
timestamp 1698431365
transform 1 0 34160 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_324
timestamp 1698431365
transform 1 0 37632 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_326
timestamp 1698431365
transform 1 0 37856 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_366
timestamp 1698431365
transform 1 0 42336 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_398
timestamp 1698431365
transform 1 0 45920 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_414
timestamp 1698431365
transform 1 0 47712 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_418
timestamp 1698431365
transform 1 0 48160 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_51
timestamp 1698431365
transform 1 0 7056 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_81
timestamp 1698431365
transform 1 0 10416 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_98
timestamp 1698431365
transform 1 0 12320 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_121
timestamp 1698431365
transform 1 0 14896 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_123
timestamp 1698431365
transform 1 0 15120 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_173
timestamp 1698431365
transform 1 0 20720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_194
timestamp 1698431365
transform 1 0 23072 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_212
timestamp 1698431365
transform 1 0 25088 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_228
timestamp 1698431365
transform 1 0 26880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_238
timestamp 1698431365
transform 1 0 28000 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_242
timestamp 1698431365
transform 1 0 28448 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_244
timestamp 1698431365
transform 1 0 28672 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_260
timestamp 1698431365
transform 1 0 30464 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_268
timestamp 1698431365
transform 1 0 31360 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_275
timestamp 1698431365
transform 1 0 32144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_277
timestamp 1698431365
transform 1 0 32368 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_291
timestamp 1698431365
transform 1 0 33936 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_295
timestamp 1698431365
transform 1 0 34384 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_338
timestamp 1698431365
transform 1 0 39200 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_375
timestamp 1698431365
transform 1 0 43344 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_383
timestamp 1698431365
transform 1 0 44240 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_391
timestamp 1698431365
transform 1 0 45136 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_407
timestamp 1698431365
transform 1 0 46928 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_415
timestamp 1698431365
transform 1 0 47824 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_18
timestamp 1698431365
transform 1 0 3360 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_26
timestamp 1698431365
transform 1 0 4256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_28
timestamp 1698431365
transform 1 0 4480 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_51
timestamp 1698431365
transform 1 0 7056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_55
timestamp 1698431365
transform 1 0 7504 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_59
timestamp 1698431365
transform 1 0 7952 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_61
timestamp 1698431365
transform 1 0 8176 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_76
timestamp 1698431365
transform 1 0 9856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_78
timestamp 1698431365
transform 1 0 10080 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_85
timestamp 1698431365
transform 1 0 10864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_89
timestamp 1698431365
transform 1 0 11312 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_107
timestamp 1698431365
transform 1 0 13328 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_111
timestamp 1698431365
transform 1 0 13776 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_113
timestamp 1698431365
transform 1 0 14000 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_116
timestamp 1698431365
transform 1 0 14336 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_138
timestamp 1698431365
transform 1 0 16800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_147
timestamp 1698431365
transform 1 0 17808 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_153
timestamp 1698431365
transform 1 0 18480 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_155
timestamp 1698431365
transform 1 0 18704 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_158
timestamp 1698431365
transform 1 0 19040 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_160
timestamp 1698431365
transform 1 0 19264 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_163
timestamp 1698431365
transform 1 0 19600 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_179
timestamp 1698431365
transform 1 0 21392 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_220
timestamp 1698431365
transform 1 0 25984 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_224
timestamp 1698431365
transform 1 0 26432 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_236
timestamp 1698431365
transform 1 0 27776 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_240
timestamp 1698431365
transform 1 0 28224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_242
timestamp 1698431365
transform 1 0 28448 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_270
timestamp 1698431365
transform 1 0 31584 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_274
timestamp 1698431365
transform 1 0 32032 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_277
timestamp 1698431365
transform 1 0 32368 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_279
timestamp 1698431365
transform 1 0 32592 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_286
timestamp 1698431365
transform 1 0 33376 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_302
timestamp 1698431365
transform 1 0 35168 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_310
timestamp 1698431365
transform 1 0 36064 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_320
timestamp 1698431365
transform 1 0 37184 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_336
timestamp 1698431365
transform 1 0 38976 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_344
timestamp 1698431365
transform 1 0 39872 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_348
timestamp 1698431365
transform 1 0 40320 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_356
timestamp 1698431365
transform 1 0 41216 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_394
timestamp 1698431365
transform 1 0 45472 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_403
timestamp 1698431365
transform 1 0 46480 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_419
timestamp 1698431365
transform 1 0 48272 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_6
timestamp 1698431365
transform 1 0 2016 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_22
timestamp 1698431365
transform 1 0 3808 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_30
timestamp 1698431365
transform 1 0 4704 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_41
timestamp 1698431365
transform 1 0 5936 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_45
timestamp 1698431365
transform 1 0 6384 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_49
timestamp 1698431365
transform 1 0 6832 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_81
timestamp 1698431365
transform 1 0 10416 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_97
timestamp 1698431365
transform 1 0 12208 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_111
timestamp 1698431365
transform 1 0 13776 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_120
timestamp 1698431365
transform 1 0 14784 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_128
timestamp 1698431365
transform 1 0 15680 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_132
timestamp 1698431365
transform 1 0 16128 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_135
timestamp 1698431365
transform 1 0 16464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_139
timestamp 1698431365
transform 1 0 16912 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_161
timestamp 1698431365
transform 1 0 19376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_209
timestamp 1698431365
transform 1 0 24752 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_213
timestamp 1698431365
transform 1 0 25200 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_236
timestamp 1698431365
transform 1 0 27776 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_240
timestamp 1698431365
transform 1 0 28224 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_244
timestamp 1698431365
transform 1 0 28672 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_278
timestamp 1698431365
transform 1 0 32480 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_286
timestamp 1698431365
transform 1 0 33376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_309
timestamp 1698431365
transform 1 0 35952 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_313
timestamp 1698431365
transform 1 0 36400 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_349
timestamp 1698431365
transform 1 0 40432 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_391
timestamp 1698431365
transform 1 0 45136 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_408
timestamp 1698431365
transform 1 0 47040 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_416
timestamp 1698431365
transform 1 0 47936 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_10
timestamp 1698431365
transform 1 0 2464 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_42
timestamp 1698431365
transform 1 0 6048 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_58
timestamp 1698431365
transform 1 0 7840 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_66
timestamp 1698431365
transform 1 0 8736 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_74
timestamp 1698431365
transform 1 0 9632 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_77
timestamp 1698431365
transform 1 0 9968 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_79
timestamp 1698431365
transform 1 0 10192 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_82
timestamp 1698431365
transform 1 0 10528 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_96
timestamp 1698431365
transform 1 0 12096 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_102
timestamp 1698431365
transform 1 0 12768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_106
timestamp 1698431365
transform 1 0 13216 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_116
timestamp 1698431365
transform 1 0 14336 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_120
timestamp 1698431365
transform 1 0 14784 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_193
timestamp 1698431365
transform 1 0 22960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_197
timestamp 1698431365
transform 1 0 23408 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_205
timestamp 1698431365
transform 1 0 24304 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_209
timestamp 1698431365
transform 1 0 24752 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_233
timestamp 1698431365
transform 1 0 27440 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_237
timestamp 1698431365
transform 1 0 27888 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_247
timestamp 1698431365
transform 1 0 29008 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_254
timestamp 1698431365
transform 1 0 29792 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_265
timestamp 1698431365
transform 1 0 31024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_267
timestamp 1698431365
transform 1 0 31248 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_270
timestamp 1698431365
transform 1 0 31584 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_274
timestamp 1698431365
transform 1 0 32032 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_278
timestamp 1698431365
transform 1 0 32480 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_298
timestamp 1698431365
transform 1 0 34720 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_318
timestamp 1698431365
transform 1 0 36960 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_322
timestamp 1698431365
transform 1 0 37408 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_324
timestamp 1698431365
transform 1 0 37632 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_347
timestamp 1698431365
transform 1 0 40208 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_349
timestamp 1698431365
transform 1 0 40432 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_368
timestamp 1698431365
transform 1 0 42560 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_370
timestamp 1698431365
transform 1 0 42784 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_375
timestamp 1698431365
transform 1 0 43344 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_379
timestamp 1698431365
transform 1 0 43792 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_405
timestamp 1698431365
transform 1 0 46704 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_413
timestamp 1698431365
transform 1 0 47600 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_415
timestamp 1698431365
transform 1 0 47824 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_50
timestamp 1698431365
transform 1 0 6944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_54
timestamp 1698431365
transform 1 0 7392 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_58
timestamp 1698431365
transform 1 0 7840 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_81
timestamp 1698431365
transform 1 0 10416 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_123
timestamp 1698431365
transform 1 0 15120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_125
timestamp 1698431365
transform 1 0 15344 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_128
timestamp 1698431365
transform 1 0 15680 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_132
timestamp 1698431365
transform 1 0 16128 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_136
timestamp 1698431365
transform 1 0 16576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_154
timestamp 1698431365
transform 1 0 18592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_172
timestamp 1698431365
transform 1 0 20608 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_174
timestamp 1698431365
transform 1 0 20832 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_187
timestamp 1698431365
transform 1 0 22288 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_203
timestamp 1698431365
transform 1 0 24080 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_211
timestamp 1698431365
transform 1 0 24976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_225
timestamp 1698431365
transform 1 0 26544 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_251
timestamp 1698431365
transform 1 0 29456 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_253
timestamp 1698431365
transform 1 0 29680 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_256
timestamp 1698431365
transform 1 0 30016 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_260
timestamp 1698431365
transform 1 0 30464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_264
timestamp 1698431365
transform 1 0 30912 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_267
timestamp 1698431365
transform 1 0 31248 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_283
timestamp 1698431365
transform 1 0 33040 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_287
timestamp 1698431365
transform 1 0 33488 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_309
timestamp 1698431365
transform 1 0 35952 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_313
timestamp 1698431365
transform 1 0 36400 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_321
timestamp 1698431365
transform 1 0 37296 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_337
timestamp 1698431365
transform 1 0 39088 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_361
timestamp 1698431365
transform 1 0 41776 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_377
timestamp 1698431365
transform 1 0 43568 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_419
timestamp 1698431365
transform 1 0 48272 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_6
timestamp 1698431365
transform 1 0 2016 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_22
timestamp 1698431365
transform 1 0 3808 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_24
timestamp 1698431365
transform 1 0 4032 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_59
timestamp 1698431365
transform 1 0 7952 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_63
timestamp 1698431365
transform 1 0 8400 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_67
timestamp 1698431365
transform 1 0 8848 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_69
timestamp 1698431365
transform 1 0 9072 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_76
timestamp 1698431365
transform 1 0 9856 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_79
timestamp 1698431365
transform 1 0 10192 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_83
timestamp 1698431365
transform 1 0 10640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_103
timestamp 1698431365
transform 1 0 12880 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_105
timestamp 1698431365
transform 1 0 13104 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_138
timestamp 1698431365
transform 1 0 16800 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_150
timestamp 1698431365
transform 1 0 18144 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_152
timestamp 1698431365
transform 1 0 18368 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_159
timestamp 1698431365
transform 1 0 19152 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_163
timestamp 1698431365
transform 1 0 19600 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_166
timestamp 1698431365
transform 1 0 19936 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_244
timestamp 1698431365
transform 1 0 28672 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_252
timestamp 1698431365
transform 1 0 29568 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_254
timestamp 1698431365
transform 1 0 29792 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_265
timestamp 1698431365
transform 1 0 31024 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_273
timestamp 1698431365
transform 1 0 31920 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_294
timestamp 1698431365
transform 1 0 34272 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_302
timestamp 1698431365
transform 1 0 35168 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_306
timestamp 1698431365
transform 1 0 35616 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_344
timestamp 1698431365
transform 1 0 39872 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_358
timestamp 1698431365
transform 1 0 41440 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_360
timestamp 1698431365
transform 1 0 41664 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_373
timestamp 1698431365
transform 1 0 43120 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_405
timestamp 1698431365
transform 1 0 46704 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_413
timestamp 1698431365
transform 1 0 47600 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_417
timestamp 1698431365
transform 1 0 48048 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_419
timestamp 1698431365
transform 1 0 48272 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_10
timestamp 1698431365
transform 1 0 2464 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_26
timestamp 1698431365
transform 1 0 4256 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_43
timestamp 1698431365
transform 1 0 6160 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_74
timestamp 1698431365
transform 1 0 9632 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_90
timestamp 1698431365
transform 1 0 11424 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_92
timestamp 1698431365
transform 1 0 11648 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_100
timestamp 1698431365
transform 1 0 12544 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_102
timestamp 1698431365
transform 1 0 12768 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_109
timestamp 1698431365
transform 1 0 13552 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_130
timestamp 1698431365
transform 1 0 15904 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_160
timestamp 1698431365
transform 1 0 19264 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_168
timestamp 1698431365
transform 1 0 20160 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_172
timestamp 1698431365
transform 1 0 20608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_174
timestamp 1698431365
transform 1 0 20832 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_179
timestamp 1698431365
transform 1 0 21392 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_209
timestamp 1698431365
transform 1 0 24752 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_217
timestamp 1698431365
transform 1 0 25648 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_221
timestamp 1698431365
transform 1 0 26096 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_223
timestamp 1698431365
transform 1 0 26320 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_234
timestamp 1698431365
transform 1 0 27552 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_238
timestamp 1698431365
transform 1 0 28000 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_242
timestamp 1698431365
transform 1 0 28448 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_244
timestamp 1698431365
transform 1 0 28672 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_259
timestamp 1698431365
transform 1 0 30352 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_263
timestamp 1698431365
transform 1 0 30800 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_267
timestamp 1698431365
transform 1 0 31248 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_301
timestamp 1698431365
transform 1 0 35056 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_317
timestamp 1698431365
transform 1 0 36848 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_344
timestamp 1698431365
transform 1 0 39872 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_348
timestamp 1698431365
transform 1 0 40320 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_360
timestamp 1698431365
transform 1 0 41664 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_369
timestamp 1698431365
transform 1 0 42672 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_403
timestamp 1698431365
transform 1 0 46480 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_411
timestamp 1698431365
transform 1 0 47376 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_415
timestamp 1698431365
transform 1 0 47824 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_34
timestamp 1698431365
transform 1 0 5152 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_42
timestamp 1698431365
transform 1 0 6048 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_46
timestamp 1698431365
transform 1 0 6496 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_53
timestamp 1698431365
transform 1 0 7280 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_69
timestamp 1698431365
transform 1 0 9072 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_103
timestamp 1698431365
transform 1 0 12880 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_111
timestamp 1698431365
transform 1 0 13776 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_124
timestamp 1698431365
transform 1 0 15232 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_128
timestamp 1698431365
transform 1 0 15680 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_132
timestamp 1698431365
transform 1 0 16128 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_156
timestamp 1698431365
transform 1 0 18816 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_164
timestamp 1698431365
transform 1 0 19712 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_168
timestamp 1698431365
transform 1 0 20160 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_176
timestamp 1698431365
transform 1 0 21056 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_198
timestamp 1698431365
transform 1 0 23520 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_206
timestamp 1698431365
transform 1 0 24416 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_214
timestamp 1698431365
transform 1 0 25312 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_230
timestamp 1698431365
transform 1 0 27104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_269
timestamp 1698431365
transform 1 0 31472 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_273
timestamp 1698431365
transform 1 0 31920 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_277
timestamp 1698431365
transform 1 0 32368 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_279
timestamp 1698431365
transform 1 0 32592 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_287
timestamp 1698431365
transform 1 0 33488 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_315
timestamp 1698431365
transform 1 0 36624 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_331
timestamp 1698431365
transform 1 0 38416 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_333
timestamp 1698431365
transform 1 0 38640 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_342
timestamp 1698431365
transform 1 0 39648 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_366
timestamp 1698431365
transform 1 0 42336 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_388
timestamp 1698431365
transform 1 0 44800 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_2
timestamp 1698431365
transform 1 0 1568 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_6
timestamp 1698431365
transform 1 0 2016 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_22
timestamp 1698431365
transform 1 0 3808 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_30
timestamp 1698431365
transform 1 0 4704 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_45
timestamp 1698431365
transform 1 0 6384 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_49
timestamp 1698431365
transform 1 0 6832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_51
timestamp 1698431365
transform 1 0 7056 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_59
timestamp 1698431365
transform 1 0 7952 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_63
timestamp 1698431365
transform 1 0 8400 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_71
timestamp 1698431365
transform 1 0 9296 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_75
timestamp 1698431365
transform 1 0 9744 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_82
timestamp 1698431365
transform 1 0 10528 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_98
timestamp 1698431365
transform 1 0 12320 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_102
timestamp 1698431365
transform 1 0 12768 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_104
timestamp 1698431365
transform 1 0 12992 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_123
timestamp 1698431365
transform 1 0 15120 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_126
timestamp 1698431365
transform 1 0 15456 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_134
timestamp 1698431365
transform 1 0 16352 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_138
timestamp 1698431365
transform 1 0 16800 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_193
timestamp 1698431365
transform 1 0 22960 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_201
timestamp 1698431365
transform 1 0 23856 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_205
timestamp 1698431365
transform 1 0 24304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_207
timestamp 1698431365
transform 1 0 24528 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_210
timestamp 1698431365
transform 1 0 24864 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_218
timestamp 1698431365
transform 1 0 25760 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_220
timestamp 1698431365
transform 1 0 25984 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_234
timestamp 1698431365
transform 1 0 27552 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_238
timestamp 1698431365
transform 1 0 28000 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_242
timestamp 1698431365
transform 1 0 28448 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_244
timestamp 1698431365
transform 1 0 28672 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_259
timestamp 1698431365
transform 1 0 30352 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_263
timestamp 1698431365
transform 1 0 30800 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_267
timestamp 1698431365
transform 1 0 31248 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_309
timestamp 1698431365
transform 1 0 35952 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_313
timestamp 1698431365
transform 1 0 36400 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_333
timestamp 1698431365
transform 1 0 38640 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_337
timestamp 1698431365
transform 1 0 39088 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_358
timestamp 1698431365
transform 1 0 41440 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_366
timestamp 1698431365
transform 1 0 42336 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_370
timestamp 1698431365
transform 1 0 42784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_372
timestamp 1698431365
transform 1 0 43008 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_381
timestamp 1698431365
transform 1 0 44016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_387
timestamp 1698431365
transform 1 0 44688 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_419
timestamp 1698431365
transform 1 0 48272 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_10
timestamp 1698431365
transform 1 0 2464 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_26
timestamp 1698431365
transform 1 0 4256 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_34
timestamp 1698431365
transform 1 0 5152 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_38
timestamp 1698431365
transform 1 0 5600 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_69
timestamp 1698431365
transform 1 0 9072 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_80
timestamp 1698431365
transform 1 0 10304 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_112
timestamp 1698431365
transform 1 0 13888 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_128
timestamp 1698431365
transform 1 0 15680 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_174
timestamp 1698431365
transform 1 0 20832 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_190
timestamp 1698431365
transform 1 0 22624 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_194
timestamp 1698431365
transform 1 0 23072 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_208
timestamp 1698431365
transform 1 0 24640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_226
timestamp 1698431365
transform 1 0 26656 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_232
timestamp 1698431365
transform 1 0 27328 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_238
timestamp 1698431365
transform 1 0 28000 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_270
timestamp 1698431365
transform 1 0 31584 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_278
timestamp 1698431365
transform 1 0 32480 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_286
timestamp 1698431365
transform 1 0 33376 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_304
timestamp 1698431365
transform 1 0 35392 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_308
timestamp 1698431365
transform 1 0 35840 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_324
timestamp 1698431365
transform 1 0 37632 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_348
timestamp 1698431365
transform 1 0 40320 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_352
timestamp 1698431365
transform 1 0 40768 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_104
timestamp 1698431365
transform 1 0 12992 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_111
timestamp 1698431365
transform 1 0 13776 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_148
timestamp 1698431365
transform 1 0 17920 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_152
timestamp 1698431365
transform 1 0 18368 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_156
timestamp 1698431365
transform 1 0 18816 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_172
timestamp 1698431365
transform 1 0 20608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_174
timestamp 1698431365
transform 1 0 20832 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_185
timestamp 1698431365
transform 1 0 22064 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_200
timestamp 1698431365
transform 1 0 23744 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_206
timestamp 1698431365
transform 1 0 24416 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_222
timestamp 1698431365
transform 1 0 26208 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_240
timestamp 1698431365
transform 1 0 28224 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_244
timestamp 1698431365
transform 1 0 28672 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_255
timestamp 1698431365
transform 1 0 29904 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_271
timestamp 1698431365
transform 1 0 31696 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_279
timestamp 1698431365
transform 1 0 32592 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_281
timestamp 1698431365
transform 1 0 32816 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_288
timestamp 1698431365
transform 1 0 33600 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_296
timestamp 1698431365
transform 1 0 34496 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_300
timestamp 1698431365
transform 1 0 34944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_304
timestamp 1698431365
transform 1 0 35392 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_308
timestamp 1698431365
transform 1 0 35840 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_310
timestamp 1698431365
transform 1 0 36064 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_342
timestamp 1698431365
transform 1 0 39648 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_358
timestamp 1698431365
transform 1 0 41440 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_372
timestamp 1698431365
transform 1 0 43008 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_380
timestamp 1698431365
transform 1 0 43904 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_384
timestamp 1698431365
transform 1 0 44352 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_419
timestamp 1698431365
transform 1 0 48272 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_6
timestamp 1698431365
transform 1 0 2016 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_22
timestamp 1698431365
transform 1 0 3808 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_24
timestamp 1698431365
transform 1 0 4032 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_54
timestamp 1698431365
transform 1 0 7392 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_58
timestamp 1698431365
transform 1 0 7840 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_74
timestamp 1698431365
transform 1 0 9632 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_83
timestamp 1698431365
transform 1 0 10640 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_91
timestamp 1698431365
transform 1 0 11536 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_95
timestamp 1698431365
transform 1 0 11984 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_126
timestamp 1698431365
transform 1 0 15456 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_134
timestamp 1698431365
transform 1 0 16352 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_166
timestamp 1698431365
transform 1 0 19936 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_170
timestamp 1698431365
transform 1 0 20384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_186
timestamp 1698431365
transform 1 0 22176 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_190
timestamp 1698431365
transform 1 0 22624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_214
timestamp 1698431365
transform 1 0 25312 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_235
timestamp 1698431365
transform 1 0 27664 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_239
timestamp 1698431365
transform 1 0 28112 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_253
timestamp 1698431365
transform 1 0 29680 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_267
timestamp 1698431365
transform 1 0 31248 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_275
timestamp 1698431365
transform 1 0 32144 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_279
timestamp 1698431365
transform 1 0 32592 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_297
timestamp 1698431365
transform 1 0 34608 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_339
timestamp 1698431365
transform 1 0 39312 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_343
timestamp 1698431365
transform 1 0 39760 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_347
timestamp 1698431365
transform 1 0 40208 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_349
timestamp 1698431365
transform 1 0 40432 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_352
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_416
timestamp 1698431365
transform 1 0 47936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_10
timestamp 1698431365
transform 1 0 2464 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_26
timestamp 1698431365
transform 1 0 4256 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_41
timestamp 1698431365
transform 1 0 5936 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_46
timestamp 1698431365
transform 1 0 6496 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_48
timestamp 1698431365
transform 1 0 6720 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_51
timestamp 1698431365
transform 1 0 7056 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_53
timestamp 1698431365
transform 1 0 7280 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_56
timestamp 1698431365
transform 1 0 7616 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_67
timestamp 1698431365
transform 1 0 8848 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_71
timestamp 1698431365
transform 1 0 9296 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_104
timestamp 1698431365
transform 1 0 12992 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_138
timestamp 1698431365
transform 1 0 16800 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_174
timestamp 1698431365
transform 1 0 20832 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_181
timestamp 1698431365
transform 1 0 21616 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_185
timestamp 1698431365
transform 1 0 22064 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_235
timestamp 1698431365
transform 1 0 27664 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_270
timestamp 1698431365
transform 1 0 31584 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_335
timestamp 1698431365
transform 1 0 38864 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_339
timestamp 1698431365
transform 1 0 39312 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_371
timestamp 1698431365
transform 1 0 42896 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_379
timestamp 1698431365
transform 1 0 43792 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_383
timestamp 1698431365
transform 1 0 44240 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_403
timestamp 1698431365
transform 1 0 46480 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_411
timestamp 1698431365
transform 1 0 47376 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_415
timestamp 1698431365
transform 1 0 47824 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_66
timestamp 1698431365
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_146
timestamp 1698431365
transform 1 0 17696 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_203
timestamp 1698431365
transform 1 0 24080 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_207
timestamp 1698431365
transform 1 0 24528 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_209
timestamp 1698431365
transform 1 0 24752 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_216
timestamp 1698431365
transform 1 0 25536 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_248
timestamp 1698431365
transform 1 0 29120 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_252
timestamp 1698431365
transform 1 0 29568 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_270
timestamp 1698431365
transform 1 0 31584 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_272
timestamp 1698431365
transform 1 0 31808 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_278
timestamp 1698431365
transform 1 0 32480 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_327
timestamp 1698431365
transform 1 0 37968 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_343
timestamp 1698431365
transform 1 0 39760 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_347
timestamp 1698431365
transform 1 0 40208 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_349
timestamp 1698431365
transform 1 0 40432 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_352
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_416
timestamp 1698431365
transform 1 0 47936 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_2
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_6
timestamp 1698431365
transform 1 0 2016 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_22
timestamp 1698431365
transform 1 0 3808 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_30
timestamp 1698431365
transform 1 0 4704 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_43
timestamp 1698431365
transform 1 0 6160 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_47
timestamp 1698431365
transform 1 0 6608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_51
timestamp 1698431365
transform 1 0 7056 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_53
timestamp 1698431365
transform 1 0 7280 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_83
timestamp 1698431365
transform 1 0 10640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_87
timestamp 1698431365
transform 1 0 11088 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_103
timestamp 1698431365
transform 1 0 12880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_123
timestamp 1698431365
transform 1 0 15120 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_131
timestamp 1698431365
transform 1 0 16016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_135
timestamp 1698431365
transform 1 0 16464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_143
timestamp 1698431365
transform 1 0 17360 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_147
timestamp 1698431365
transform 1 0 17808 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_179
timestamp 1698431365
transform 1 0 21392 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_194
timestamp 1698431365
transform 1 0 23072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_196
timestamp 1698431365
transform 1 0 23296 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_215
timestamp 1698431365
transform 1 0 25424 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_219
timestamp 1698431365
transform 1 0 25872 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_235
timestamp 1698431365
transform 1 0 27664 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_243
timestamp 1698431365
transform 1 0 28560 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_255
timestamp 1698431365
transform 1 0 29904 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_271
timestamp 1698431365
transform 1 0 31696 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_273
timestamp 1698431365
transform 1 0 31920 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_294
timestamp 1698431365
transform 1 0 34272 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_310
timestamp 1698431365
transform 1 0 36064 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_314
timestamp 1698431365
transform 1 0 36512 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_419
timestamp 1698431365
transform 1 0 48272 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_10
timestamp 1698431365
transform 1 0 2464 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_18
timestamp 1698431365
transform 1 0 3360 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_22
timestamp 1698431365
transform 1 0 3808 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_52
timestamp 1698431365
transform 1 0 7168 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_56
timestamp 1698431365
transform 1 0 7616 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_64
timestamp 1698431365
transform 1 0 8512 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_78
timestamp 1698431365
transform 1 0 10080 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_85
timestamp 1698431365
transform 1 0 10864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_89
timestamp 1698431365
transform 1 0 11312 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_105
timestamp 1698431365
transform 1 0 13104 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_138
timestamp 1698431365
transform 1 0 16800 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_146
timestamp 1698431365
transform 1 0 17696 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_192
timestamp 1698431365
transform 1 0 22848 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_196
timestamp 1698431365
transform 1 0 23296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_220
timestamp 1698431365
transform 1 0 25984 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_224
timestamp 1698431365
transform 1 0 26432 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_228
timestamp 1698431365
transform 1 0 26880 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_232
timestamp 1698431365
transform 1 0 27328 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_240
timestamp 1698431365
transform 1 0 28224 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_244
timestamp 1698431365
transform 1 0 28672 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_250
timestamp 1698431365
transform 1 0 29344 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_258
timestamp 1698431365
transform 1 0 30240 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_266
timestamp 1698431365
transform 1 0 31136 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_274
timestamp 1698431365
transform 1 0 32032 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_278
timestamp 1698431365
transform 1 0 32480 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_346
timestamp 1698431365
transform 1 0 40096 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_6
timestamp 1698431365
transform 1 0 2016 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_14
timestamp 1698431365
transform 1 0 2912 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_16
timestamp 1698431365
transform 1 0 3136 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_19
timestamp 1698431365
transform 1 0 3472 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_27
timestamp 1698431365
transform 1 0 4368 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_31
timestamp 1698431365
transform 1 0 4816 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_41
timestamp 1698431365
transform 1 0 5936 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_57
timestamp 1698431365
transform 1 0 7728 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_65
timestamp 1698431365
transform 1 0 8624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_67
timestamp 1698431365
transform 1 0 8848 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_97
timestamp 1698431365
transform 1 0 12208 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_101
timestamp 1698431365
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_136
timestamp 1698431365
transform 1 0 16576 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_158
timestamp 1698431365
transform 1 0 19040 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_166
timestamp 1698431365
transform 1 0 19936 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_170
timestamp 1698431365
transform 1 0 20384 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_174
timestamp 1698431365
transform 1 0 20832 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_185
timestamp 1698431365
transform 1 0 22064 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_189
timestamp 1698431365
transform 1 0 22512 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_228
timestamp 1698431365
transform 1 0 26880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_236
timestamp 1698431365
transform 1 0 27776 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_238
timestamp 1698431365
transform 1 0 28000 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_249
timestamp 1698431365
transform 1 0 29232 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_279
timestamp 1698431365
transform 1 0 32592 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_281
timestamp 1698431365
transform 1 0 32816 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_288
timestamp 1698431365
transform 1 0 33600 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_304
timestamp 1698431365
transform 1 0 35392 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_312
timestamp 1698431365
transform 1 0 36288 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_314
timestamp 1698431365
transform 1 0 36512 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_419
timestamp 1698431365
transform 1 0 48272 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_33
timestamp 1698431365
transform 1 0 5040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_37
timestamp 1698431365
transform 1 0 5488 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_68
timestamp 1698431365
transform 1 0 8960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_76
timestamp 1698431365
transform 1 0 9856 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_80
timestamp 1698431365
transform 1 0 10304 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_110
timestamp 1698431365
transform 1 0 13664 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_200
timestamp 1698431365
transform 1 0 23744 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_204
timestamp 1698431365
transform 1 0 24192 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_294
timestamp 1698431365
transform 1 0 34272 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_326
timestamp 1698431365
transform 1 0 37856 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_342
timestamp 1698431365
transform 1 0 39648 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_416
timestamp 1698431365
transform 1 0 47936 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_18
timestamp 1698431365
transform 1 0 3360 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_22
timestamp 1698431365
transform 1 0 3808 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_30
timestamp 1698431365
transform 1 0 4704 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_53
timestamp 1698431365
transform 1 0 7280 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_61
timestamp 1698431365
transform 1 0 8176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_65
timestamp 1698431365
transform 1 0 8624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_67
timestamp 1698431365
transform 1 0 8848 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_70
timestamp 1698431365
transform 1 0 9184 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_102
timestamp 1698431365
transform 1 0 12768 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_104
timestamp 1698431365
transform 1 0 12992 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_109
timestamp 1698431365
transform 1 0 13552 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_112
timestamp 1698431365
transform 1 0 13888 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_128
timestamp 1698431365
transform 1 0 15680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_135
timestamp 1698431365
transform 1 0 16464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_139
timestamp 1698431365
transform 1 0 16912 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_142
timestamp 1698431365
transform 1 0 17248 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_160
timestamp 1698431365
transform 1 0 19264 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_168
timestamp 1698431365
transform 1 0 20160 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_170
timestamp 1698431365
transform 1 0 20384 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_173
timestamp 1698431365
transform 1 0 20720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_177
timestamp 1698431365
transform 1 0 21168 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_193
timestamp 1698431365
transform 1 0 22960 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_201
timestamp 1698431365
transform 1 0 23856 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_217
timestamp 1698431365
transform 1 0 25648 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_221
timestamp 1698431365
transform 1 0 26096 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_237
timestamp 1698431365
transform 1 0 27888 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_251
timestamp 1698431365
transform 1 0 29456 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_267
timestamp 1698431365
transform 1 0 31248 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_300
timestamp 1698431365
transform 1 0 34944 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_308
timestamp 1698431365
transform 1 0 35840 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_312
timestamp 1698431365
transform 1 0 36288 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_314
timestamp 1698431365
transform 1 0 36512 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_333
timestamp 1698431365
transform 1 0 38640 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_339
timestamp 1698431365
transform 1 0 39312 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_371
timestamp 1698431365
transform 1 0 42896 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_379
timestamp 1698431365
transform 1 0 43792 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_383
timestamp 1698431365
transform 1 0 44240 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_403
timestamp 1698431365
transform 1 0 46480 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_411
timestamp 1698431365
transform 1 0 47376 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_415
timestamp 1698431365
transform 1 0 47824 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_36
timestamp 1698431365
transform 1 0 5376 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_70
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_88
timestamp 1698431365
transform 1 0 11200 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_106
timestamp 1698431365
transform 1 0 13216 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_117
timestamp 1698431365
transform 1 0 14448 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_121
timestamp 1698431365
transform 1 0 14896 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_132
timestamp 1698431365
transform 1 0 16128 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_153
timestamp 1698431365
transform 1 0 18480 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_169
timestamp 1698431365
transform 1 0 20272 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_182
timestamp 1698431365
transform 1 0 21728 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_186
timestamp 1698431365
transform 1 0 22176 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_201
timestamp 1698431365
transform 1 0 23856 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_203
timestamp 1698431365
transform 1 0 24080 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_214
timestamp 1698431365
transform 1 0 25312 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_218
timestamp 1698431365
transform 1 0 25760 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_233
timestamp 1698431365
transform 1 0 27440 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_237
timestamp 1698431365
transform 1 0 27888 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_240
timestamp 1698431365
transform 1 0 28224 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_254
timestamp 1698431365
transform 1 0 29792 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_268
timestamp 1698431365
transform 1 0 31360 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_288
timestamp 1698431365
transform 1 0 33600 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_290
timestamp 1698431365
transform 1 0 33824 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_305
timestamp 1698431365
transform 1 0 35504 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_308
timestamp 1698431365
transform 1 0 35840 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_312
timestamp 1698431365
transform 1 0 36288 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_321
timestamp 1698431365
transform 1 0 37296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_325
timestamp 1698431365
transform 1 0 37744 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_337
timestamp 1698431365
transform 1 0 39088 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_339
timestamp 1698431365
transform 1 0 39312 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_356
timestamp 1698431365
transform 1 0 41216 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_360
timestamp 1698431365
transform 1 0 41664 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_369
timestamp 1698431365
transform 1 0 42672 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_373
timestamp 1698431365
transform 1 0 43120 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_376
timestamp 1698431365
transform 1 0 43456 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_385
timestamp 1698431365
transform 1 0 44464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_389
timestamp 1698431365
transform 1 0 44912 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_401
timestamp 1698431365
transform 1 0 46256 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_405
timestamp 1698431365
transform 1 0 46704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_407
timestamp 1698431365
transform 1 0 46928 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_410
timestamp 1698431365
transform 1 0 47264 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_414
timestamp 1698431365
transform 1 0 47712 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 2800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform 1 0 6832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input4
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 15568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input6
timestamp 1698431365
transform 1 0 2464 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input7
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform 1 0 3136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input11
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input12
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input14
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input15
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input16
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input17
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input18
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input19
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input21
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input24
timestamp 1698431365
transform -1 0 23632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input25
timestamp 1698431365
transform -1 0 27664 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698431365
transform -1 0 31696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 10864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 18928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input29
timestamp 1698431365
transform -1 0 46256 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input30
timestamp 1698431365
transform -1 0 44464 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input31
timestamp 1698431365
transform -1 0 42672 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input32
timestamp 1698431365
transform -1 0 41216 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input33
timestamp 1698431365
transform -1 0 39088 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input34
timestamp 1698431365
transform -1 0 37296 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input35
timestamp 1698431365
transform -1 0 35504 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input36
timestamp 1698431365
transform 1 0 33376 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_97 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_98
timestamp 1698431365
transform 1 0 47936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_99
timestamp 1698431365
transform 1 0 47936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_100
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_101
timestamp 1698431365
transform 1 0 47936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_102
timestamp 1698431365
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_103
timestamp 1698431365
transform 1 0 47936 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_104
timestamp 1698431365
transform 1 0 47936 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_105
timestamp 1698431365
transform 1 0 47936 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_106
timestamp 1698431365
transform 1 0 47936 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_107
timestamp 1698431365
transform 1 0 47936 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_108
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_109
timestamp 1698431365
transform 1 0 47936 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  interp_tri_110
timestamp 1698431365
transform 1 0 47936 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3584 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38
timestamp 1698431365
transform 1 0 45472 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output39
timestamp 1698431365
transform 1 0 46816 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output40
timestamp 1698431365
transform 1 0 46816 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output41
timestamp 1698431365
transform 1 0 46816 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output42
timestamp 1698431365
transform 1 0 46816 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output43
timestamp 1698431365
transform 1 0 46816 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output44
timestamp 1698431365
transform 1 0 46816 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output45
timestamp 1698431365
transform 1 0 46816 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output46
timestamp 1698431365
transform 1 0 46816 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output47
timestamp 1698431365
transform 1 0 46816 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output48
timestamp 1698431365
transform 1 0 46816 0 1 58016
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output49
timestamp 1698431365
transform 1 0 46816 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output50
timestamp 1698431365
transform 1 0 46816 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output51
timestamp 1698431365
transform 1 0 46816 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output52
timestamp 1698431365
transform 1 0 46816 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698431365
transform 1 0 46816 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output54
timestamp 1698431365
transform 1 0 46816 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output55
timestamp 1698431365
transform 1 0 46816 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output56
timestamp 1698431365
transform 1 0 46816 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output57
timestamp 1698431365
transform 1 0 16912 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output58
timestamp 1698431365
transform 1 0 15008 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output59
timestamp 1698431365
transform 1 0 13328 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output60
timestamp 1698431365
transform -1 0 12768 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698431365
transform -1 0 11200 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output62
timestamp 1698431365
transform -1 0 8960 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output63
timestamp 1698431365
transform -1 0 7392 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output64
timestamp 1698431365
transform 1 0 3584 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output65
timestamp 1698431365
transform -1 0 33600 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output66
timestamp 1698431365
transform -1 0 31360 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output67
timestamp 1698431365
transform 1 0 28672 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output68
timestamp 1698431365
transform -1 0 27440 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output69
timestamp 1698431365
transform -1 0 25648 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output70
timestamp 1698431365
transform 1 0 22288 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output71
timestamp 1698431365
transform 1 0 20608 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output72
timestamp 1698431365
transform -1 0 20272 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 48608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 48608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 48608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 48608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 48608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 48608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 48608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 48608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 48608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 48608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 48608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 48608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 48608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 48608 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 48608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 48608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 48608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 48608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 48608 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 48608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 48608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 48608 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 48608 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 48608 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 48608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 48608 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 48608 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 48608 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 48608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 48608 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 48608 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 48608 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 48608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 48608 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 48608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 48608 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 48608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 48608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer1
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer2
timestamp 1698431365
transform -1 0 23856 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer3
timestamp 1698431365
transform -1 0 37744 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer4
timestamp 1698431365
transform -1 0 39312 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer5
timestamp 1698431365
transform -1 0 33488 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer6
timestamp 1698431365
transform -1 0 32144 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer7
timestamp 1698431365
transform -1 0 40208 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer8
timestamp 1698431365
transform -1 0 11424 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer9
timestamp 1698431365
transform -1 0 22288 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer10
timestamp 1698431365
transform -1 0 17920 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer11
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer12
timestamp 1698431365
transform -1 0 23632 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer13
timestamp 1698431365
transform 1 0 27104 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  rebuffer14 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18704 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer15
timestamp 1698431365
transform -1 0 19264 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer16
timestamp 1698431365
transform -1 0 22960 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer17
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer18
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer19
timestamp 1698431365
transform 1 0 37184 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer20
timestamp 1698431365
transform -1 0 15008 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer21
timestamp 1698431365
transform -1 0 10528 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer22
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer23
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer24
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39536 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer26
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer27
timestamp 1698431365
transform 1 0 12656 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer28
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer29
timestamp 1698431365
transform 1 0 16016 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_200
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_201
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_202
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_203
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_204
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_205
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_206
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_207
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_208
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_209
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_210
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_211
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_212
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_213
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_214
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_215
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_216
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_217
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_218
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_219
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_220
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_221
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_222
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_223
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_224
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_225
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_226
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_227
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_228
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_229
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_230
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_231
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_232
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_233
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_234
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_235
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_236
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_237
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_238
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_239
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_240
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_241
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_242
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_243
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_244
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_245
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_246
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_247
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_248
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_249
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_250
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_251
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_252
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_253
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_254
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_255
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_256
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_257
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_258
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_259
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_260
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_261
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_262
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_263
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_264
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_265
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_266
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_267
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_268
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_269
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_270
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_271
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_272
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_273
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_274
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_275
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_276
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_277
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_278
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_279
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_280
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_281
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_282
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_283
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_284
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_285
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_286
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_287
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_288
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_289
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_290
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_291
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_292
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_293
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_294
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_295
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_296
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_297
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_298
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_299
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_300
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_301
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_302
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_303
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_304
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_305
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_306
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_307
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_308
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_309
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_310
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_311
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_312
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_313
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_314
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_315
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_316
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_317
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_318
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_319
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_320
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_321
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_322
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_323
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_324
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_325
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_326
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_327
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_328
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_329
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_330
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_331
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_332
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_333
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_334
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_335
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_336
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_337
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_338
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_339
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_340
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_341
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_342
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_343
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_344
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_345
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_346
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_347
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_348
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_349
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_350
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_351
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_352
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_353
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_354
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_355
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_356
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_357
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_358
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_360
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_361
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_362
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_363
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_364
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_367
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_368
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_369
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_374
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_375
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_387
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_392
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_393
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_394
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_398
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_399
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_400
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_401
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_403
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_404
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_405
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_406
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_407
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_408
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_409
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_410
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_411
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_412
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_413
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_414
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_415
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_416
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_417
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_418
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_419
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_420
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_421
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_422
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_423
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_424
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_425
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_426
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_427
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_428
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_429
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_430
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_431
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_432
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_433
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_434
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_435
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_436
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_437
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_438
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_439
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_440
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_441
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_442
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_443
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_444
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_445
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_446
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_447
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_448
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_449
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_450
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_451
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_452
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_453
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_454
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_455
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_456
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_457
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_458
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_459
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_460
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_461
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_462
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_463
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_464
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_465
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_466
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_467
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_468
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_469
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_470
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_471
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_472
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_473
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_474
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_475
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_476
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_477
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_478
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_479
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_480
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_481
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_482
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_483
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_484
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_485
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_486
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_487
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_488
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_489
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_490
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_491
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_492
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_493
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_494
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_495
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_496
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_497
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_498
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_499
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_500
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_501
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_502
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_503
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_504
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_505
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_506
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_507
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_508
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_509
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_510
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_511
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_512
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_513
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_514
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_515
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_516
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_517
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_518
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_519
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_520
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_521
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_522
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_523
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_524
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_525
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_526
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_527
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_528
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_529
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_530
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_531
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_532
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_533
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_534
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_535
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_536
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_537
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_538
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_539
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_540
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_541
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_542
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_543
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_544
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_545
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_546
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_547
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_548
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_549
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_550
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_551
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_552
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_553
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_554
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_555
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_556
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_557
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_558
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_559
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_560
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_561
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_562
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_563
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_564
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_565
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_566
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_567
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_568
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_569
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_570
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_571
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_572
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_573
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_574
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_575
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_576
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_577
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_578
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_579
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_580
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_581
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_582
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_583
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_584
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_585
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_586
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_587
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_588
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_589
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_590
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_591
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_592
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_593
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_594
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_595
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_596
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_597
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_598
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_599
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_600
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_601
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_602
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_603
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_604
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_605
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_606
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_607
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_608
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_609
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_610
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_611
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_612
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_613
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_614
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_615
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_616
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_617
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_618
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_619
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_620
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_621
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_622
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_623
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_624
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_625
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_626
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_627
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_628
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_629
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_630
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_631
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_632
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_633
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_634
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_635
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_636
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_637
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_638
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_639
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_640
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_641
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_642
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_643
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_644
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_645
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_646
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_647
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_648
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_649
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_650
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_651
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_652
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_653
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_654
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_655
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_656
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_657
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_658
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_659
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_660
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_661
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_662
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_663
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_664
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_665
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_666
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_667
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_668
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_669
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_670
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_671
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_672
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_673
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_674
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_675
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_676
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_677
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_678
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_679
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_680
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_681
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_682
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_683
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_684
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_685
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_686
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_687
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_688
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_689
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_690
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_691
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_692
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_693
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_694
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_695
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_696
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_697
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_698
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_699
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_700
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_701
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_702
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_703
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_704
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_705
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_706
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_707
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_708
timestamp 1698431365
transform 1 0 12768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_709
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_710
timestamp 1698431365
transform 1 0 20384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_711
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_712
timestamp 1698431365
transform 1 0 28000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_713
timestamp 1698431365
transform 1 0 31808 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_714
timestamp 1698431365
transform 1 0 35616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_715
timestamp 1698431365
transform 1 0 39424 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_716
timestamp 1698431365
transform 1 0 43232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_717
timestamp 1698431365
transform 1 0 47040 0 -1 76832
box -86 -86 310 870
<< labels >>
flabel metal2 s 2464 79200 2576 80000 0 FreeSans 448 90 0 0 active
port 0 nsew signal tristate
flabel metal2 s 47264 79200 47376 80000 0 FreeSans 448 90 0 0 clk
port 1 nsew signal input
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 2 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 2 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 3 nsew ground bidirectional
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 wb_clk_i
port 4 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 wb_rst_i
port 5 nsew signal input
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 6 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 7 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 8 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 9 nsew signal input
flabel metal3 s 0 77952 800 78064 0 FreeSans 448 0 0 0 wbs_dat_i[0]
port 10 nsew signal input
flabel metal3 s 0 53312 800 53424 0 FreeSans 448 0 0 0 wbs_dat_i[10]
port 11 nsew signal input
flabel metal3 s 0 50848 800 50960 0 FreeSans 448 0 0 0 wbs_dat_i[11]
port 12 nsew signal input
flabel metal3 s 0 48384 800 48496 0 FreeSans 448 0 0 0 wbs_dat_i[12]
port 13 nsew signal input
flabel metal3 s 0 45920 800 46032 0 FreeSans 448 0 0 0 wbs_dat_i[13]
port 14 nsew signal input
flabel metal3 s 0 43456 800 43568 0 FreeSans 448 0 0 0 wbs_dat_i[14]
port 15 nsew signal input
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 wbs_dat_i[15]
port 16 nsew signal input
flabel metal3 s 0 38528 800 38640 0 FreeSans 448 0 0 0 wbs_dat_i[16]
port 17 nsew signal input
flabel metal3 s 0 36064 800 36176 0 FreeSans 448 0 0 0 wbs_dat_i[17]
port 18 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 wbs_dat_i[18]
port 19 nsew signal input
flabel metal3 s 0 31136 800 31248 0 FreeSans 448 0 0 0 wbs_dat_i[19]
port 20 nsew signal input
flabel metal3 s 0 75488 800 75600 0 FreeSans 448 0 0 0 wbs_dat_i[1]
port 21 nsew signal input
flabel metal3 s 0 28672 800 28784 0 FreeSans 448 0 0 0 wbs_dat_i[20]
port 22 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 wbs_dat_i[21]
port 23 nsew signal input
flabel metal3 s 0 23744 800 23856 0 FreeSans 448 0 0 0 wbs_dat_i[22]
port 24 nsew signal input
flabel metal3 s 0 21280 800 21392 0 FreeSans 448 0 0 0 wbs_dat_i[23]
port 25 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 wbs_dat_i[24]
port 26 nsew signal input
flabel metal3 s 0 16352 800 16464 0 FreeSans 448 0 0 0 wbs_dat_i[25]
port 27 nsew signal input
flabel metal3 s 0 13888 800 14000 0 FreeSans 448 0 0 0 wbs_dat_i[26]
port 28 nsew signal input
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 wbs_dat_i[27]
port 29 nsew signal input
flabel metal3 s 0 8960 800 9072 0 FreeSans 448 0 0 0 wbs_dat_i[28]
port 30 nsew signal input
flabel metal3 s 0 6496 800 6608 0 FreeSans 448 0 0 0 wbs_dat_i[29]
port 31 nsew signal input
flabel metal3 s 0 73024 800 73136 0 FreeSans 448 0 0 0 wbs_dat_i[2]
port 32 nsew signal input
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 wbs_dat_i[30]
port 33 nsew signal input
flabel metal3 s 0 1568 800 1680 0 FreeSans 448 0 0 0 wbs_dat_i[31]
port 34 nsew signal input
flabel metal3 s 0 70560 800 70672 0 FreeSans 448 0 0 0 wbs_dat_i[3]
port 35 nsew signal input
flabel metal3 s 0 68096 800 68208 0 FreeSans 448 0 0 0 wbs_dat_i[4]
port 36 nsew signal input
flabel metal3 s 0 65632 800 65744 0 FreeSans 448 0 0 0 wbs_dat_i[5]
port 37 nsew signal input
flabel metal3 s 0 63168 800 63280 0 FreeSans 448 0 0 0 wbs_dat_i[6]
port 38 nsew signal input
flabel metal3 s 0 60704 800 60816 0 FreeSans 448 0 0 0 wbs_dat_i[7]
port 39 nsew signal input
flabel metal3 s 0 58240 800 58352 0 FreeSans 448 0 0 0 wbs_dat_i[8]
port 40 nsew signal input
flabel metal3 s 0 55776 800 55888 0 FreeSans 448 0 0 0 wbs_dat_i[9]
port 41 nsew signal input
flabel metal3 s 49200 1568 50000 1680 0 FreeSans 448 0 0 0 wbs_dat_o[0]
port 42 nsew signal tristate
flabel metal3 s 49200 26208 50000 26320 0 FreeSans 448 0 0 0 wbs_dat_o[10]
port 43 nsew signal tristate
flabel metal3 s 49200 28672 50000 28784 0 FreeSans 448 0 0 0 wbs_dat_o[11]
port 44 nsew signal tristate
flabel metal3 s 49200 31136 50000 31248 0 FreeSans 448 0 0 0 wbs_dat_o[12]
port 45 nsew signal tristate
flabel metal3 s 49200 33600 50000 33712 0 FreeSans 448 0 0 0 wbs_dat_o[13]
port 46 nsew signal tristate
flabel metal3 s 49200 36064 50000 36176 0 FreeSans 448 0 0 0 wbs_dat_o[14]
port 47 nsew signal tristate
flabel metal3 s 49200 38528 50000 38640 0 FreeSans 448 0 0 0 wbs_dat_o[15]
port 48 nsew signal tristate
flabel metal3 s 49200 40992 50000 41104 0 FreeSans 448 0 0 0 wbs_dat_o[16]
port 49 nsew signal tristate
flabel metal3 s 49200 43456 50000 43568 0 FreeSans 448 0 0 0 wbs_dat_o[17]
port 50 nsew signal tristate
flabel metal3 s 49200 45920 50000 46032 0 FreeSans 448 0 0 0 wbs_dat_o[18]
port 51 nsew signal tristate
flabel metal3 s 49200 48384 50000 48496 0 FreeSans 448 0 0 0 wbs_dat_o[19]
port 52 nsew signal tristate
flabel metal3 s 49200 4032 50000 4144 0 FreeSans 448 0 0 0 wbs_dat_o[1]
port 53 nsew signal tristate
flabel metal3 s 49200 50848 50000 50960 0 FreeSans 448 0 0 0 wbs_dat_o[20]
port 54 nsew signal tristate
flabel metal3 s 49200 53312 50000 53424 0 FreeSans 448 0 0 0 wbs_dat_o[21]
port 55 nsew signal tristate
flabel metal3 s 49200 55776 50000 55888 0 FreeSans 448 0 0 0 wbs_dat_o[22]
port 56 nsew signal tristate
flabel metal3 s 49200 58240 50000 58352 0 FreeSans 448 0 0 0 wbs_dat_o[23]
port 57 nsew signal tristate
flabel metal3 s 49200 60704 50000 60816 0 FreeSans 448 0 0 0 wbs_dat_o[24]
port 58 nsew signal tristate
flabel metal3 s 49200 63168 50000 63280 0 FreeSans 448 0 0 0 wbs_dat_o[25]
port 59 nsew signal tristate
flabel metal3 s 49200 65632 50000 65744 0 FreeSans 448 0 0 0 wbs_dat_o[26]
port 60 nsew signal tristate
flabel metal3 s 49200 68096 50000 68208 0 FreeSans 448 0 0 0 wbs_dat_o[27]
port 61 nsew signal tristate
flabel metal3 s 49200 70560 50000 70672 0 FreeSans 448 0 0 0 wbs_dat_o[28]
port 62 nsew signal tristate
flabel metal3 s 49200 73024 50000 73136 0 FreeSans 448 0 0 0 wbs_dat_o[29]
port 63 nsew signal tristate
flabel metal3 s 49200 6496 50000 6608 0 FreeSans 448 0 0 0 wbs_dat_o[2]
port 64 nsew signal tristate
flabel metal3 s 49200 75488 50000 75600 0 FreeSans 448 0 0 0 wbs_dat_o[30]
port 65 nsew signal tristate
flabel metal3 s 49200 77952 50000 78064 0 FreeSans 448 0 0 0 wbs_dat_o[31]
port 66 nsew signal tristate
flabel metal3 s 49200 8960 50000 9072 0 FreeSans 448 0 0 0 wbs_dat_o[3]
port 67 nsew signal tristate
flabel metal3 s 49200 11424 50000 11536 0 FreeSans 448 0 0 0 wbs_dat_o[4]
port 68 nsew signal tristate
flabel metal3 s 49200 13888 50000 14000 0 FreeSans 448 0 0 0 wbs_dat_o[5]
port 69 nsew signal tristate
flabel metal3 s 49200 16352 50000 16464 0 FreeSans 448 0 0 0 wbs_dat_o[6]
port 70 nsew signal tristate
flabel metal3 s 49200 18816 50000 18928 0 FreeSans 448 0 0 0 wbs_dat_o[7]
port 71 nsew signal tristate
flabel metal3 s 49200 21280 50000 21392 0 FreeSans 448 0 0 0 wbs_dat_o[8]
port 72 nsew signal tristate
flabel metal3 s 49200 23744 50000 23856 0 FreeSans 448 0 0 0 wbs_dat_o[9]
port 73 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 74 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 75 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 76 nsew signal input
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 77 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 78 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_we_i
port 79 nsew signal input
flabel metal2 s 16800 79200 16912 80000 0 FreeSans 448 90 0 0 x_end[0]
port 80 nsew signal tristate
flabel metal2 s 15008 79200 15120 80000 0 FreeSans 448 90 0 0 x_end[1]
port 81 nsew signal tristate
flabel metal2 s 13216 79200 13328 80000 0 FreeSans 448 90 0 0 x_end[2]
port 82 nsew signal tristate
flabel metal2 s 11424 79200 11536 80000 0 FreeSans 448 90 0 0 x_end[3]
port 83 nsew signal tristate
flabel metal2 s 9632 79200 9744 80000 0 FreeSans 448 90 0 0 x_end[4]
port 84 nsew signal tristate
flabel metal2 s 7840 79200 7952 80000 0 FreeSans 448 90 0 0 x_end[5]
port 85 nsew signal tristate
flabel metal2 s 6048 79200 6160 80000 0 FreeSans 448 90 0 0 x_end[6]
port 86 nsew signal tristate
flabel metal2 s 4256 79200 4368 80000 0 FreeSans 448 90 0 0 x_end[7]
port 87 nsew signal tristate
flabel metal2 s 31136 79200 31248 80000 0 FreeSans 448 90 0 0 x_start[0]
port 88 nsew signal tristate
flabel metal2 s 29344 79200 29456 80000 0 FreeSans 448 90 0 0 x_start[1]
port 89 nsew signal tristate
flabel metal2 s 27552 79200 27664 80000 0 FreeSans 448 90 0 0 x_start[2]
port 90 nsew signal tristate
flabel metal2 s 25760 79200 25872 80000 0 FreeSans 448 90 0 0 x_start[3]
port 91 nsew signal tristate
flabel metal2 s 23968 79200 24080 80000 0 FreeSans 448 90 0 0 x_start[4]
port 92 nsew signal tristate
flabel metal2 s 22176 79200 22288 80000 0 FreeSans 448 90 0 0 x_start[5]
port 93 nsew signal tristate
flabel metal2 s 20384 79200 20496 80000 0 FreeSans 448 90 0 0 x_start[6]
port 94 nsew signal tristate
flabel metal2 s 18592 79200 18704 80000 0 FreeSans 448 90 0 0 x_start[7]
port 95 nsew signal tristate
flabel metal2 s 45472 79200 45584 80000 0 FreeSans 448 90 0 0 y[0]
port 96 nsew signal input
flabel metal2 s 43680 79200 43792 80000 0 FreeSans 448 90 0 0 y[1]
port 97 nsew signal input
flabel metal2 s 41888 79200 42000 80000 0 FreeSans 448 90 0 0 y[2]
port 98 nsew signal input
flabel metal2 s 40096 79200 40208 80000 0 FreeSans 448 90 0 0 y[3]
port 99 nsew signal input
flabel metal2 s 38304 79200 38416 80000 0 FreeSans 448 90 0 0 y[4]
port 100 nsew signal input
flabel metal2 s 36512 79200 36624 80000 0 FreeSans 448 90 0 0 y[5]
port 101 nsew signal input
flabel metal2 s 34720 79200 34832 80000 0 FreeSans 448 90 0 0 y[6]
port 102 nsew signal input
flabel metal2 s 32928 79200 33040 80000 0 FreeSans 448 90 0 0 y[7]
port 103 nsew signal input
rlabel metal1 24976 76048 24976 76048 0 vdd
rlabel metal1 24976 76832 24976 76832 0 vss
rlabel metal2 5992 68432 5992 68432 0 _0000_
rlabel metal2 33096 74760 33096 74760 0 _0001_
rlabel metal2 30632 73752 30632 73752 0 _0002_
rlabel metal2 26712 74144 26712 74144 0 _0003_
rlabel metal2 28616 74368 28616 74368 0 _0004_
rlabel metal3 24584 74200 24584 74200 0 _0005_
rlabel metal2 27272 74368 27272 74368 0 _0006_
rlabel metal2 19432 74368 19432 74368 0 _0007_
rlabel metal2 25816 31808 25816 31808 0 _0008_
rlabel metal2 14728 75320 14728 75320 0 _0009_
rlabel metal2 26376 74144 26376 74144 0 _0010_
rlabel metal2 11592 74760 11592 74760 0 _0011_
rlabel metal2 9968 73976 9968 73976 0 _0012_
rlabel metal2 8344 73024 8344 73024 0 _0013_
rlabel metal3 6048 74984 6048 74984 0 _0014_
rlabel metal2 5656 72800 5656 72800 0 _0015_
rlabel metal2 4256 73976 4256 73976 0 _0016_
rlabel metal2 5096 65800 5096 65800 0 _0017_
rlabel metal2 4088 61208 4088 61208 0 _0018_
rlabel metal2 2744 57344 2744 57344 0 _0019_
rlabel metal2 2408 52808 2408 52808 0 _0020_
rlabel metal2 6440 46368 6440 46368 0 _0021_
rlabel metal2 5656 39004 5656 39004 0 _0022_
rlabel metal2 2520 35168 2520 35168 0 _0023_
rlabel metal2 2632 30464 2632 30464 0 _0024_
rlabel metal2 6440 26600 6440 26600 0 _0025_
rlabel metal2 5768 21056 5768 21056 0 _0026_
rlabel metal2 2520 29288 2520 29288 0 _0027_
rlabel metal2 2800 26376 2800 26376 0 _0028_
rlabel metal2 9688 58408 9688 58408 0 _0029_
rlabel metal2 9800 56616 9800 56616 0 _0030_
rlabel metal2 2576 50792 2576 50792 0 _0031_
rlabel metal2 9800 53368 9800 53368 0 _0032_
rlabel metal2 2520 48664 2520 48664 0 _0033_
rlabel metal2 2408 40488 2408 40488 0 _0034_
rlabel metal2 2576 39704 2576 39704 0 _0035_
rlabel metal2 9632 40040 9632 40040 0 _0036_
rlabel metal2 8736 66136 8736 66136 0 _0037_
rlabel metal2 10864 43624 10864 43624 0 _0038_
rlabel metal2 11648 38920 11648 38920 0 _0039_
rlabel metal2 12264 45416 12264 45416 0 _0040_
rlabel metal2 16072 42728 16072 42728 0 _0041_
rlabel metal2 12488 41188 12488 41188 0 _0042_
rlabel metal2 14336 39704 14336 39704 0 _0043_
rlabel metal2 16072 39788 16072 39788 0 _0044_
rlabel metal2 18200 40656 18200 40656 0 _0045_
rlabel metal2 12040 61096 12040 61096 0 _0046_
rlabel metal2 11368 68152 11368 68152 0 _0047_
rlabel metal2 12264 65688 12264 65688 0 _0048_
rlabel metal2 11368 65016 11368 65016 0 _0049_
rlabel metal2 16744 60592 16744 60592 0 _0050_
rlabel metal2 21896 60368 21896 60368 0 _0051_
rlabel metal2 22568 62188 22568 62188 0 _0052_
rlabel metal2 20104 60368 20104 60368 0 _0053_
rlabel metal3 25704 59976 25704 59976 0 _0054_
rlabel metal2 26152 58632 26152 58632 0 _0055_
rlabel metal3 28560 53704 28560 53704 0 _0056_
rlabel metal3 25816 54432 25816 54432 0 _0057_
rlabel metal2 28168 53256 28168 53256 0 _0058_
rlabel metal2 24360 48664 24360 48664 0 _0059_
rlabel metal2 25368 36064 25368 36064 0 _0060_
rlabel metal2 24920 16240 24920 16240 0 _0061_
rlabel metal2 13160 68992 13160 68992 0 _0062_
rlabel metal2 14560 70840 14560 70840 0 _0063_
rlabel metal2 14952 67648 14952 67648 0 _0064_
rlabel metal2 14504 72128 14504 72128 0 _0065_
rlabel metal2 17024 66136 17024 66136 0 _0066_
rlabel metal3 22120 66136 22120 66136 0 _0067_
rlabel metal2 20888 65520 20888 65520 0 _0068_
rlabel metal2 18704 67704 18704 67704 0 _0069_
rlabel metal2 25368 49056 25368 49056 0 _0070_
rlabel metal3 26432 46536 26432 46536 0 _0071_
rlabel metal3 26544 45192 26544 45192 0 _0072_
rlabel metal3 26320 43400 26320 43400 0 _0073_
rlabel metal3 26432 41832 26432 41832 0 _0074_
rlabel metal2 26600 40432 26600 40432 0 _0075_
rlabel metal2 26264 18088 26264 18088 0 _0076_
rlabel metal2 22624 18424 22624 18424 0 _0077_
rlabel metal2 14168 48384 14168 48384 0 _0078_
rlabel metal2 15624 52696 15624 52696 0 _0079_
rlabel metal2 15064 54096 15064 54096 0 _0080_
rlabel metal2 14336 57848 14336 57848 0 _0081_
rlabel metal2 12152 57008 12152 57008 0 _0082_
rlabel metal2 11928 54936 11928 54936 0 _0083_
rlabel metal2 11816 51688 11816 51688 0 _0084_
rlabel metal2 10808 48664 10808 48664 0 _0085_
rlabel metal2 21784 6216 21784 6216 0 _0086_
rlabel metal2 19880 5488 19880 5488 0 _0087_
rlabel metal2 18536 6496 18536 6496 0 _0088_
rlabel metal2 18592 6664 18592 6664 0 _0089_
rlabel metal2 15960 7784 15960 7784 0 _0090_
rlabel metal2 16016 12152 16016 12152 0 _0091_
rlabel metal2 13496 6160 13496 6160 0 _0092_
rlabel metal2 15064 5488 15064 5488 0 _0093_
rlabel metal2 16744 5936 16744 5936 0 _0094_
rlabel metal2 15512 12936 15512 12936 0 _0095_
rlabel metal2 21112 13664 21112 13664 0 _0096_
rlabel metal2 21224 13944 21224 13944 0 _0097_
rlabel metal2 20384 13720 20384 13720 0 _0098_
rlabel metal3 20048 21336 20048 21336 0 _0099_
rlabel metal2 17640 9632 17640 9632 0 _0100_
rlabel metal2 18424 6048 18424 6048 0 _0101_
rlabel metal2 18816 5208 18816 5208 0 _0102_
rlabel metal2 19152 5320 19152 5320 0 _0103_
rlabel metal2 20552 5264 20552 5264 0 _0104_
rlabel metal2 21560 5152 21560 5152 0 _0105_
rlabel metal2 23800 4760 23800 4760 0 _0106_
rlabel metal2 27888 6776 27888 6776 0 _0107_
rlabel metal2 24696 12824 24696 12824 0 _0108_
rlabel metal2 26936 10080 26936 10080 0 _0109_
rlabel metal2 26936 7672 26936 7672 0 _0110_
rlabel metal2 27776 7336 27776 7336 0 _0111_
rlabel metal2 28056 4928 28056 4928 0 _0112_
rlabel metal3 41272 5992 41272 5992 0 _0113_
rlabel metal2 42840 20104 42840 20104 0 _0114_
rlabel metal2 29904 11480 29904 11480 0 _0115_
rlabel metal3 39256 18424 39256 18424 0 _0116_
rlabel metal3 41048 18536 41048 18536 0 _0117_
rlabel metal2 42112 16744 42112 16744 0 _0118_
rlabel metal2 41944 5880 41944 5880 0 _0119_
rlabel metal2 43512 7504 43512 7504 0 _0120_
rlabel metal2 44968 18760 44968 18760 0 _0121_
rlabel metal2 45584 20104 45584 20104 0 _0122_
rlabel metal2 28616 20384 28616 20384 0 _0123_
rlabel metal2 27048 21224 27048 21224 0 _0124_
rlabel metal2 1288 47040 1288 47040 0 _0125_
rlabel metal2 45192 20048 45192 20048 0 _0126_
rlabel metal3 25816 19208 25816 19208 0 _0127_
rlabel metal2 25592 19712 25592 19712 0 _0128_
rlabel metal2 42672 9016 42672 9016 0 _0129_
rlabel metal3 43736 9016 43736 9016 0 _0130_
rlabel metal2 41496 6888 41496 6888 0 _0131_
rlabel metal2 22680 4256 22680 4256 0 _0132_
rlabel metal2 23576 4536 23576 4536 0 _0133_
rlabel metal2 20552 5880 20552 5880 0 _0134_
rlabel metal2 22344 5768 22344 5768 0 _0135_
rlabel metal2 22904 6944 22904 6944 0 _0136_
rlabel metal2 23128 5488 23128 5488 0 _0137_
rlabel metal2 16072 12768 16072 12768 0 _0138_
rlabel metal3 23744 15288 23744 15288 0 _0139_
rlabel metal3 22736 15400 22736 15400 0 _0140_
rlabel metal2 22848 14280 22848 14280 0 _0141_
rlabel metal2 22904 14784 22904 14784 0 _0142_
rlabel metal2 17080 13720 17080 13720 0 _0143_
rlabel metal2 16184 12600 16184 12600 0 _0144_
rlabel metal2 16520 6384 16520 6384 0 _0145_
rlabel metal2 15960 5600 15960 5600 0 _0146_
rlabel metal2 17304 5376 17304 5376 0 _0147_
rlabel metal2 17976 5096 17976 5096 0 _0148_
rlabel metal2 28728 5656 28728 5656 0 _0149_
rlabel metal2 27832 7896 27832 7896 0 _0150_
rlabel metal3 28392 7672 28392 7672 0 _0151_
rlabel metal2 27272 7560 27272 7560 0 _0152_
rlabel metal3 29932 8008 29932 8008 0 _0153_
rlabel metal2 41384 6776 41384 6776 0 _0154_
rlabel metal2 42000 7672 42000 7672 0 _0155_
rlabel metal3 38864 9688 38864 9688 0 _0156_
rlabel metal2 35560 11424 35560 11424 0 _0157_
rlabel metal3 38136 15512 38136 15512 0 _0158_
rlabel metal2 39704 5208 39704 5208 0 _0159_
rlabel metal2 38752 4536 38752 4536 0 _0160_
rlabel metal2 39256 5096 39256 5096 0 _0161_
rlabel metal2 38976 4312 38976 4312 0 _0162_
rlabel metal2 39256 10136 39256 10136 0 _0163_
rlabel metal2 41160 17836 41160 17836 0 _0164_
rlabel metal2 40152 8904 40152 8904 0 _0165_
rlabel metal2 39928 7280 39928 7280 0 _0166_
rlabel metal2 39032 10808 39032 10808 0 _0167_
rlabel metal3 26768 20552 26768 20552 0 _0168_
rlabel metal2 26040 20328 26040 20328 0 _0169_
rlabel metal2 3696 73976 3696 73976 0 _0170_
rlabel metal2 25032 69832 25032 69832 0 _0171_
rlabel metal2 6104 62328 6104 62328 0 _0172_
rlabel metal2 6776 60200 6776 60200 0 _0173_
rlabel metal2 5768 62188 5768 62188 0 _0174_
rlabel metal2 4928 62328 4928 62328 0 _0175_
rlabel metal2 5992 58408 5992 58408 0 _0176_
rlabel metal2 6104 58576 6104 58576 0 _0177_
rlabel metal2 4648 57904 4648 57904 0 _0178_
rlabel metal2 3752 57624 3752 57624 0 _0179_
rlabel metal3 7952 57512 7952 57512 0 _0180_
rlabel metal2 6664 57176 6664 57176 0 _0181_
rlabel metal2 5992 53256 5992 53256 0 _0182_
rlabel metal2 2744 51744 2744 51744 0 _0183_
rlabel metal2 4424 47376 4424 47376 0 _0184_
rlabel metal2 6664 52584 6664 52584 0 _0185_
rlabel metal2 4984 52640 4984 52640 0 _0186_
rlabel metal2 4872 46872 4872 46872 0 _0187_
rlabel metal3 5600 46760 5600 46760 0 _0188_
rlabel metal3 4704 42728 4704 42728 0 _0189_
rlabel metal2 4984 46424 4984 46424 0 _0190_
rlabel metal2 4368 45864 4368 45864 0 _0191_
rlabel metal2 4536 43680 4536 43680 0 _0192_
rlabel metal2 4984 41776 4984 41776 0 _0193_
rlabel metal2 5096 42000 5096 42000 0 _0194_
rlabel metal2 4704 42056 4704 42056 0 _0195_
rlabel metal2 5152 41720 5152 41720 0 _0196_
rlabel metal2 2296 35224 2296 35224 0 _0197_
rlabel metal2 6888 31472 6888 31472 0 _0198_
rlabel metal2 4760 35112 4760 35112 0 _0199_
rlabel metal3 5656 36232 5656 36232 0 _0200_
rlabel metal2 5544 32928 5544 32928 0 _0201_
rlabel metal2 2968 30520 2968 30520 0 _0202_
rlabel metal3 5152 25480 5152 25480 0 _0203_
rlabel metal2 5656 29792 5656 29792 0 _0204_
rlabel metal2 5992 29904 5992 29904 0 _0205_
rlabel metal2 5208 24976 5208 24976 0 _0206_
rlabel metal2 5152 25592 5152 25592 0 _0207_
rlabel metal2 6440 24360 6440 24360 0 _0208_
rlabel metal2 4928 24696 4928 24696 0 _0209_
rlabel metal2 4816 23128 4816 23128 0 _0210_
rlabel metal3 5040 20776 5040 20776 0 _0211_
rlabel metal2 6216 65016 6216 65016 0 _0212_
rlabel metal2 5992 65520 5992 65520 0 _0213_
rlabel metal2 35168 64568 35168 64568 0 _0214_
rlabel metal2 33768 58324 33768 58324 0 _0215_
rlabel metal3 34888 63112 34888 63112 0 _0216_
rlabel metal3 34944 64792 34944 64792 0 _0217_
rlabel metal2 33656 65072 33656 65072 0 _0218_
rlabel metal3 32816 60872 32816 60872 0 _0219_
rlabel metal2 33880 60704 33880 60704 0 _0220_
rlabel metal3 32872 65352 32872 65352 0 _0221_
rlabel metal2 34328 66304 34328 66304 0 _0222_
rlabel metal2 32424 65576 32424 65576 0 _0223_
rlabel metal2 33432 69048 33432 69048 0 _0224_
rlabel metal2 35336 66920 35336 66920 0 _0225_
rlabel metal2 35896 65912 35896 65912 0 _0226_
rlabel metal2 35672 63952 35672 63952 0 _0227_
rlabel metal2 33768 55076 33768 55076 0 _0228_
rlabel metal2 33320 54600 33320 54600 0 _0229_
rlabel metal3 33040 55272 33040 55272 0 _0230_
rlabel metal3 34944 63784 34944 63784 0 _0231_
rlabel metal2 36120 64624 36120 64624 0 _0232_
rlabel metal2 35896 67032 35896 67032 0 _0233_
rlabel metal2 32984 67760 32984 67760 0 _0234_
rlabel metal2 33096 68488 33096 68488 0 _0235_
rlabel metal2 32536 66780 32536 66780 0 _0236_
rlabel metal2 33544 61040 33544 61040 0 _0237_
rlabel metal2 32872 60816 32872 60816 0 _0238_
rlabel metal2 32536 60312 32536 60312 0 _0239_
rlabel metal2 31528 61208 31528 61208 0 _0240_
rlabel metal2 33376 60984 33376 60984 0 _0241_
rlabel metal2 32872 64120 32872 64120 0 _0242_
rlabel metal2 33656 67900 33656 67900 0 _0243_
rlabel metal2 33768 69496 33768 69496 0 _0244_
rlabel metal2 33656 70168 33656 70168 0 _0245_
rlabel metal2 34440 68096 34440 68096 0 _0246_
rlabel metal2 36232 67536 36232 67536 0 _0247_
rlabel metal2 36008 70784 36008 70784 0 _0248_
rlabel metal2 36792 64624 36792 64624 0 _0249_
rlabel metal2 36344 68936 36344 68936 0 _0250_
rlabel metal2 37688 70112 37688 70112 0 _0251_
rlabel metal3 36008 52920 36008 52920 0 _0252_
rlabel metal2 38024 52080 38024 52080 0 _0253_
rlabel metal2 35728 56840 35728 56840 0 _0254_
rlabel metal2 33936 54712 33936 54712 0 _0255_
rlabel metal2 34664 54768 34664 54768 0 _0256_
rlabel metal3 34944 55048 34944 55048 0 _0257_
rlabel metal2 35784 50288 35784 50288 0 _0258_
rlabel metal3 33880 49896 33880 49896 0 _0259_
rlabel metal3 33656 50680 33656 50680 0 _0260_
rlabel metal2 35224 50680 35224 50680 0 _0261_
rlabel metal2 35952 55160 35952 55160 0 _0262_
rlabel metal2 36512 56168 36512 56168 0 _0263_
rlabel metal2 37128 69328 37128 69328 0 _0264_
rlabel metal2 34888 71008 34888 71008 0 _0265_
rlabel metal2 32984 70560 32984 70560 0 _0266_
rlabel metal2 33992 71736 33992 71736 0 _0267_
rlabel metal2 32648 71176 32648 71176 0 _0268_
rlabel metal2 33096 72464 33096 72464 0 _0269_
rlabel metal2 31192 72240 31192 72240 0 _0270_
rlabel metal2 30520 70560 30520 70560 0 _0271_
rlabel metal2 38024 69720 38024 69720 0 _0272_
rlabel metal2 38920 70448 38920 70448 0 _0273_
rlabel metal3 36176 71624 36176 71624 0 _0274_
rlabel metal2 38024 54824 38024 54824 0 _0275_
rlabel metal2 35784 56056 35784 56056 0 _0276_
rlabel metal2 37072 55832 37072 55832 0 _0277_
rlabel metal2 38024 56336 38024 56336 0 _0278_
rlabel metal2 35896 49336 35896 49336 0 _0279_
rlabel metal2 36120 48944 36120 48944 0 _0280_
rlabel metal2 37240 48272 37240 48272 0 _0281_
rlabel metal3 34440 47432 34440 47432 0 _0282_
rlabel metal3 33320 47544 33320 47544 0 _0283_
rlabel metal2 34384 47544 34384 47544 0 _0284_
rlabel metal2 34440 48048 34440 48048 0 _0285_
rlabel metal2 37184 47432 37184 47432 0 _0286_
rlabel metal2 38696 48272 38696 48272 0 _0287_
rlabel metal2 33208 41160 33208 41160 0 _0288_
rlabel metal2 35504 41384 35504 41384 0 _0289_
rlabel metal3 36792 41944 36792 41944 0 _0290_
rlabel metal2 37240 41608 37240 41608 0 _0291_
rlabel metal2 38584 46088 38584 46088 0 _0292_
rlabel metal2 38304 53816 38304 53816 0 _0293_
rlabel metal2 39256 55160 39256 55160 0 _0294_
rlabel metal2 39144 70224 39144 70224 0 _0295_
rlabel metal2 30968 70560 30968 70560 0 _0296_
rlabel metal2 31416 72184 31416 72184 0 _0297_
rlabel metal2 30520 72968 30520 72968 0 _0298_
rlabel metal2 30072 71008 30072 71008 0 _0299_
rlabel metal2 30744 71680 30744 71680 0 _0300_
rlabel metal2 29064 70280 29064 70280 0 _0301_
rlabel metal2 37632 50400 37632 50400 0 _0302_
rlabel metal2 38808 54656 38808 54656 0 _0303_
rlabel metal2 38696 54040 38696 54040 0 _0304_
rlabel metal2 39088 41160 39088 41160 0 _0305_
rlabel metal2 32984 41552 32984 41552 0 _0306_
rlabel metal3 34272 41048 34272 41048 0 _0307_
rlabel metal3 36512 40376 36512 40376 0 _0308_
rlabel metal2 37352 40600 37352 40600 0 _0309_
rlabel metal2 37856 40152 37856 40152 0 _0310_
rlabel metal2 37800 20216 37800 20216 0 _0311_
rlabel metal2 38696 22288 38696 22288 0 _0312_
rlabel metal2 39816 29792 39816 29792 0 _0313_
rlabel metal2 37688 48048 37688 48048 0 _0314_
rlabel metal2 37912 44240 37912 44240 0 _0315_
rlabel metal2 35168 46872 35168 46872 0 _0316_
rlabel metal2 34776 45584 34776 45584 0 _0317_
rlabel metal2 31864 44184 31864 44184 0 _0318_
rlabel metal2 30856 45136 30856 45136 0 _0319_
rlabel metal2 30744 45024 30744 45024 0 _0320_
rlabel metal2 31080 45304 31080 45304 0 _0321_
rlabel metal2 34328 44688 34328 44688 0 _0322_
rlabel metal2 35224 45248 35224 45248 0 _0323_
rlabel metal2 34440 41272 34440 41272 0 _0324_
rlabel metal3 35504 40936 35504 40936 0 _0325_
rlabel metal2 35448 40712 35448 40712 0 _0326_
rlabel metal2 35896 40432 35896 40432 0 _0327_
rlabel metal2 36008 39984 36008 39984 0 _0328_
rlabel metal3 36792 44296 36792 44296 0 _0329_
rlabel metal2 38248 44296 38248 44296 0 _0330_
rlabel metal2 39312 44184 39312 44184 0 _0331_
rlabel metal3 39368 38024 39368 38024 0 _0332_
rlabel metal2 29512 66640 29512 66640 0 _0333_
rlabel metal2 35112 71064 35112 71064 0 _0334_
rlabel metal2 30352 64456 30352 64456 0 _0335_
rlabel metal2 29400 69832 29400 69832 0 _0336_
rlabel metal2 28504 70952 28504 70952 0 _0337_
rlabel metal2 30184 66472 30184 66472 0 _0338_
rlabel metal2 29960 69496 29960 69496 0 _0339_
rlabel metal3 30408 67816 30408 67816 0 _0340_
rlabel metal2 29400 63504 29400 63504 0 _0341_
rlabel metal2 38136 34832 38136 34832 0 _0342_
rlabel metal2 40040 36120 40040 36120 0 _0343_
rlabel metal2 38360 37296 38360 37296 0 _0344_
rlabel metal3 39536 36344 39536 36344 0 _0345_
rlabel metal2 38416 32648 38416 32648 0 _0346_
rlabel metal2 38416 43288 38416 43288 0 _0347_
rlabel metal3 36960 32536 36960 32536 0 _0348_
rlabel metal3 36064 45192 36064 45192 0 _0349_
rlabel metal2 36568 45136 36568 45136 0 _0350_
rlabel metal2 35560 31696 35560 31696 0 _0351_
rlabel metal3 31360 44296 31360 44296 0 _0352_
rlabel metal2 30968 44968 30968 44968 0 _0353_
rlabel metal2 31136 40824 31136 40824 0 _0354_
rlabel metal2 29624 37520 29624 37520 0 _0355_
rlabel metal3 27944 45192 27944 45192 0 _0356_
rlabel metal3 28840 37128 28840 37128 0 _0357_
rlabel metal3 32368 37016 32368 37016 0 _0358_
rlabel metal2 33320 34496 33320 34496 0 _0359_
rlabel metal3 33096 39592 33096 39592 0 _0360_
rlabel metal2 33096 41104 33096 41104 0 _0361_
rlabel metal2 33656 39200 33656 39200 0 _0362_
rlabel metal2 33432 36792 33432 36792 0 _0363_
rlabel metal2 35224 34552 35224 34552 0 _0364_
rlabel metal2 35672 32872 35672 32872 0 _0365_
rlabel metal3 36736 31640 36736 31640 0 _0366_
rlabel metal3 35224 30072 35224 30072 0 _0367_
rlabel metal2 36120 27776 36120 27776 0 _0368_
rlabel metal2 36232 39396 36232 39396 0 _0369_
rlabel metal3 36512 19208 36512 19208 0 _0370_
rlabel metal3 36736 19320 36736 19320 0 _0371_
rlabel metal2 35336 19376 35336 19376 0 _0372_
rlabel metal2 36120 25452 36120 25452 0 _0373_
rlabel metal2 36120 30016 36120 30016 0 _0374_
rlabel metal2 37128 33488 37128 33488 0 _0375_
rlabel metal2 31192 62608 31192 62608 0 _0376_
rlabel metal2 30520 65240 30520 65240 0 _0377_
rlabel metal2 29176 69216 29176 69216 0 _0378_
rlabel metal2 29512 61264 29512 61264 0 _0379_
rlabel metal2 29176 62608 29176 62608 0 _0380_
rlabel metal2 30240 63784 30240 63784 0 _0381_
rlabel metal2 38024 34552 38024 34552 0 _0382_
rlabel metal2 32088 32816 32088 32816 0 _0383_
rlabel metal3 36624 30184 36624 30184 0 _0384_
rlabel metal2 33320 31192 33320 31192 0 _0385_
rlabel metal2 35560 28000 35560 28000 0 _0386_
rlabel metal2 36232 27720 36232 27720 0 _0387_
rlabel metal2 32760 27832 32760 27832 0 _0388_
rlabel metal3 35112 30184 35112 30184 0 _0389_
rlabel metal2 33824 28504 33824 28504 0 _0390_
rlabel metal2 31304 37072 31304 37072 0 _0391_
rlabel metal2 31080 35280 31080 35280 0 _0392_
rlabel metal2 32312 36008 32312 36008 0 _0393_
rlabel metal2 32424 25368 32424 25368 0 _0394_
rlabel metal3 29232 35784 29232 35784 0 _0395_
rlabel metal2 30408 39816 30408 39816 0 _0396_
rlabel metal2 29960 36848 29960 36848 0 _0397_
rlabel metal2 30520 35896 30520 35896 0 _0398_
rlabel metal2 30520 38668 30520 38668 0 _0399_
rlabel metal2 31360 35560 31360 35560 0 _0400_
rlabel metal2 33880 35560 33880 35560 0 _0401_
rlabel metal2 34888 33208 34888 33208 0 _0402_
rlabel metal2 34104 26236 34104 26236 0 _0403_
rlabel metal2 31864 24808 31864 24808 0 _0404_
rlabel metal2 32312 25200 32312 25200 0 _0405_
rlabel metal2 33040 23912 33040 23912 0 _0406_
rlabel metal2 33992 24192 33992 24192 0 _0407_
rlabel metal2 36456 20160 36456 20160 0 _0408_
rlabel metal2 36120 19320 36120 19320 0 _0409_
rlabel metal2 37576 19488 37576 19488 0 _0410_
rlabel metal2 35112 19656 35112 19656 0 _0411_
rlabel metal2 33208 39872 33208 39872 0 _0412_
rlabel metal2 35224 20160 35224 20160 0 _0413_
rlabel metal2 35168 14728 35168 14728 0 _0414_
rlabel metal2 35560 14336 35560 14336 0 _0415_
rlabel metal2 34776 14112 34776 14112 0 _0416_
rlabel metal2 34048 14280 34048 14280 0 _0417_
rlabel metal2 33656 22400 33656 22400 0 _0418_
rlabel metal2 31640 30184 31640 30184 0 _0419_
rlabel metal3 30352 31752 30352 31752 0 _0420_
rlabel metal3 31584 62328 31584 62328 0 _0421_
rlabel metal2 31528 63448 31528 63448 0 _0422_
rlabel metal2 30968 63504 30968 63504 0 _0423_
rlabel metal2 25928 75432 25928 75432 0 _0424_
rlabel metal2 28504 30912 28504 30912 0 _0425_
rlabel metal2 28840 31080 28840 31080 0 _0426_
rlabel metal2 29288 30128 29288 30128 0 _0427_
rlabel metal2 15288 43792 15288 43792 0 _0428_
rlabel metal2 32536 29848 32536 29848 0 _0429_
rlabel metal2 28056 28840 28056 28840 0 _0430_
rlabel metal3 33376 27048 33376 27048 0 _0431_
rlabel metal2 33208 28448 33208 28448 0 _0432_
rlabel metal2 33096 28168 33096 28168 0 _0433_
rlabel metal2 30912 26488 30912 26488 0 _0434_
rlabel metal2 33992 19264 33992 19264 0 _0435_
rlabel metal2 33432 18928 33432 18928 0 _0436_
rlabel metal2 33040 20776 33040 20776 0 _0437_
rlabel metal2 32816 24696 32816 24696 0 _0438_
rlabel metal3 33208 20888 33208 20888 0 _0439_
rlabel metal2 31136 14616 31136 14616 0 _0440_
rlabel metal2 32312 11424 32312 11424 0 _0441_
rlabel metal2 30184 14840 30184 14840 0 _0442_
rlabel metal2 31864 12544 31864 12544 0 _0443_
rlabel metal2 31192 16464 31192 16464 0 _0444_
rlabel metal2 31976 18704 31976 18704 0 _0445_
rlabel metal2 32592 19320 32592 19320 0 _0446_
rlabel metal2 31864 16072 31864 16072 0 _0447_
rlabel metal2 31640 12600 31640 12600 0 _0448_
rlabel metal2 32872 12096 32872 12096 0 _0449_
rlabel metal3 33376 11368 33376 11368 0 _0450_
rlabel metal2 35000 13664 35000 13664 0 _0451_
rlabel metal2 35336 12992 35336 12992 0 _0452_
rlabel metal3 35336 10696 35336 10696 0 _0453_
rlabel metal2 34440 33656 34440 33656 0 _0454_
rlabel metal2 34776 33656 34776 33656 0 _0455_
rlabel metal2 34328 8232 34328 8232 0 _0456_
rlabel metal2 35896 4368 35896 4368 0 _0457_
rlabel metal2 36904 6272 36904 6272 0 _0458_
rlabel metal2 35336 6216 35336 6216 0 _0459_
rlabel metal2 35560 6776 35560 6776 0 _0460_
rlabel metal2 34216 11088 34216 11088 0 _0461_
rlabel metal2 33376 11256 33376 11256 0 _0462_
rlabel metal2 31472 26376 31472 26376 0 _0463_
rlabel metal2 29736 28672 29736 28672 0 _0464_
rlabel metal3 28952 30072 28952 30072 0 _0465_
rlabel metal2 28504 72520 28504 72520 0 _0466_
rlabel metal2 27552 27944 27552 27944 0 _0467_
rlabel metal2 28728 29288 28728 29288 0 _0468_
rlabel metal2 25480 28728 25480 28728 0 _0469_
rlabel metal2 31080 26824 31080 26824 0 _0470_
rlabel metal2 31864 26768 31864 26768 0 _0471_
rlabel metal2 29848 23632 29848 23632 0 _0472_
rlabel metal2 31360 20216 31360 20216 0 _0473_
rlabel metal2 32088 20048 32088 20048 0 _0474_
rlabel metal2 30184 20496 30184 20496 0 _0475_
rlabel metal2 35000 6272 35000 6272 0 _0476_
rlabel metal3 34832 8456 34832 8456 0 _0477_
rlabel metal2 34664 9128 34664 9128 0 _0478_
rlabel metal2 34832 8232 34832 8232 0 _0479_
rlabel metal2 33432 7840 33432 7840 0 _0480_
rlabel metal2 32928 10696 32928 10696 0 _0481_
rlabel metal2 33320 10864 33320 10864 0 _0482_
rlabel metal2 33880 6664 33880 6664 0 _0483_
rlabel metal2 36008 5544 36008 5544 0 _0484_
rlabel metal2 29848 6384 29848 6384 0 _0485_
rlabel metal2 29792 16744 29792 16744 0 _0486_
rlabel metal2 30072 4816 30072 4816 0 _0487_
rlabel metal2 25704 11816 25704 11816 0 _0488_
rlabel metal2 26040 10920 26040 10920 0 _0489_
rlabel metal2 27048 6356 27048 6356 0 _0490_
rlabel metal3 29064 4312 29064 4312 0 _0491_
rlabel metal2 31976 6720 31976 6720 0 _0492_
rlabel metal2 31360 12376 31360 12376 0 _0493_
rlabel metal2 31528 8316 31528 8316 0 _0494_
rlabel metal2 30408 17136 30408 17136 0 _0495_
rlabel metal2 30184 13888 30184 13888 0 _0496_
rlabel metal2 31864 10584 31864 10584 0 _0497_
rlabel metal3 31472 9128 31472 9128 0 _0498_
rlabel metal2 32200 6608 32200 6608 0 _0499_
rlabel metal3 33432 6664 33432 6664 0 _0500_
rlabel metal2 31808 6664 31808 6664 0 _0501_
rlabel metal2 29736 23632 29736 23632 0 _0502_
rlabel metal2 25480 25088 25480 25088 0 _0503_
rlabel metal2 25312 24808 25312 24808 0 _0504_
rlabel metal2 20832 73976 20832 73976 0 _0505_
rlabel metal2 25816 26292 25816 26292 0 _0506_
rlabel metal2 25928 28672 25928 28672 0 _0507_
rlabel metal2 30464 19992 30464 19992 0 _0508_
rlabel metal2 29960 20608 29960 20608 0 _0509_
rlabel metal2 30632 22400 30632 22400 0 _0510_
rlabel metal3 30016 21560 30016 21560 0 _0511_
rlabel metal2 34552 7112 34552 7112 0 _0512_
rlabel metal2 31640 7056 31640 7056 0 _0513_
rlabel metal2 28504 9856 28504 9856 0 _0514_
rlabel metal2 26712 11760 26712 11760 0 _0515_
rlabel metal2 26824 10976 26824 10976 0 _0516_
rlabel metal2 27384 10360 27384 10360 0 _0517_
rlabel metal2 26992 10808 26992 10808 0 _0518_
rlabel metal2 27776 11368 27776 11368 0 _0519_
rlabel metal2 30744 9856 30744 9856 0 _0520_
rlabel metal2 31864 8344 31864 8344 0 _0521_
rlabel metal2 31304 9576 31304 9576 0 _0522_
rlabel metal2 29960 4704 29960 4704 0 _0523_
rlabel metal2 29568 5208 29568 5208 0 _0524_
rlabel metal2 30128 4088 30128 4088 0 _0525_
rlabel metal2 29288 6272 29288 6272 0 _0526_
rlabel metal2 29792 12936 29792 12936 0 _0527_
rlabel metal2 29400 13272 29400 13272 0 _0528_
rlabel metal2 29960 7140 29960 7140 0 _0529_
rlabel metal2 30296 6608 30296 6608 0 _0530_
rlabel metal2 29568 9576 29568 9576 0 _0531_
rlabel metal2 29848 15848 29848 15848 0 _0532_
rlabel metal2 29064 23296 29064 23296 0 _0533_
rlabel metal2 25592 30240 25592 30240 0 _0534_
rlabel metal2 33264 72632 33264 72632 0 _0535_
rlabel metal2 19040 20664 19040 20664 0 _0536_
rlabel metal2 19208 41496 19208 41496 0 _0537_
rlabel metal2 2184 33712 2184 33712 0 _0538_
rlabel metal2 2744 32032 2744 32032 0 _0539_
rlabel metal2 15176 46648 15176 46648 0 _0540_
rlabel metal2 2968 49728 2968 49728 0 _0541_
rlabel metal2 2744 32760 2744 32760 0 _0542_
rlabel metal2 20496 42728 20496 42728 0 _0543_
rlabel metal3 17612 42616 17612 42616 0 _0544_
rlabel metal2 10304 43624 10304 43624 0 _0545_
rlabel metal3 9912 57792 9912 57792 0 _0546_
rlabel metal2 20328 43904 20328 43904 0 _0547_
rlabel metal2 18536 47936 18536 47936 0 _0548_
rlabel metal2 9408 57624 9408 57624 0 _0549_
rlabel metal2 15176 45472 15176 45472 0 _0550_
rlabel metal2 15960 46368 15960 46368 0 _0551_
rlabel metal2 9744 56840 9744 56840 0 _0552_
rlabel metal2 9240 57512 9240 57512 0 _0553_
rlabel metal2 2184 49056 2184 49056 0 _0554_
rlabel metal2 2240 47656 2240 47656 0 _0555_
rlabel metal2 2576 49784 2576 49784 0 _0556_
rlabel metal3 10136 52920 10136 52920 0 _0557_
rlabel metal2 9352 53032 9352 53032 0 _0558_
rlabel metal2 2576 47656 2576 47656 0 _0559_
rlabel metal2 11648 46872 11648 46872 0 _0560_
rlabel metal2 2744 47628 2744 47628 0 _0561_
rlabel metal2 2632 43792 2632 43792 0 _0562_
rlabel metal2 2800 44520 2800 44520 0 _0563_
rlabel metal2 9912 43120 9912 43120 0 _0564_
rlabel metal2 19544 50904 19544 50904 0 _0565_
rlabel metal2 19208 52472 19208 52472 0 _0566_
rlabel metal2 9632 64904 9632 64904 0 _0567_
rlabel metal2 11816 41776 11816 41776 0 _0568_
rlabel metal2 16856 44240 16856 44240 0 _0569_
rlabel metal2 11704 43120 11704 43120 0 _0570_
rlabel metal3 11592 45752 11592 45752 0 _0571_
rlabel metal2 11312 43512 11312 43512 0 _0572_
rlabel metal2 11088 42952 11088 42952 0 _0573_
rlabel metal2 17080 45416 17080 45416 0 _0574_
rlabel metal2 15848 46144 15848 46144 0 _0575_
rlabel metal3 16632 45080 16632 45080 0 _0576_
rlabel metal2 15400 45584 15400 45584 0 _0577_
rlabel metal2 15960 43568 15960 43568 0 _0578_
rlabel metal2 16352 43624 16352 43624 0 _0579_
rlabel metal2 15400 48860 15400 48860 0 _0580_
rlabel metal2 15568 43624 15568 43624 0 _0581_
rlabel metal2 12376 43792 12376 43792 0 _0582_
rlabel metal2 14168 43960 14168 43960 0 _0583_
rlabel metal2 14168 46928 14168 46928 0 _0584_
rlabel metal2 16968 39704 16968 39704 0 _0585_
rlabel metal2 15848 41048 15848 41048 0 _0586_
rlabel metal2 16968 40880 16968 40880 0 _0587_
rlabel metal2 16744 41552 16744 41552 0 _0588_
rlabel metal2 17920 45864 17920 45864 0 _0589_
rlabel metal2 17584 46088 17584 46088 0 _0590_
rlabel metal3 13552 61544 13552 61544 0 _0591_
rlabel metal2 13720 61488 13720 61488 0 _0592_
rlabel metal2 16968 60256 16968 60256 0 _0593_
rlabel metal2 11536 63896 11536 63896 0 _0594_
rlabel metal2 13496 61320 13496 61320 0 _0595_
rlabel metal2 12040 64792 12040 64792 0 _0596_
rlabel metal2 11032 64792 11032 64792 0 _0597_
rlabel metal2 15624 63112 15624 63112 0 _0598_
rlabel metal2 12488 66024 12488 66024 0 _0599_
rlabel metal2 12096 64120 12096 64120 0 _0600_
rlabel metal3 12096 64568 12096 64568 0 _0601_
rlabel metal2 10584 64344 10584 64344 0 _0602_
rlabel metal2 22680 60648 22680 60648 0 _0603_
rlabel metal3 17360 62328 17360 62328 0 _0604_
rlabel metal2 18648 61320 18648 61320 0 _0605_
rlabel metal2 17136 62328 17136 62328 0 _0606_
rlabel metal2 22792 60144 22792 60144 0 _0607_
rlabel metal3 21000 59976 21000 59976 0 _0608_
rlabel metal3 21448 59864 21448 59864 0 _0609_
rlabel metal2 22792 61712 22792 61712 0 _0610_
rlabel metal2 21672 61488 21672 61488 0 _0611_
rlabel metal2 20216 60648 20216 60648 0 _0612_
rlabel metal3 19432 59976 19432 59976 0 _0613_
rlabel metal2 23912 53032 23912 53032 0 _0614_
rlabel metal2 24416 54600 24416 54600 0 _0615_
rlabel metal2 25312 59416 25312 59416 0 _0616_
rlabel metal2 22456 53704 22456 53704 0 _0617_
rlabel metal2 24024 58408 24024 58408 0 _0618_
rlabel metal2 24248 59696 24248 59696 0 _0619_
rlabel metal2 26264 58520 26264 58520 0 _0620_
rlabel metal2 25816 58352 25816 58352 0 _0621_
rlabel metal2 26376 58296 26376 58296 0 _0622_
rlabel metal2 24808 53592 24808 53592 0 _0623_
rlabel metal2 26152 54880 26152 54880 0 _0624_
rlabel metal2 26040 54376 26040 54376 0 _0625_
rlabel metal2 25536 54488 25536 54488 0 _0626_
rlabel metal2 24696 47936 24696 47936 0 _0627_
rlabel metal2 26096 53032 26096 53032 0 _0628_
rlabel metal2 23576 41216 23576 41216 0 _0629_
rlabel metal2 21896 52752 21896 52752 0 _0630_
rlabel metal2 24360 47824 24360 47824 0 _0631_
rlabel metal3 23688 47208 23688 47208 0 _0632_
rlabel metal2 16632 45808 16632 45808 0 _0633_
rlabel metal2 24696 38864 24696 38864 0 _0634_
rlabel metal2 25592 38864 25592 38864 0 _0635_
rlabel metal2 25256 39536 25256 39536 0 _0636_
rlabel metal2 24920 38304 24920 38304 0 _0637_
rlabel metal3 23184 38808 23184 38808 0 _0638_
rlabel metal2 13944 65800 13944 65800 0 _0639_
rlabel metal2 18424 62944 18424 62944 0 _0640_
rlabel metal2 15288 66640 15288 66640 0 _0641_
rlabel metal2 16296 64904 16296 64904 0 _0642_
rlabel metal2 13832 64512 13832 64512 0 _0643_
rlabel metal2 14168 66640 14168 66640 0 _0644_
rlabel metal2 14280 65072 14280 65072 0 _0645_
rlabel metal3 16408 65296 16408 65296 0 _0646_
rlabel metal2 17640 64904 17640 64904 0 _0647_
rlabel metal3 17864 64568 17864 64568 0 _0648_
rlabel metal2 19992 63392 19992 63392 0 _0649_
rlabel metal2 17752 64064 17752 64064 0 _0650_
rlabel metal3 21000 63224 21000 63224 0 _0651_
rlabel metal2 20440 65072 20440 65072 0 _0652_
rlabel metal2 18872 63616 18872 63616 0 _0653_
rlabel metal2 22792 44072 22792 44072 0 _0654_
rlabel metal2 26040 45024 26040 45024 0 _0655_
rlabel metal2 25424 47432 25424 47432 0 _0656_
rlabel metal2 20328 47824 20328 47824 0 _0657_
rlabel metal2 22120 44352 22120 44352 0 _0658_
rlabel metal3 23632 46760 23632 46760 0 _0659_
rlabel metal2 23408 46872 23408 46872 0 _0660_
rlabel metal2 25592 46536 25592 46536 0 _0661_
rlabel metal3 24864 46648 24864 46648 0 _0662_
rlabel metal2 25872 41944 25872 41944 0 _0663_
rlabel metal2 25480 45080 25480 45080 0 _0664_
rlabel metal2 24472 42056 24472 42056 0 _0665_
rlabel metal2 27048 43232 27048 43232 0 _0666_
rlabel metal2 25200 43512 25200 43512 0 _0667_
rlabel metal2 24808 41272 24808 41272 0 _0668_
rlabel metal3 24752 41944 24752 41944 0 _0669_
rlabel metal3 24136 44520 24136 44520 0 _0670_
rlabel metal2 23912 39648 23912 39648 0 _0671_
rlabel metal3 24360 40488 24360 40488 0 _0672_
rlabel metal2 23128 39872 23128 39872 0 _0673_
rlabel metal2 21616 40152 21616 40152 0 _0674_
rlabel metal2 22008 40488 22008 40488 0 _0675_
rlabel metal3 17696 49784 17696 49784 0 _0676_
rlabel metal2 16072 56000 16072 56000 0 _0677_
rlabel metal2 15064 49280 15064 49280 0 _0678_
rlabel metal2 13608 48664 13608 48664 0 _0679_
rlabel metal3 13720 54600 13720 54600 0 _0680_
rlabel metal2 14616 48888 14616 48888 0 _0681_
rlabel metal3 16184 52920 16184 52920 0 _0682_
rlabel metal3 14896 52920 14896 52920 0 _0683_
rlabel metal2 15288 54040 15288 54040 0 _0684_
rlabel metal3 14056 53704 14056 53704 0 _0685_
rlabel metal2 14616 57344 14616 57344 0 _0686_
rlabel metal2 14168 56952 14168 56952 0 _0687_
rlabel metal2 14392 47432 14392 47432 0 _0688_
rlabel metal2 13720 56000 13720 56000 0 _0689_
rlabel metal3 12880 56728 12880 56728 0 _0690_
rlabel metal2 11480 55048 11480 55048 0 _0691_
rlabel metal2 11928 56728 11928 56728 0 _0692_
rlabel metal2 12152 55048 12152 55048 0 _0693_
rlabel metal2 11816 55328 11816 55328 0 _0694_
rlabel metal3 12992 52136 12992 52136 0 _0695_
rlabel metal2 12264 52528 12264 52528 0 _0696_
rlabel metal2 11088 48328 11088 48328 0 _0697_
rlabel metal2 10808 48216 10808 48216 0 _0698_
rlabel metal2 14224 4312 14224 4312 0 _0699_
rlabel metal2 6104 69664 6104 69664 0 _0700_
rlabel metal3 17192 49000 17192 49000 0 _0701_
rlabel metal2 22344 69720 22344 69720 0 _0702_
rlabel metal2 22624 69608 22624 69608 0 _0703_
rlabel metal2 22792 70056 22792 70056 0 _0704_
rlabel metal2 23408 68712 23408 68712 0 _0705_
rlabel metal2 23464 69776 23464 69776 0 _0706_
rlabel metal2 18424 70448 18424 70448 0 _0707_
rlabel metal2 19712 70280 19712 70280 0 _0708_
rlabel metal2 19936 71176 19936 71176 0 _0709_
rlabel metal2 19936 70952 19936 70952 0 _0710_
rlabel metal2 8232 70224 8232 70224 0 _0711_
rlabel metal3 8064 48440 8064 48440 0 _0712_
rlabel metal3 8848 45080 8848 45080 0 _0713_
rlabel metal2 23576 71232 23576 71232 0 _0714_
rlabel metal2 22624 73192 22624 73192 0 _0715_
rlabel metal2 24584 70616 24584 70616 0 _0716_
rlabel metal2 25088 72408 25088 72408 0 _0717_
rlabel metal3 23128 71120 23128 71120 0 _0718_
rlabel metal2 18872 71064 18872 71064 0 _0719_
rlabel metal2 19432 72128 19432 72128 0 _0720_
rlabel metal2 21336 72464 21336 72464 0 _0721_
rlabel metal3 19824 72856 19824 72856 0 _0722_
rlabel metal2 18536 71176 18536 71176 0 _0723_
rlabel metal2 1512 54656 1512 54656 0 _0724_
rlabel metal2 8344 45136 8344 45136 0 _0725_
rlabel metal2 7224 40880 7224 40880 0 _0726_
rlabel metal2 7504 22344 7504 22344 0 _0727_
rlabel metal2 5768 44744 5768 44744 0 _0728_
rlabel metal2 1400 46816 1400 46816 0 _0729_
rlabel metal2 8736 70280 8736 70280 0 _0730_
rlabel metal2 9016 70504 9016 70504 0 _0731_
rlabel metal2 8680 69496 8680 69496 0 _0732_
rlabel metal2 10920 22512 10920 22512 0 _0733_
rlabel metal3 20216 42336 20216 42336 0 _0734_
rlabel metal2 22232 49392 22232 49392 0 _0735_
rlabel metal2 20664 45528 20664 45528 0 _0736_
rlabel metal3 23492 49784 23492 49784 0 _0737_
rlabel metal2 25760 50008 25760 50008 0 _0738_
rlabel metal2 25816 50792 25816 50792 0 _0739_
rlabel metal2 41160 48608 41160 48608 0 _0740_
rlabel metal2 39984 41944 39984 41944 0 _0741_
rlabel metal2 38808 60816 38808 60816 0 _0742_
rlabel metal2 25592 59472 25592 59472 0 _0743_
rlabel metal2 21560 45864 21560 45864 0 _0744_
rlabel metal2 21448 52080 21448 52080 0 _0745_
rlabel metal2 25368 51352 25368 51352 0 _0746_
rlabel metal2 26488 49448 26488 49448 0 _0747_
rlabel metal2 25984 57848 25984 57848 0 _0748_
rlabel metal2 32816 52136 32816 52136 0 _0749_
rlabel metal3 32144 52024 32144 52024 0 _0750_
rlabel metal3 30128 55384 30128 55384 0 _0751_
rlabel metal2 19880 52528 19880 52528 0 _0752_
rlabel metal2 20104 50792 20104 50792 0 _0753_
rlabel metal2 21000 42504 21000 42504 0 _0754_
rlabel metal2 20944 50344 20944 50344 0 _0755_
rlabel metal2 23240 47544 23240 47544 0 _0756_
rlabel metal2 23576 56112 23576 56112 0 _0757_
rlabel metal2 26040 56504 26040 56504 0 _0758_
rlabel metal2 10808 24304 10808 24304 0 _0759_
rlabel metal2 10584 19208 10584 19208 0 _0760_
rlabel metal2 29120 70728 29120 70728 0 _0761_
rlabel metal2 40936 41888 40936 41888 0 _0762_
rlabel metal3 39368 41160 39368 41160 0 _0763_
rlabel metal2 26936 57792 26936 57792 0 _0764_
rlabel metal2 27720 56336 27720 56336 0 _0765_
rlabel metal2 33544 54824 33544 54824 0 _0766_
rlabel metal2 35560 49336 35560 49336 0 _0767_
rlabel metal2 26264 47208 26264 47208 0 _0768_
rlabel metal2 22680 58016 22680 58016 0 _0769_
rlabel metal2 26488 56392 26488 56392 0 _0770_
rlabel metal3 32648 47320 32648 47320 0 _0771_
rlabel metal2 30408 45696 30408 45696 0 _0772_
rlabel metal2 20440 51744 20440 51744 0 _0773_
rlabel metal2 41496 41160 41496 41160 0 _0774_
rlabel metal2 41832 39480 41832 39480 0 _0775_
rlabel metal2 24640 53032 24640 53032 0 _0776_
rlabel metal2 23464 52304 23464 52304 0 _0777_
rlabel metal2 26936 51632 26936 51632 0 _0778_
rlabel metal2 12376 13832 12376 13832 0 _0779_
rlabel metal2 13272 11872 13272 11872 0 _0780_
rlabel metal2 26376 19320 26376 19320 0 _0781_
rlabel metal2 30744 67396 30744 67396 0 _0782_
rlabel metal3 28560 50456 28560 50456 0 _0783_
rlabel metal2 30632 40488 30632 40488 0 _0784_
rlabel metal2 27048 42672 27048 42672 0 _0785_
rlabel metal2 41720 39872 41720 39872 0 _0786_
rlabel metal2 41608 23408 41608 23408 0 _0787_
rlabel metal2 23464 50960 23464 50960 0 _0788_
rlabel metal3 28784 50344 28784 50344 0 _0789_
rlabel metal2 15736 37184 15736 37184 0 _0790_
rlabel metal2 28952 63392 28952 63392 0 _0791_
rlabel metal2 28448 62888 28448 62888 0 _0792_
rlabel metal2 26264 50400 26264 50400 0 _0793_
rlabel metal2 14840 25648 14840 25648 0 _0794_
rlabel metal2 14056 12600 14056 12600 0 _0795_
rlabel metal2 14952 13496 14952 13496 0 _0796_
rlabel metal3 26152 47152 26152 47152 0 _0797_
rlabel metal2 41160 32536 41160 32536 0 _0798_
rlabel metal3 26376 49896 26376 49896 0 _0799_
rlabel metal2 26824 49000 26824 49000 0 _0800_
rlabel metal2 34944 40600 34944 40600 0 _0801_
rlabel metal2 26824 44296 26824 44296 0 _0802_
rlabel metal2 26488 48552 26488 48552 0 _0803_
rlabel metal2 17304 21280 17304 21280 0 _0804_
rlabel metal2 25928 22512 25928 22512 0 _0805_
rlabel metal2 18088 44632 18088 44632 0 _0806_
rlabel metal2 18144 46872 18144 46872 0 _0807_
rlabel metal3 19376 33544 19376 33544 0 _0808_
rlabel metal2 19992 33824 19992 33824 0 _0809_
rlabel metal3 40824 32648 40824 32648 0 _0810_
rlabel metal2 25704 42504 25704 42504 0 _0811_
rlabel metal2 31696 17752 31696 17752 0 _0812_
rlabel metal3 30856 17416 30856 17416 0 _0813_
rlabel metal2 25088 24024 25088 24024 0 _0814_
rlabel metal2 23688 41440 23688 41440 0 _0815_
rlabel metal2 22288 41832 22288 41832 0 _0816_
rlabel metal2 24136 42280 24136 42280 0 _0817_
rlabel metal2 25368 40600 25368 40600 0 _0818_
rlabel metal2 18536 20944 18536 20944 0 _0819_
rlabel metal2 21672 17640 21672 17640 0 _0820_
rlabel metal2 24360 15680 24360 15680 0 _0821_
rlabel metal2 25816 21168 25816 21168 0 _0822_
rlabel metal3 37800 11368 37800 11368 0 _0823_
rlabel metal2 27608 10248 27608 10248 0 _0824_
rlabel metal2 29120 14504 29120 14504 0 _0825_
rlabel metal3 29344 14616 29344 14616 0 _0826_
rlabel metal2 22680 36624 22680 36624 0 _0827_
rlabel via2 21336 45752 21336 45752 0 _0828_
rlabel metal2 22456 48860 22456 48860 0 _0829_
rlabel metal2 47096 16408 47096 16408 0 _0830_
rlabel metal2 20888 25032 20888 25032 0 _0831_
rlabel metal2 22904 19992 22904 19992 0 _0832_
rlabel metal3 24584 20104 24584 20104 0 _0833_
rlabel metal2 27608 13496 27608 13496 0 _0834_
rlabel metal2 26488 19432 26488 19432 0 _0835_
rlabel metal2 47152 19880 47152 19880 0 _0836_
rlabel metal2 2520 31696 2520 31696 0 _0837_
rlabel metal3 21168 29624 21168 29624 0 _0838_
rlabel metal2 19432 27216 19432 27216 0 _0839_
rlabel metal2 18424 49168 18424 49168 0 _0840_
rlabel metal3 17472 54600 17472 54600 0 _0841_
rlabel metal2 24584 55888 24584 55888 0 _0842_
rlabel metal2 20104 57008 20104 57008 0 _0843_
rlabel metal2 18648 54264 18648 54264 0 _0844_
rlabel metal2 18480 54488 18480 54488 0 _0845_
rlabel metal3 19656 55832 19656 55832 0 _0846_
rlabel metal2 19376 57176 19376 57176 0 _0847_
rlabel metal2 17864 53816 17864 53816 0 _0848_
rlabel metal2 17528 55496 17528 55496 0 _0849_
rlabel metal2 18648 56336 18648 56336 0 _0850_
rlabel metal2 17248 72296 17248 72296 0 _0851_
rlabel metal3 17304 59304 17304 59304 0 _0852_
rlabel metal2 18200 58520 18200 58520 0 _0853_
rlabel metal2 19208 56840 19208 56840 0 _0854_
rlabel metal2 17528 57064 17528 57064 0 _0855_
rlabel metal2 19880 57176 19880 57176 0 _0856_
rlabel metal2 18872 57680 18872 57680 0 _0857_
rlabel metal3 23240 64568 23240 64568 0 _0858_
rlabel metal2 18200 55440 18200 55440 0 _0859_
rlabel metal2 22120 56504 22120 56504 0 _0860_
rlabel metal2 23016 65856 23016 65856 0 _0861_
rlabel metal2 21000 53368 21000 53368 0 _0862_
rlabel metal2 22568 55720 22568 55720 0 _0863_
rlabel metal2 19544 64512 19544 64512 0 _0864_
rlabel metal2 20832 51576 20832 51576 0 _0865_
rlabel metal3 21112 57624 21112 57624 0 _0866_
rlabel metal4 12600 25424 12600 25424 0 _0867_
rlabel metal2 18536 34776 18536 34776 0 _0868_
rlabel metal2 42112 49112 42112 49112 0 _0869_
rlabel metal2 7616 68488 7616 68488 0 _0870_
rlabel metal2 8288 47096 8288 47096 0 _0871_
rlabel metal2 7168 56280 7168 56280 0 _0872_
rlabel metal2 8512 40488 8512 40488 0 _0873_
rlabel metal2 8456 38416 8456 38416 0 _0874_
rlabel metal3 8008 42952 8008 42952 0 _0875_
rlabel metal2 2408 43932 2408 43932 0 _0876_
rlabel metal2 10584 39816 10584 39816 0 _0877_
rlabel metal2 8008 35672 8008 35672 0 _0878_
rlabel metal3 3248 49784 3248 49784 0 _0879_
rlabel metal2 7336 52416 7336 52416 0 _0880_
rlabel metal2 11088 52248 11088 52248 0 _0881_
rlabel metal2 10248 53256 10248 53256 0 _0882_
rlabel metal2 4200 45752 4200 45752 0 _0883_
rlabel metal2 4984 48664 4984 48664 0 _0884_
rlabel metal2 6888 53480 6888 53480 0 _0885_
rlabel metal2 8904 51632 8904 51632 0 _0886_
rlabel metal2 8008 47992 8008 47992 0 _0887_
rlabel metal2 5656 50624 5656 50624 0 _0888_
rlabel metal2 6104 52304 6104 52304 0 _0889_
rlabel metal2 7672 48216 7672 48216 0 _0890_
rlabel metal2 6440 49364 6440 49364 0 _0891_
rlabel metal2 8232 47824 8232 47824 0 _0892_
rlabel metal2 7504 48888 7504 48888 0 _0893_
rlabel metal2 7280 39592 7280 39592 0 _0894_
rlabel metal2 9128 43064 9128 43064 0 _0895_
rlabel metal2 6608 42952 6608 42952 0 _0896_
rlabel metal3 7896 39480 7896 39480 0 _0897_
rlabel metal2 8344 36792 8344 36792 0 _0898_
rlabel metal2 5880 43568 5880 43568 0 _0899_
rlabel metal2 6888 43848 6888 43848 0 _0900_
rlabel metal2 7784 37856 7784 37856 0 _0901_
rlabel metal2 8456 35896 8456 35896 0 _0902_
rlabel metal2 8680 34440 8680 34440 0 _0903_
rlabel metal2 18312 21728 18312 21728 0 _0904_
rlabel metal2 20440 39004 20440 39004 0 _0905_
rlabel metal2 33096 48776 33096 48776 0 _0906_
rlabel metal2 31304 58072 31304 58072 0 _0907_
rlabel metal2 16072 33936 16072 33936 0 _0908_
rlabel metal2 21392 39368 21392 39368 0 _0909_
rlabel metal3 30184 71848 30184 71848 0 _0910_
rlabel metal2 16968 25872 16968 25872 0 _0911_
rlabel metal3 17920 21560 17920 21560 0 _0912_
rlabel metal2 20888 24864 20888 24864 0 _0913_
rlabel metal2 31248 57512 31248 57512 0 _0914_
rlabel metal2 30184 57512 30184 57512 0 _0915_
rlabel metal3 17472 21336 17472 21336 0 _0916_
rlabel metal3 9128 40936 9128 40936 0 _0917_
rlabel metal2 7784 32648 7784 32648 0 _0918_
rlabel metal2 11032 47320 11032 47320 0 _0919_
rlabel metal2 7448 32648 7448 32648 0 _0920_
rlabel metal2 6552 33656 6552 33656 0 _0921_
rlabel metal3 5152 34888 5152 34888 0 _0922_
rlabel metal3 8960 30968 8960 30968 0 _0923_
rlabel metal3 8792 33208 8792 33208 0 _0924_
rlabel metal2 10584 29400 10584 29400 0 _0925_
rlabel metal3 11508 29512 11508 29512 0 _0926_
rlabel metal2 16744 22960 16744 22960 0 _0927_
rlabel metal2 17752 35952 17752 35952 0 _0928_
rlabel metal2 18312 37744 18312 37744 0 _0929_
rlabel metal2 19768 36904 19768 36904 0 _0930_
rlabel metal2 28672 45640 28672 45640 0 _0931_
rlabel via2 32088 66248 32088 66248 0 _0932_
rlabel metal2 34440 66192 34440 66192 0 _0933_
rlabel metal2 32200 52864 32200 52864 0 _0934_
rlabel metal2 22568 20384 22568 20384 0 _0935_
rlabel metal3 41328 60760 41328 60760 0 _0936_
rlabel metal3 39480 57624 39480 57624 0 _0937_
rlabel metal2 39480 61096 39480 61096 0 _0938_
rlabel metal2 40376 43904 40376 43904 0 _0939_
rlabel metal2 38808 47152 38808 47152 0 _0940_
rlabel metal2 41608 40768 41608 40768 0 _0941_
rlabel metal2 39816 60256 39816 60256 0 _0942_
rlabel metal2 38696 63896 38696 63896 0 _0943_
rlabel metal2 38808 44072 38808 44072 0 _0944_
rlabel metal2 38920 59528 38920 59528 0 _0945_
rlabel metal2 37856 59416 37856 59416 0 _0946_
rlabel metal2 22008 19376 22008 19376 0 _0947_
rlabel metal2 38024 24920 38024 24920 0 _0948_
rlabel metal2 36344 60816 36344 60816 0 _0949_
rlabel metal2 37408 61544 37408 61544 0 _0950_
rlabel metal2 37912 63840 37912 63840 0 _0951_
rlabel metal2 36624 14616 36624 14616 0 _0952_
rlabel metal2 38192 63672 38192 63672 0 _0953_
rlabel metal2 38360 64120 38360 64120 0 _0954_
rlabel metal2 38696 65128 38696 65128 0 _0955_
rlabel metal2 39200 65688 39200 65688 0 _0956_
rlabel metal2 39480 66360 39480 66360 0 _0957_
rlabel metal2 29008 46760 29008 46760 0 _0958_
rlabel metal2 20888 37128 20888 37128 0 _0959_
rlabel metal3 18480 35560 18480 35560 0 _0960_
rlabel metal2 18872 35392 18872 35392 0 _0961_
rlabel metal3 20104 35784 20104 35784 0 _0962_
rlabel metal2 12712 33880 12712 33880 0 _0963_
rlabel metal3 8848 33320 8848 33320 0 _0964_
rlabel metal2 5656 32088 5656 32088 0 _0965_
rlabel metal3 7952 32648 7952 32648 0 _0966_
rlabel metal2 11032 32704 11032 32704 0 _0967_
rlabel metal2 10248 32704 10248 32704 0 _0968_
rlabel metal2 11704 24080 11704 24080 0 _0969_
rlabel metal3 11984 33208 11984 33208 0 _0970_
rlabel metal2 14728 33768 14728 33768 0 _0971_
rlabel metal2 20216 34888 20216 34888 0 _0972_
rlabel metal2 27048 37688 27048 37688 0 _0973_
rlabel metal3 36624 68488 36624 68488 0 _0974_
rlabel metal2 40712 64400 40712 64400 0 _0975_
rlabel metal2 41832 62244 41832 62244 0 _0976_
rlabel metal2 40208 60200 40208 60200 0 _0977_
rlabel metal2 41048 60256 41048 60256 0 _0978_
rlabel metal3 42784 61656 42784 61656 0 _0979_
rlabel metal2 41160 54208 41160 54208 0 _0980_
rlabel metal2 40768 55272 40768 55272 0 _0981_
rlabel metal2 12096 26488 12096 26488 0 _0982_
rlabel metal2 14560 23240 14560 23240 0 _0983_
rlabel metal2 13944 21840 13944 21840 0 _0984_
rlabel metal2 38696 45024 38696 45024 0 _0985_
rlabel metal2 40432 47320 40432 47320 0 _0986_
rlabel metal2 41272 49840 41272 49840 0 _0987_
rlabel metal2 41272 56560 41272 56560 0 _0988_
rlabel metal2 42168 58800 42168 58800 0 _0989_
rlabel metal2 40040 64400 40040 64400 0 _0990_
rlabel metal2 39704 66304 39704 66304 0 _0991_
rlabel metal2 39592 65744 39592 65744 0 _0992_
rlabel metal2 33768 60480 33768 60480 0 _0993_
rlabel metal2 36120 60760 36120 60760 0 _0994_
rlabel metal3 36848 60536 36848 60536 0 _0995_
rlabel metal2 37016 60816 37016 60816 0 _0996_
rlabel metal2 32536 72408 32536 72408 0 _0997_
rlabel metal3 35840 60872 35840 60872 0 _0998_
rlabel metal2 37576 62552 37576 62552 0 _0999_
rlabel metal2 36792 63056 36792 63056 0 _1000_
rlabel metal2 38360 65968 38360 65968 0 _1001_
rlabel metal2 39816 68656 39816 68656 0 _1002_
rlabel metal3 39144 68600 39144 68600 0 _1003_
rlabel metal2 22120 34776 22120 34776 0 _1004_
rlabel metal3 16184 30184 16184 30184 0 _1005_
rlabel metal3 15792 30296 15792 30296 0 _1006_
rlabel metal2 16072 31360 16072 31360 0 _1007_
rlabel metal2 14392 33432 14392 33432 0 _1008_
rlabel metal2 16856 33880 16856 33880 0 _1009_
rlabel metal2 15848 33320 15848 33320 0 _1010_
rlabel metal2 12264 29232 12264 29232 0 _1011_
rlabel metal2 10808 29848 10808 29848 0 _1012_
rlabel metal3 7280 32312 7280 32312 0 _1013_
rlabel metal2 8904 30408 8904 30408 0 _1014_
rlabel via2 4872 30968 4872 30968 0 _1015_
rlabel metal2 6664 32480 6664 32480 0 _1016_
rlabel metal2 7784 31360 7784 31360 0 _1017_
rlabel metal2 8344 24976 8344 24976 0 _1018_
rlabel metal2 8456 27440 8456 27440 0 _1019_
rlabel metal2 5880 25536 5880 25536 0 _1020_
rlabel metal2 8344 25480 8344 25480 0 _1021_
rlabel metal2 10360 26768 10360 26768 0 _1022_
rlabel metal2 11928 24080 11928 24080 0 _1023_
rlabel metal2 12936 30576 12936 30576 0 _1024_
rlabel metal2 16352 30744 16352 30744 0 _1025_
rlabel metal3 23072 31528 23072 31528 0 _1026_
rlabel metal2 20664 35336 20664 35336 0 _1027_
rlabel metal2 21672 35280 21672 35280 0 _1028_
rlabel metal2 23240 30464 23240 30464 0 _1029_
rlabel metal3 35112 69160 35112 69160 0 _1030_
rlabel metal2 41720 60648 41720 60648 0 _1031_
rlabel metal2 42280 62244 42280 62244 0 _1032_
rlabel metal3 42336 62328 42336 62328 0 _1033_
rlabel metal2 42840 54544 42840 54544 0 _1034_
rlabel metal2 43176 54432 43176 54432 0 _1035_
rlabel metal2 43736 56784 43736 56784 0 _1036_
rlabel metal3 40880 48888 40880 48888 0 _1037_
rlabel metal2 40544 49112 40544 49112 0 _1038_
rlabel metal2 40880 51128 40880 51128 0 _1039_
rlabel metal2 43176 55832 43176 55832 0 _1040_
rlabel metal2 41832 47544 41832 47544 0 _1041_
rlabel metal3 12544 12936 12544 12936 0 _1042_
rlabel metal2 12768 12712 12768 12712 0 _1043_
rlabel metal2 28728 20328 28728 20328 0 _1044_
rlabel metal3 41552 45864 41552 45864 0 _1045_
rlabel metal2 42280 46928 42280 46928 0 _1046_
rlabel metal2 43568 49224 43568 49224 0 _1047_
rlabel metal2 43512 58072 43512 58072 0 _1048_
rlabel metal2 43736 62272 43736 62272 0 _1049_
rlabel metal2 42504 62552 42504 62552 0 _1050_
rlabel metal2 43064 64736 43064 64736 0 _1051_
rlabel metal2 42392 66584 42392 66584 0 _1052_
rlabel metal2 41272 65576 41272 65576 0 _1053_
rlabel metal2 40040 65744 40040 65744 0 _1054_
rlabel metal2 41384 66640 41384 66640 0 _1055_
rlabel metal2 40488 68208 40488 68208 0 _1056_
rlabel metal2 39144 68152 39144 68152 0 _1057_
rlabel metal2 25928 69552 25928 69552 0 _1058_
rlabel metal2 25928 70672 25928 70672 0 _1059_
rlabel metal2 40600 68096 40600 68096 0 _1060_
rlabel via2 42280 67704 42280 67704 0 _1061_
rlabel metal2 42616 66640 42616 66640 0 _1062_
rlabel metal2 44184 54880 44184 54880 0 _1063_
rlabel metal3 21336 32536 21336 32536 0 _1064_
rlabel metal3 23072 31752 23072 31752 0 _1065_
rlabel metal2 22064 31752 22064 31752 0 _1066_
rlabel metal2 18200 29960 18200 29960 0 _1067_
rlabel metal2 16408 31640 16408 31640 0 _1068_
rlabel metal3 17528 30856 17528 30856 0 _1069_
rlabel metal2 18088 30576 18088 30576 0 _1070_
rlabel metal2 16240 25480 16240 25480 0 _1071_
rlabel metal3 15568 27832 15568 27832 0 _1072_
rlabel metal2 15176 25928 15176 25928 0 _1073_
rlabel metal2 15848 25816 15848 25816 0 _1074_
rlabel metal2 16968 26992 16968 26992 0 _1075_
rlabel metal2 11480 24024 11480 24024 0 _1076_
rlabel metal2 11704 28000 11704 28000 0 _1077_
rlabel metal2 12936 27496 12936 27496 0 _1078_
rlabel metal2 13832 27384 13832 27384 0 _1079_
rlabel metal2 10920 25032 10920 25032 0 _1080_
rlabel metal2 9800 27272 9800 27272 0 _1081_
rlabel metal2 7728 22344 7728 22344 0 _1082_
rlabel metal2 7224 24696 7224 24696 0 _1083_
rlabel metal2 8400 22344 8400 22344 0 _1084_
rlabel metal2 10136 19600 10136 19600 0 _1085_
rlabel metal2 10808 22400 10808 22400 0 _1086_
rlabel metal3 13160 27048 13160 27048 0 _1087_
rlabel metal2 17752 27048 17752 27048 0 _1088_
rlabel metal3 18648 29512 18648 29512 0 _1089_
rlabel metal2 23576 30576 23576 30576 0 _1090_
rlabel metal2 43456 44520 43456 44520 0 _1091_
rlabel metal2 44968 55216 44968 55216 0 _1092_
rlabel metal2 43400 57512 43400 57512 0 _1093_
rlabel metal2 43960 57568 43960 57568 0 _1094_
rlabel metal2 44520 57904 44520 57904 0 _1095_
rlabel metal2 42616 47544 42616 47544 0 _1096_
rlabel metal2 42896 46088 42896 46088 0 _1097_
rlabel metal3 43288 46648 43288 46648 0 _1098_
rlabel metal2 41496 44688 41496 44688 0 _1099_
rlabel metal2 42056 43596 42056 43596 0 _1100_
rlabel metal2 9576 22792 9576 22792 0 _1101_
rlabel metal2 14560 20104 14560 20104 0 _1102_
rlabel metal2 15176 19656 15176 19656 0 _1103_
rlabel metal2 41552 43512 41552 43512 0 _1104_
rlabel metal2 42616 43624 42616 43624 0 _1105_
rlabel metal2 44072 46200 44072 46200 0 _1106_
rlabel metal2 44520 47544 44520 47544 0 _1107_
rlabel metal2 43736 49672 43736 49672 0 _1108_
rlabel metal3 42336 51352 42336 51352 0 _1109_
rlabel metal2 40712 44464 40712 44464 0 _1110_
rlabel metal2 42728 51576 42728 51576 0 _1111_
rlabel metal2 43064 50456 43064 50456 0 _1112_
rlabel metal2 44184 49336 44184 49336 0 _1113_
rlabel metal2 44296 49504 44296 49504 0 _1114_
rlabel metal2 45192 58128 45192 58128 0 _1115_
rlabel metal2 44968 59976 44968 59976 0 _1116_
rlabel metal2 44296 62608 44296 62608 0 _1117_
rlabel metal2 44072 62888 44072 62888 0 _1118_
rlabel metal2 43288 65072 43288 65072 0 _1119_
rlabel metal2 43176 68600 43176 68600 0 _1120_
rlabel metal2 27384 70224 27384 70224 0 _1121_
rlabel metal2 26544 70280 26544 70280 0 _1122_
rlabel metal2 26544 74088 26544 74088 0 _1123_
rlabel metal2 27328 69272 27328 69272 0 _1124_
rlabel metal2 26152 68880 26152 68880 0 _1125_
rlabel metal2 44800 61768 44800 61768 0 _1126_
rlabel metal2 45416 62832 45416 62832 0 _1127_
rlabel metal2 43848 67452 43848 67452 0 _1128_
rlabel metal2 46032 62552 46032 62552 0 _1129_
rlabel metal2 42952 53816 42952 53816 0 _1130_
rlabel metal2 45304 54040 45304 54040 0 _1131_
rlabel metal2 46032 57848 46032 57848 0 _1132_
rlabel metal2 45192 57008 45192 57008 0 _1133_
rlabel metal2 45640 55496 45640 55496 0 _1134_
rlabel metal2 43960 50904 43960 50904 0 _1135_
rlabel metal2 43512 50624 43512 50624 0 _1136_
rlabel metal3 44968 50232 44968 50232 0 _1137_
rlabel metal2 38808 27664 38808 27664 0 _1138_
rlabel metal2 21784 30744 21784 30744 0 _1139_
rlabel metal2 39144 29680 39144 29680 0 _1140_
rlabel metal2 39032 27552 39032 27552 0 _1141_
rlabel metal3 22176 27944 22176 27944 0 _1142_
rlabel metal2 19320 29288 19320 29288 0 _1143_
rlabel metal2 18872 28952 18872 28952 0 _1144_
rlabel metal3 20384 28616 20384 28616 0 _1145_
rlabel metal2 23072 25144 23072 25144 0 _1146_
rlabel metal2 16800 26040 16800 26040 0 _1147_
rlabel metal3 19488 25480 19488 25480 0 _1148_
rlabel metal2 18424 25256 18424 25256 0 _1149_
rlabel metal2 19096 25312 19096 25312 0 _1150_
rlabel metal2 13888 26488 13888 26488 0 _1151_
rlabel metal2 18536 26488 18536 26488 0 _1152_
rlabel metal2 15736 21168 15736 21168 0 _1153_
rlabel metal2 14616 22680 14616 22680 0 _1154_
rlabel metal2 14728 22680 14728 22680 0 _1155_
rlabel metal2 15848 21504 15848 21504 0 _1156_
rlabel metal2 16968 21168 16968 21168 0 _1157_
rlabel metal3 12488 23912 12488 23912 0 _1158_
rlabel metal3 11480 22456 11480 22456 0 _1159_
rlabel metal2 10696 23744 10696 23744 0 _1160_
rlabel metal3 11928 20104 11928 20104 0 _1161_
rlabel metal2 11256 19880 11256 19880 0 _1162_
rlabel metal3 11480 18536 11480 18536 0 _1163_
rlabel metal3 11928 18200 11928 18200 0 _1164_
rlabel metal3 12208 18424 12208 18424 0 _1165_
rlabel metal2 17192 19712 17192 19712 0 _1166_
rlabel metal2 18760 23968 18760 23968 0 _1167_
rlabel metal2 20888 26628 20888 26628 0 _1168_
rlabel metal2 37016 27440 37016 27440 0 _1169_
rlabel metal2 45360 48104 45360 48104 0 _1170_
rlabel metal2 44856 45080 44856 45080 0 _1171_
rlabel metal2 44744 46704 44744 46704 0 _1172_
rlabel metal2 45080 45024 45080 45024 0 _1173_
rlabel metal2 46536 44520 46536 44520 0 _1174_
rlabel metal2 43120 42840 43120 42840 0 _1175_
rlabel metal2 42112 31864 42112 31864 0 _1176_
rlabel metal3 36120 48776 36120 48776 0 _1177_
rlabel metal2 42728 42952 42728 42952 0 _1178_
rlabel metal2 45304 40600 45304 40600 0 _1179_
rlabel metal2 39368 41664 39368 41664 0 _1180_
rlabel metal2 40040 40600 40040 40600 0 _1181_
rlabel metal2 41440 34888 41440 34888 0 _1182_
rlabel metal2 43400 36456 43400 36456 0 _1183_
rlabel metal3 41496 37240 41496 37240 0 _1184_
rlabel metal2 43512 37184 43512 37184 0 _1185_
rlabel metal2 44856 38360 44856 38360 0 _1186_
rlabel metal2 46088 40768 46088 40768 0 _1187_
rlabel metal3 41328 40376 41328 40376 0 _1188_
rlabel metal2 42616 39872 42616 39872 0 _1189_
rlabel metal2 43064 39648 43064 39648 0 _1190_
rlabel via2 43624 39928 43624 39928 0 _1191_
rlabel metal2 45416 40824 45416 40824 0 _1192_
rlabel metal2 45080 41440 45080 41440 0 _1193_
rlabel metal2 45864 41552 45864 41552 0 _1194_
rlabel metal2 46424 43512 46424 43512 0 _1195_
rlabel metal2 46872 43904 46872 43904 0 _1196_
rlabel metal2 46312 54040 46312 54040 0 _1197_
rlabel metal3 46144 63112 46144 63112 0 _1198_
rlabel metal2 27384 68152 27384 68152 0 _1199_
rlabel metal2 26264 68152 26264 68152 0 _1200_
rlabel metal2 25536 68712 25536 68712 0 _1201_
rlabel metal2 26936 67816 26936 67816 0 _1202_
rlabel metal2 25928 65016 25928 65016 0 _1203_
rlabel metal2 45752 62720 45752 62720 0 _1204_
rlabel metal2 46312 62608 46312 62608 0 _1205_
rlabel metal2 45864 62188 45864 62188 0 _1206_
rlabel metal2 46200 49392 46200 49392 0 _1207_
rlabel metal2 46144 53704 46144 53704 0 _1208_
rlabel metal2 46536 54376 46536 54376 0 _1209_
rlabel metal2 45976 51744 45976 51744 0 _1210_
rlabel metal3 46928 43512 46928 43512 0 _1211_
rlabel metal2 47432 43568 47432 43568 0 _1212_
rlabel metal2 46984 42056 46984 42056 0 _1213_
rlabel metal2 44968 39004 44968 39004 0 _1214_
rlabel metal3 42280 24696 42280 24696 0 _1215_
rlabel metal2 43288 34832 43288 34832 0 _1216_
rlabel metal2 38864 23352 38864 23352 0 _1217_
rlabel metal3 41888 34888 41888 34888 0 _1218_
rlabel metal2 43456 34104 43456 34104 0 _1219_
rlabel metal2 42112 22344 42112 22344 0 _1220_
rlabel metal2 43624 33824 43624 33824 0 _1221_
rlabel metal3 21840 16968 21840 16968 0 _1222_
rlabel metal2 40040 29848 40040 29848 0 _1223_
rlabel metal2 41608 31248 41608 31248 0 _1224_
rlabel metal2 41832 33992 41832 33992 0 _1225_
rlabel metal2 40712 29736 40712 29736 0 _1226_
rlabel metal3 41776 30184 41776 30184 0 _1227_
rlabel metal2 41272 30184 41272 30184 0 _1228_
rlabel metal2 42616 31248 42616 31248 0 _1229_
rlabel metal2 42952 32536 42952 32536 0 _1230_
rlabel metal2 44856 34104 44856 34104 0 _1231_
rlabel metal2 45416 36456 45416 36456 0 _1232_
rlabel metal2 39368 28280 39368 28280 0 _1233_
rlabel metal2 43400 29176 43400 29176 0 _1234_
rlabel metal2 43344 38808 43344 38808 0 _1235_
rlabel metal3 43904 38920 43904 38920 0 _1236_
rlabel metal2 42616 29848 42616 29848 0 _1237_
rlabel metal2 22904 24696 22904 24696 0 _1238_
rlabel metal2 23632 24920 23632 24920 0 _1239_
rlabel metal2 22232 26544 22232 26544 0 _1240_
rlabel metal2 24024 26572 24024 26572 0 _1241_
rlabel metal2 25704 24080 25704 24080 0 _1242_
rlabel metal2 33992 23072 33992 23072 0 _1243_
rlabel metal2 21336 22792 21336 22792 0 _1244_
rlabel metal2 20104 24808 20104 24808 0 _1245_
rlabel metal2 19432 24640 19432 24640 0 _1246_
rlabel metal2 21392 23800 21392 23800 0 _1247_
rlabel metal2 16072 21448 16072 21448 0 _1248_
rlabel metal3 20384 20776 20384 20776 0 _1249_
rlabel metal2 18984 21224 18984 21224 0 _1250_
rlabel metal2 19712 19992 19712 19992 0 _1251_
rlabel metal2 19992 20608 19992 20608 0 _1252_
rlabel metal2 20328 19096 20328 19096 0 _1253_
rlabel metal2 12936 18816 12936 18816 0 _1254_
rlabel metal3 11256 19208 11256 19208 0 _1255_
rlabel metal2 11816 19684 11816 19684 0 _1256_
rlabel metal3 13160 18984 13160 18984 0 _1257_
rlabel metal2 11816 13552 11816 13552 0 _1258_
rlabel metal3 12432 19096 12432 19096 0 _1259_
rlabel metal2 14056 19712 14056 19712 0 _1260_
rlabel metal3 18200 18424 18200 18424 0 _1261_
rlabel metal2 15624 18312 15624 18312 0 _1262_
rlabel metal2 15848 17976 15848 17976 0 _1263_
rlabel metal2 15960 17696 15960 17696 0 _1264_
rlabel metal2 17416 16324 17416 16324 0 _1265_
rlabel metal3 12264 15400 12264 15400 0 _1266_
rlabel metal2 11144 14784 11144 14784 0 _1267_
rlabel metal2 11592 14840 11592 14840 0 _1268_
rlabel metal2 12320 14616 12320 14616 0 _1269_
rlabel metal2 13552 6664 13552 6664 0 _1270_
rlabel metal2 17976 15148 17976 15148 0 _1271_
rlabel metal2 18760 18088 18760 18088 0 _1272_
rlabel metal3 19656 18312 19656 18312 0 _1273_
rlabel metal2 20104 22232 20104 22232 0 _1274_
rlabel metal3 23240 23800 23240 23800 0 _1275_
rlabel metal2 34216 23856 34216 23856 0 _1276_
rlabel metal2 37800 22344 37800 22344 0 _1277_
rlabel metal2 38696 20440 38696 20440 0 _1278_
rlabel metal2 38416 22232 38416 22232 0 _1279_
rlabel metal2 37128 23520 37128 23520 0 _1280_
rlabel metal2 43960 29848 43960 29848 0 _1281_
rlabel metal2 46088 34328 46088 34328 0 _1282_
rlabel metal3 47768 49784 47768 49784 0 _1283_
rlabel metal3 47040 49896 47040 49896 0 _1284_
rlabel metal2 28056 62664 28056 62664 0 _1285_
rlabel metal2 26040 64344 26040 64344 0 _1286_
rlabel metal3 21056 64792 21056 64792 0 _1287_
rlabel metal2 25480 63616 25480 63616 0 _1288_
rlabel metal2 26992 62440 26992 62440 0 _1289_
rlabel metal2 46088 49952 46088 49952 0 _1290_
rlabel metal2 46760 57176 46760 57176 0 _1291_
rlabel metal2 47096 33824 47096 33824 0 _1292_
rlabel metal2 45528 35504 45528 35504 0 _1293_
rlabel metal2 46760 35784 46760 35784 0 _1294_
rlabel metal2 47208 34664 47208 34664 0 _1295_
rlabel metal2 47320 33208 47320 33208 0 _1296_
rlabel metal2 44016 29400 44016 29400 0 _1297_
rlabel metal3 44576 28504 44576 28504 0 _1298_
rlabel metal2 44744 29288 44744 29288 0 _1299_
rlabel metal3 45976 28728 45976 28728 0 _1300_
rlabel metal2 45304 31808 45304 31808 0 _1301_
rlabel metal3 45416 34216 45416 34216 0 _1302_
rlabel metal2 45192 26628 45192 26628 0 _1303_
rlabel metal2 43792 26264 43792 26264 0 _1304_
rlabel metal2 42336 24808 42336 24808 0 _1305_
rlabel metal2 41944 24304 41944 24304 0 _1306_
rlabel metal2 36680 13552 36680 13552 0 _1307_
rlabel metal2 40600 25312 40600 25312 0 _1308_
rlabel metal2 34496 48776 34496 48776 0 _1309_
rlabel metal3 33936 17080 33936 17080 0 _1310_
rlabel metal3 40712 24696 40712 24696 0 _1311_
rlabel metal2 39368 22736 39368 22736 0 _1312_
rlabel metal3 40880 24808 40880 24808 0 _1313_
rlabel metal2 42504 25088 42504 25088 0 _1314_
rlabel metal2 43680 25592 43680 25592 0 _1315_
rlabel metal3 44520 26152 44520 26152 0 _1316_
rlabel metal2 37688 24248 37688 24248 0 _1317_
rlabel metal2 38472 22680 38472 22680 0 _1318_
rlabel metal2 42280 21728 42280 21728 0 _1319_
rlabel metal2 42784 21560 42784 21560 0 _1320_
rlabel metal2 23016 23632 23016 23632 0 _1321_
rlabel metal3 24360 23912 24360 23912 0 _1322_
rlabel metal2 24024 23520 24024 23520 0 _1323_
rlabel metal2 26600 19768 26600 19768 0 _1324_
rlabel metal2 35448 14448 35448 14448 0 _1325_
rlabel metal3 20944 22456 20944 22456 0 _1326_
rlabel metal2 21784 23016 21784 23016 0 _1327_
rlabel metal2 23408 15624 23408 15624 0 _1328_
rlabel metal2 22456 19208 22456 19208 0 _1329_
rlabel metal2 22792 19600 22792 19600 0 _1330_
rlabel metal2 23184 18984 23184 18984 0 _1331_
rlabel metal3 19544 17528 19544 17528 0 _1332_
rlabel metal2 20440 16268 20440 16268 0 _1333_
rlabel metal2 17976 11088 17976 11088 0 _1334_
rlabel metal2 14280 6272 14280 6272 0 _1335_
rlabel metal2 14056 5768 14056 5768 0 _1336_
rlabel metal2 12264 11536 12264 11536 0 _1337_
rlabel metal2 12712 12264 12712 12264 0 _1338_
rlabel metal2 13496 14672 13496 14672 0 _1339_
rlabel metal2 14392 10136 14392 10136 0 _1340_
rlabel metal2 14392 9352 14392 9352 0 _1341_
rlabel metal2 19712 10584 19712 10584 0 _1342_
rlabel metal2 16016 16856 16016 16856 0 _1343_
rlabel metal2 16632 17640 16632 17640 0 _1344_
rlabel metal3 19936 16856 19936 16856 0 _1345_
rlabel metal2 17080 21224 17080 21224 0 _1346_
rlabel metal3 21000 16072 21000 16072 0 _1347_
rlabel metal2 22120 17976 22120 17976 0 _1348_
rlabel metal2 19208 11088 19208 11088 0 _1349_
rlabel metal2 20776 10528 20776 10528 0 _1350_
rlabel metal2 22792 10920 22792 10920 0 _1351_
rlabel metal2 24472 12264 24472 12264 0 _1352_
rlabel metal3 37128 14616 37128 14616 0 _1353_
rlabel metal2 39592 13720 39592 13720 0 _1354_
rlabel metal3 37072 14504 37072 14504 0 _1355_
rlabel metal2 38472 13664 38472 13664 0 _1356_
rlabel metal2 40152 15260 40152 15260 0 _1357_
rlabel metal2 41832 19096 41832 19096 0 _1358_
rlabel metal3 45864 25592 45864 25592 0 _1359_
rlabel metal2 47432 26432 47432 26432 0 _1360_
rlabel metal2 47096 30632 47096 30632 0 _1361_
rlabel metal2 46760 33880 46760 33880 0 _1362_
rlabel metal2 26488 48888 26488 48888 0 _1363_
rlabel metal2 26264 64064 26264 64064 0 _1364_
rlabel metal2 28336 27048 28336 27048 0 _1365_
rlabel metal2 27944 26096 27944 26096 0 _1366_
rlabel metal2 29064 25760 29064 25760 0 _1367_
rlabel metal3 46368 33320 46368 33320 0 _1368_
rlabel metal2 45472 21784 45472 21784 0 _1369_
rlabel metal2 45864 25648 45864 25648 0 _1370_
rlabel metal2 45976 26432 45976 26432 0 _1371_
rlabel metal3 46536 25480 46536 25480 0 _1372_
rlabel metal3 46032 23352 46032 23352 0 _1373_
rlabel via2 40152 14504 40152 14504 0 _1374_
rlabel metal2 41888 14616 41888 14616 0 _1375_
rlabel metal2 42952 16016 42952 16016 0 _1376_
rlabel metal2 42896 19880 42896 19880 0 _1377_
rlabel metal2 43344 16296 43344 16296 0 _1378_
rlabel metal2 44856 16520 44856 16520 0 _1379_
rlabel metal2 44576 24696 44576 24696 0 _1380_
rlabel metal3 44464 24472 44464 24472 0 _1381_
rlabel metal2 43288 18592 43288 18592 0 _1382_
rlabel metal2 40264 21056 40264 21056 0 _1383_
rlabel metal2 39480 19992 39480 19992 0 _1384_
rlabel metal2 39928 19152 39928 19152 0 _1385_
rlabel metal2 40264 19264 40264 19264 0 _1386_
rlabel metal2 41608 20608 41608 20608 0 _1387_
rlabel metal2 42896 17528 42896 17528 0 _1388_
rlabel metal2 44072 12936 44072 12936 0 _1389_
rlabel metal3 39592 12936 39592 12936 0 _1390_
rlabel metal2 40320 12936 40320 12936 0 _1391_
rlabel metal3 42000 12824 42000 12824 0 _1392_
rlabel metal2 40824 23632 40824 23632 0 _1393_
rlabel metal2 40376 24192 40376 24192 0 _1394_
rlabel metal2 41048 12656 41048 12656 0 _1395_
rlabel metal2 24024 13888 24024 13888 0 _1396_
rlabel metal2 27160 13664 27160 13664 0 _1397_
rlabel metal2 33880 6048 33880 6048 0 _1398_
rlabel metal2 22232 10304 22232 10304 0 _1399_
rlabel metal2 23576 8372 23576 8372 0 _1400_
rlabel metal2 21336 16352 21336 16352 0 _1401_
rlabel metal2 21784 8288 21784 8288 0 _1402_
rlabel metal3 19208 9688 19208 9688 0 _1403_
rlabel metal3 20384 8008 20384 8008 0 _1404_
rlabel metal2 16520 8288 16520 8288 0 _1405_
rlabel metal2 14840 14112 14840 14112 0 _1406_
rlabel metal2 15848 13048 15848 13048 0 _1407_
rlabel metal2 14728 12600 14728 12600 0 _1408_
rlabel metal2 15064 11648 15064 11648 0 _1409_
rlabel metal2 15176 10304 15176 10304 0 _1410_
rlabel metal2 16632 8288 16632 8288 0 _1411_
rlabel metal2 18648 8176 18648 8176 0 _1412_
rlabel metal2 11704 11368 11704 11368 0 _1413_
rlabel metal2 12712 11648 12712 11648 0 _1414_
rlabel metal2 18200 11648 18200 11648 0 _1415_
rlabel metal2 18760 12768 18760 12768 0 _1416_
rlabel metal2 19264 12264 19264 12264 0 _1417_
rlabel metal2 20440 26880 20440 26880 0 _1418_
rlabel metal2 19992 11648 19992 11648 0 _1419_
rlabel metal2 18984 13104 18984 13104 0 _1420_
rlabel metal2 18760 8848 18760 8848 0 _1421_
rlabel metal3 19992 8120 19992 8120 0 _1422_
rlabel metal2 21896 7952 21896 7952 0 _1423_
rlabel metal3 23072 8232 23072 8232 0 _1424_
rlabel metal2 33656 5824 33656 5824 0 _1425_
rlabel metal2 37688 11256 37688 11256 0 _1426_
rlabel metal2 28224 11368 28224 11368 0 _1427_
rlabel metal3 36904 9016 36904 9016 0 _1428_
rlabel metal2 38472 5096 38472 5096 0 _1429_
rlabel metal3 40264 11928 40264 11928 0 _1430_
rlabel metal2 45080 14112 45080 14112 0 _1431_
rlabel metal2 45192 16016 45192 16016 0 _1432_
rlabel metal2 45976 19712 45976 19712 0 _1433_
rlabel metal2 45528 22904 45528 22904 0 _1434_
rlabel metal2 28616 25200 28616 25200 0 _1435_
rlabel metal2 27608 25256 27608 25256 0 _1436_
rlabel metal2 28336 26264 28336 26264 0 _1437_
rlabel metal3 27160 23128 27160 23128 0 _1438_
rlabel metal2 26264 22512 26264 22512 0 _1439_
rlabel metal2 45304 21952 45304 21952 0 _1440_
rlabel metal2 45864 22232 45864 22232 0 _1441_
rlabel metal2 45416 21112 45416 21112 0 _1442_
rlabel metal2 43456 11928 43456 11928 0 _1443_
rlabel metal3 44856 14504 44856 14504 0 _1444_
rlabel metal3 44744 15848 44744 15848 0 _1445_
rlabel metal2 45528 15848 45528 15848 0 _1446_
rlabel metal2 45416 19040 45416 19040 0 _1447_
rlabel metal3 41944 12040 41944 12040 0 _1448_
rlabel metal2 41944 11648 41944 11648 0 _1449_
rlabel metal2 42504 11480 42504 11480 0 _1450_
rlabel metal2 42168 10472 42168 10472 0 _1451_
rlabel metal2 43288 16072 43288 16072 0 _1452_
rlabel metal2 44072 10248 44072 10248 0 _1453_
rlabel metal2 35672 5824 35672 5824 0 _1454_
rlabel metal2 37800 5936 37800 5936 0 _1455_
rlabel metal2 38920 4760 38920 4760 0 _1456_
rlabel metal2 38696 19488 38696 19488 0 _1457_
rlabel metal2 39872 17528 39872 17528 0 _1458_
rlabel metal2 24136 7728 24136 7728 0 _1459_
rlabel metal2 24360 6776 24360 6776 0 _1460_
rlabel metal2 25704 6608 25704 6608 0 _1461_
rlabel metal2 21336 7952 21336 7952 0 _1462_
rlabel metal2 11592 36176 11592 36176 0 a\[0\]\[0\]
rlabel metal2 9520 28616 9520 28616 0 a\[0\]\[1\]
rlabel metal2 10584 16072 10584 16072 0 a\[0\]\[2\]
rlabel metal2 15008 37352 15008 37352 0 a\[0\]\[3\]
rlabel metal2 14448 37128 14448 37128 0 a\[0\]\[4\]
rlabel metal2 16408 39172 16408 39172 0 a\[0\]\[5\]
rlabel metal2 18424 22064 18424 22064 0 a\[0\]\[6\]
rlabel metal2 20440 40264 20440 40264 0 a\[0\]\[7\]
rlabel metal2 15232 49784 15232 49784 0 a\[1\]\[0\]
rlabel metal2 22232 72464 22232 72464 0 a\[1\]\[1\]
rlabel metal2 20664 69832 20664 69832 0 a\[1\]\[2\]
rlabel metal2 17976 72744 17976 72744 0 a\[1\]\[3\]
rlabel metal2 18144 62552 18144 62552 0 a\[1\]\[4\]
rlabel metal2 24360 73192 24360 73192 0 a\[1\]\[5\]
rlabel metal3 24304 62216 24304 62216 0 a\[1\]\[6\]
rlabel metal2 20328 69944 20328 69944 0 a\[1\]\[7\]
rlabel metal2 2520 77882 2520 77882 0 active
rlabel metal2 28840 55776 28840 55776 0 b\[0\]\[0\]
rlabel metal2 40208 46536 40208 46536 0 b\[0\]\[1\]
rlabel metal2 40040 48048 40040 48048 0 b\[0\]\[2\]
rlabel metal2 41048 53088 41048 53088 0 b\[0\]\[3\]
rlabel metal2 41720 42280 41720 42280 0 b\[0\]\[4\]
rlabel metal3 40320 49896 40320 49896 0 b\[0\]\[5\]
rlabel metal2 37240 25144 37240 25144 0 b\[0\]\[6\]
rlabel metal2 37688 14532 37688 14532 0 b\[0\]\[7\]
rlabel metal2 15512 66864 15512 66864 0 b\[1\]\[0\]
rlabel metal2 16632 71232 16632 71232 0 b\[1\]\[1\]
rlabel metal2 17080 70392 17080 70392 0 b\[1\]\[2\]
rlabel metal3 17136 73192 17136 73192 0 b\[1\]\[3\]
rlabel metal2 19040 66360 19040 66360 0 b\[1\]\[4\]
rlabel metal2 24584 66920 24584 66920 0 b\[1\]\[5\]
rlabel metal3 23688 67144 23688 67144 0 b\[1\]\[6\]
rlabel metal2 20776 68656 20776 68656 0 b\[1\]\[7\]
rlabel metal3 7168 67592 7168 67592 0 bflip
rlabel metal2 33320 42280 33320 42280 0 c\[0\]\[0\]
rlabel metal2 31528 46984 31528 46984 0 c\[0\]\[1\]
rlabel metal2 29960 45472 29960 45472 0 c\[0\]\[2\]
rlabel metal2 29848 43736 29848 43736 0 c\[0\]\[3\]
rlabel metal2 31976 41888 31976 41888 0 c\[0\]\[4\]
rlabel metal2 32424 39312 32424 39312 0 c\[0\]\[5\]
rlabel metal3 32704 18424 32704 18424 0 c\[0\]\[6\]
rlabel metal2 37072 13944 37072 13944 0 c\[0\]\[7\]
rlabel metal2 16296 48496 16296 48496 0 c\[1\]\[0\]
rlabel metal2 17752 52864 17752 52864 0 c\[1\]\[1\]
rlabel metal2 16968 54376 16968 54376 0 c\[1\]\[2\]
rlabel metal2 16688 57736 16688 57736 0 c\[1\]\[3\]
rlabel metal2 13832 57624 13832 57624 0 c\[1\]\[4\]
rlabel metal2 13608 54992 13608 54992 0 c\[1\]\[5\]
rlabel metal2 20664 53144 20664 53144 0 c\[1\]\[6\]
rlabel metal2 20720 50904 20720 50904 0 c\[1\]\[7\]
rlabel metal2 23800 47880 23800 47880 0 clk
rlabel metal3 21112 48104 21112 48104 0 clknet_0_clk
rlabel metal2 1904 35672 1904 35672 0 clknet_1_0__leaf_clk
rlabel metal3 6664 73976 6664 73976 0 clknet_1_1__leaf_clk
rlabel metal2 7336 61712 7336 61712 0 delta_t\[0\]
rlabel metal2 7952 60088 7952 60088 0 delta_t\[1\]
rlabel metal3 4928 52136 4928 52136 0 delta_t\[2\]
rlabel metal2 8344 52808 8344 52808 0 delta_t\[3\]
rlabel metal2 23744 49672 23744 49672 0 delta_t\[4\]
rlabel metal2 3192 42280 3192 42280 0 delta_t\[5\]
rlabel metal3 4312 39032 4312 39032 0 delta_t\[6\]
rlabel metal3 20328 35896 20328 35896 0 delta_t\[7\]
rlabel metal2 6496 25480 6496 25480 0 delta_t\[8\]
rlabel metal2 6104 24864 6104 24864 0 delta_t\[9\]
rlabel metal2 3136 20160 3136 20160 0 net1
rlabel metal2 15904 64792 15904 64792 0 net10
rlabel metal2 48216 33936 48216 33936 0 net100
rlabel metal2 48216 36176 48216 36176 0 net101
rlabel metal2 48216 38808 48216 38808 0 net102
rlabel metal2 48216 61040 48216 61040 0 net103
rlabel metal2 48216 63616 48216 63616 0 net104
rlabel metal2 48216 65856 48216 65856 0 net105
rlabel metal2 48216 68432 48216 68432 0 net106
rlabel metal2 48216 70672 48216 70672 0 net107
rlabel metal2 48216 73248 48216 73248 0 net108
rlabel metal3 48762 75544 48762 75544 0 net109
rlabel metal2 2184 73528 2184 73528 0 net11
rlabel metal2 48216 77336 48216 77336 0 net110
rlabel metal2 21448 30632 21448 30632 0 net111
rlabel metal2 22680 31472 22680 31472 0 net112
rlabel metal2 36568 31808 36568 31808 0 net113
rlabel metal2 38584 35896 38584 35896 0 net114
rlabel metal2 32984 30856 32984 30856 0 net115
rlabel metal2 31640 61544 31640 61544 0 net116
rlabel metal2 39704 37576 39704 37576 0 net117
rlabel metal2 10920 30240 10920 30240 0 net118
rlabel metal2 21784 28672 21784 28672 0 net119
rlabel metal2 16408 62832 16408 62832 0 net12
rlabel metal2 17416 32200 17416 32200 0 net120
rlabel metal2 9912 32984 9912 32984 0 net121
rlabel metal2 23128 25816 23128 25816 0 net122
rlabel metal2 27384 21840 27384 21840 0 net123
rlabel metal2 20328 22736 20328 22736 0 net124
rlabel metal2 17080 27328 17080 27328 0 net125
rlabel metal2 22456 28672 22456 28672 0 net126
rlabel metal2 19880 27496 19880 27496 0 net127
rlabel metal3 10360 31640 10360 31640 0 net128
rlabel metal2 38696 27888 38696 27888 0 net129
rlabel metal2 19992 62888 19992 62888 0 net13
rlabel metal2 13552 27944 13552 27944 0 net130
rlabel metal2 9912 26544 9912 26544 0 net131
rlabel metal3 11592 26936 11592 26936 0 net132
rlabel metal2 20216 25816 20216 25816 0 net133
rlabel metal2 13888 23800 13888 23800 0 net134
rlabel metal2 38584 31248 38584 31248 0 net135
rlabel metal2 10248 22008 10248 22008 0 net136
rlabel metal2 13944 19432 13944 19432 0 net137
rlabel metal2 13608 24192 13608 24192 0 net138
rlabel metal2 17640 32816 17640 32816 0 net139
rlabel metal3 1960 24024 1960 24024 0 net14
rlabel metal2 2296 21672 2296 21672 0 net15
rlabel metal2 1960 50288 1960 50288 0 net16
rlabel metal2 2240 70840 2240 70840 0 net17
rlabel metal2 2912 47432 2912 47432 0 net18
rlabel metal3 1960 66248 1960 66248 0 net19
rlabel metal3 8064 3416 8064 3416 0 net2
rlabel metal3 2184 45304 2184 45304 0 net20
rlabel metal2 16016 41832 16016 41832 0 net21
rlabel metal2 2744 34832 2744 34832 0 net22
rlabel metal2 1960 49896 1960 49896 0 net23
rlabel metal2 21336 40936 21336 40936 0 net24
rlabel metal2 21000 40040 21000 40040 0 net25
rlabel metal3 31192 3360 31192 3360 0 net26
rlabel metal2 11368 3808 11368 3808 0 net27
rlabel metal2 19376 3416 19376 3416 0 net28
rlabel metal2 45528 75152 45528 75152 0 net29
rlabel metal4 22456 40432 22456 40432 0 net3
rlabel metal2 22792 74312 22792 74312 0 net30
rlabel metal3 37016 72016 37016 72016 0 net31
rlabel metal2 20216 74816 20216 74816 0 net32
rlabel metal2 38360 76104 38360 76104 0 net33
rlabel metal2 36568 74760 36568 74760 0 net34
rlabel metal2 34328 74424 34328 74424 0 net35
rlabel metal2 33992 74200 33992 74200 0 net36
rlabel metal2 3304 74872 3304 74872 0 net37
rlabel metal2 18984 4144 18984 4144 0 net38
rlabel metal3 45752 41944 45752 41944 0 net39
rlabel metal2 23576 40040 23576 40040 0 net4
rlabel metal2 47264 41160 47264 41160 0 net40
rlabel metal2 45976 46312 45976 46312 0 net41
rlabel metal2 46648 47376 46648 47376 0 net42
rlabel metal3 46256 49000 46256 49000 0 net43
rlabel metal3 30212 4536 30212 4536 0 net44
rlabel metal2 19208 56112 19208 56112 0 net45
rlabel metal3 24472 56168 24472 56168 0 net46
rlabel metal3 25368 53424 25368 53424 0 net47
rlabel metal2 46984 58072 46984 58072 0 net48
rlabel metal2 26824 51464 26824 51464 0 net49
rlabel metal2 15064 3752 15064 3752 0 net5
rlabel metal2 46984 9856 46984 9856 0 net50
rlabel metal2 28448 12152 28448 12152 0 net51
rlabel metal3 35000 14784 35000 14784 0 net52
rlabel metal2 47432 16408 47432 16408 0 net53
rlabel metal2 47264 19208 47264 19208 0 net54
rlabel metal2 46984 21168 46984 21168 0 net55
rlabel metal2 46760 24080 46760 24080 0 net56
rlabel metal2 16856 75600 16856 75600 0 net57
rlabel metal2 13552 74200 13552 74200 0 net58
rlabel metal2 13496 75600 13496 75600 0 net59
rlabel metal3 4200 75656 4200 75656 0 net6
rlabel metal2 12040 75320 12040 75320 0 net60
rlabel metal2 10696 76440 10696 76440 0 net61
rlabel metal2 8792 75600 8792 75600 0 net62
rlabel metal2 7000 74816 7000 74816 0 net63
rlabel metal2 1960 75600 1960 75600 0 net64
rlabel metal2 34776 76104 34776 76104 0 net65
rlabel metal2 32424 75320 32424 75320 0 net66
rlabel metal2 28840 75600 28840 75600 0 net67
rlabel metal3 28224 76440 28224 76440 0 net68
rlabel metal2 26096 74200 26096 74200 0 net69
rlabel metal3 1904 38696 1904 38696 0 net7
rlabel metal2 20664 75208 20664 75208 0 net70
rlabel metal2 20328 75600 20328 75600 0 net71
rlabel metal2 20104 76384 20104 76384 0 net72
rlabel metal3 25368 17640 25368 17640 0 net73
rlabel metal2 2632 39144 2632 39144 0 net74
rlabel metal2 2856 39872 2856 39872 0 net75
rlabel metal3 26600 41944 26600 41944 0 net76
rlabel metal3 25312 39144 25312 39144 0 net77
rlabel metal2 3192 40376 3192 40376 0 net78
rlabel metal2 21448 18200 21448 18200 0 net79
rlabel metal2 14672 43960 14672 43960 0 net8
rlabel metal2 13944 55216 13944 55216 0 net80
rlabel metal2 10472 56560 10472 56560 0 net81
rlabel metal2 1736 53760 1736 53760 0 net82
rlabel metal2 1736 48720 1736 48720 0 net83
rlabel metal2 27832 49392 27832 49392 0 net84
rlabel metal2 28504 54824 28504 54824 0 net85
rlabel metal3 25928 47264 25928 47264 0 net86
rlabel metal2 12488 70280 12488 70280 0 net87
rlabel metal2 14168 71344 14168 71344 0 net88
rlabel metal3 9800 66248 9800 66248 0 net89
rlabel metal2 12320 44968 12320 44968 0 net9
rlabel metal2 10136 60984 10136 60984 0 net90
rlabel metal2 21840 62328 21840 62328 0 net91
rlabel metal2 21616 66248 21616 66248 0 net92
rlabel metal3 19992 67144 19992 67144 0 net93
rlabel metal2 18312 65296 18312 65296 0 net94
rlabel metal3 6272 51912 6272 51912 0 net95
rlabel metal2 3248 46312 3248 46312 0 net96
rlabel metal2 48216 26544 48216 26544 0 net97
rlabel metal3 48216 28616 48216 28616 0 net98
rlabel metal2 48216 31360 48216 31360 0 net99
rlabel metal2 7056 56840 7056 56840 0 t_reg\[0\]
rlabel metal3 5936 58408 5936 58408 0 t_reg\[1\]
rlabel metal2 4872 55776 4872 55776 0 t_reg\[2\]
rlabel metal2 4480 53816 4480 53816 0 t_reg\[3\]
rlabel metal3 6328 44072 6328 44072 0 t_reg\[4\]
rlabel metal2 7336 37968 7336 37968 0 t_reg\[5\]
rlabel metal2 6720 34776 6720 34776 0 t_reg\[6\]
rlabel metal3 5320 33208 5320 33208 0 t_reg\[7\]
rlabel metal2 8568 26516 8568 26516 0 t_reg\[8\]
rlabel metal2 7784 21448 7784 21448 0 t_reg\[9\]
rlabel metal2 2744 2086 2744 2086 0 wb_clk_i
rlabel metal2 6776 2086 6776 2086 0 wb_rst_i
rlabel metal2 47096 2058 47096 2058 0 wbs_ack_o
rlabel metal2 39200 2184 39200 2184 0 wbs_adr_i[2]
rlabel metal2 43064 2058 43064 2058 0 wbs_adr_i[3]
rlabel metal2 14840 2086 14840 2086 0 wbs_cyc_i
rlabel metal2 2632 76832 2632 76832 0 wbs_dat_i[0]
rlabel metal3 1246 38584 1246 38584 0 wbs_dat_i[16]
rlabel metal2 1736 36176 1736 36176 0 wbs_dat_i[17]
rlabel metal2 1736 33880 1736 33880 0 wbs_dat_i[18]
rlabel metal2 1960 30240 1960 30240 0 wbs_dat_i[19]
rlabel metal3 1246 75544 1246 75544 0 wbs_dat_i[1]
rlabel metal2 1736 29232 1736 29232 0 wbs_dat_i[20]
rlabel metal3 1246 26264 1246 26264 0 wbs_dat_i[21]
rlabel metal3 1246 23800 1246 23800 0 wbs_dat_i[22]
rlabel metal2 1736 21448 1736 21448 0 wbs_dat_i[23]
rlabel metal2 1736 73192 1736 73192 0 wbs_dat_i[2]
rlabel metal2 1736 70672 1736 70672 0 wbs_dat_i[3]
rlabel metal2 1848 68040 1848 68040 0 wbs_dat_i[4]
rlabel metal3 1302 65688 1302 65688 0 wbs_dat_i[5]
rlabel metal3 1302 63224 1302 63224 0 wbs_dat_i[6]
rlabel metal3 1246 60760 1246 60760 0 wbs_dat_i[7]
rlabel metal3 1246 58296 1246 58296 0 wbs_dat_i[8]
rlabel metal2 1736 55944 1736 55944 0 wbs_dat_i[9]
rlabel metal3 48538 1624 48538 1624 0 wbs_dat_o[0]
rlabel metal3 48706 41048 48706 41048 0 wbs_dat_o[16]
rlabel metal3 48538 43512 48538 43512 0 wbs_dat_o[17]
rlabel metal2 48104 46256 48104 46256 0 wbs_dat_o[18]
rlabel metal3 48538 48440 48538 48440 0 wbs_dat_o[19]
rlabel metal2 48104 4144 48104 4144 0 wbs_dat_o[1]
rlabel metal2 48104 51072 48104 51072 0 wbs_dat_o[20]
rlabel metal3 48706 53368 48706 53368 0 wbs_dat_o[21]
rlabel metal2 48104 55888 48104 55888 0 wbs_dat_o[22]
rlabel metal3 48706 58296 48706 58296 0 wbs_dat_o[23]
rlabel metal3 48706 6552 48706 6552 0 wbs_dat_o[2]
rlabel metal3 48706 9016 48706 9016 0 wbs_dat_o[3]
rlabel metal2 47768 11704 47768 11704 0 wbs_dat_o[4]
rlabel metal3 48706 13944 48706 13944 0 wbs_dat_o[5]
rlabel metal2 47768 16632 47768 16632 0 wbs_dat_o[6]
rlabel metal3 48706 18872 48706 18872 0 wbs_dat_o[7]
rlabel metal2 48104 21392 48104 21392 0 wbs_dat_o[8]
rlabel metal3 48706 23800 48706 23800 0 wbs_dat_o[9]
rlabel metal2 23128 2184 23128 2184 0 wbs_sel_i[0]
rlabel metal2 27384 2856 27384 2856 0 wbs_sel_i[1]
rlabel metal2 30968 2086 30968 2086 0 wbs_sel_i[2]
rlabel metal2 10808 2086 10808 2086 0 wbs_stb_i
rlabel metal2 18984 3416 18984 3416 0 wbs_we_i
rlabel metal2 17976 76776 17976 76776 0 x_end[0]
rlabel metal2 15624 76776 15624 76776 0 x_end[1]
rlabel metal2 13944 76496 13944 76496 0 x_end[2]
rlabel metal2 11648 76664 11648 76664 0 x_end[3]
rlabel metal2 10248 76944 10248 76944 0 x_end[4]
rlabel metal2 7896 77882 7896 77882 0 x_end[5]
rlabel metal2 6160 76328 6160 76328 0 x_end[6]
rlabel metal2 4368 76328 4368 76328 0 x_end[7]
rlabel metal2 31192 77938 31192 77938 0 x_start[0]
rlabel metal2 30408 76944 30408 76944 0 x_start[1]
rlabel metal2 29288 76496 29288 76496 0 x_start[2]
rlabel metal2 26376 76776 26376 76776 0 x_start[3]
rlabel metal2 24472 76608 24472 76608 0 x_start[4]
rlabel metal2 23128 76664 23128 76664 0 x_start[5]
rlabel metal2 21560 76832 21560 76832 0 x_start[6]
rlabel metal2 19208 76776 19208 76776 0 x_start[7]
rlabel metal2 46088 76832 46088 76832 0 y[0]
rlabel metal2 44296 76832 44296 76832 0 y[1]
rlabel metal2 42392 76832 42392 76832 0 y[2]
rlabel metal2 40824 76496 40824 76496 0 y[3]
rlabel metal2 38808 76720 38808 76720 0 y[4]
rlabel metal2 36960 76440 36960 76440 0 y[5]
rlabel metal2 35112 76888 35112 76888 0 y[6]
rlabel metal2 33320 75712 33320 75712 0 y[7]
<< properties >>
string FIXED_BBOX 0 0 50000 80000
<< end >>
