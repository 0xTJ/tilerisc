// This is the unpowered netlist.
module interp_tri (active,
    clk,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i,
    x_end,
    x_start,
    y);
 output active;
 input clk;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [3:2] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;
 output [7:0] x_end;
 output [7:0] x_start;
 input [7:0] y;

 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire \a[0][0] ;
 wire \a[0][1] ;
 wire \a[0][2] ;
 wire \a[0][3] ;
 wire \a[0][4] ;
 wire \a[0][5] ;
 wire \a[0][6] ;
 wire \a[0][7] ;
 wire \a[1][0] ;
 wire \a[1][1] ;
 wire \a[1][2] ;
 wire \a[1][3] ;
 wire \a[1][4] ;
 wire \a[1][5] ;
 wire \a[1][6] ;
 wire \a[1][7] ;
 wire \b[0][0] ;
 wire \b[0][1] ;
 wire \b[0][2] ;
 wire \b[0][3] ;
 wire \b[0][4] ;
 wire \b[0][5] ;
 wire \b[0][6] ;
 wire \b[0][7] ;
 wire \b[1][0] ;
 wire \b[1][1] ;
 wire \b[1][2] ;
 wire \b[1][3] ;
 wire \b[1][4] ;
 wire \b[1][5] ;
 wire \b[1][6] ;
 wire \b[1][7] ;
 wire bflip;
 wire \c[0][0] ;
 wire \c[0][1] ;
 wire \c[0][2] ;
 wire \c[0][3] ;
 wire \c[0][4] ;
 wire \c[0][5] ;
 wire \c[0][6] ;
 wire \c[0][7] ;
 wire \c[1][0] ;
 wire \c[1][1] ;
 wire \c[1][2] ;
 wire \c[1][3] ;
 wire \c[1][4] ;
 wire \c[1][5] ;
 wire \c[1][6] ;
 wire \c[1][7] ;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \delta_t[0] ;
 wire \delta_t[1] ;
 wire \delta_t[2] ;
 wire \delta_t[3] ;
 wire \delta_t[4] ;
 wire \delta_t[5] ;
 wire \delta_t[6] ;
 wire \delta_t[7] ;
 wire \delta_t[8] ;
 wire \delta_t[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire \t_reg[0] ;
 wire \t_reg[1] ;
 wire \t_reg[2] ;
 wire \t_reg[3] ;
 wire \t_reg[4] ;
 wire \t_reg[5] ;
 wire \t_reg[6] ;
 wire \t_reg[7] ;
 wire \t_reg[8] ;
 wire \t_reg[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A1 (.I(\a[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__A1 (.I(\a[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1468__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(\a[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__A1 (.I(\a[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A1 (.I(\a[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__I (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A1 (.I(\b[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__I (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1496__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__I (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__I (.I(\b[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__B2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__I (.I(\b[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__B2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__B2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__I (.I(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__I (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__B2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__C2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__I (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__I (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__I (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__I (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__B2 (.I(\delta_t[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__I (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__I (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__I (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__B (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__B2 (.I(\delta_t[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__I (.I(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__I0 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__I1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__I2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__I3 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__S0 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__S1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__I0 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__I1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__I2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__I3 (.I(\delta_t[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__S0 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__S1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__I0 (.I(\a[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__I1 (.I(\b[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__I3 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__S0 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__S1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__I (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__I (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(\a[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(\a[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A1 (.I(\a[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(\a[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__B2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__B2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__B2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A4 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A3 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A4 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A1 (.I(\delta_t[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A1 (.I(\delta_t[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A1 (.I(\delta_t[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A4 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__I (.I(\delta_t[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__I (.I(\delta_t[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A3 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__I (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__B1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A3 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A4 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__B2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A1 (.I(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(\delta_t[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A3 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__I (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__I (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A1 (.I(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__B2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A1 (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__I (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A1 (.I(\b[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A1 (.I(\b[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A1 (.I(\b[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(\b[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A1 (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__I (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__I (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__I (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__I (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__B (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A1 (.I(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__I (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__I (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A3 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__I (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A3 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__I (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A2 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A3 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A3 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A3 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__I (.I(\delta_t[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(\delta_t[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A3 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__I (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A3 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A3 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__B (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A3 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__B (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__I (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__B (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A3 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__B (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__I0 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__I1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__I (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__C (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__C (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__I (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__I (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__I (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__I (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__C (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__C (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__C (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__C (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__B (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__C (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__C (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__B (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__B (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A1 (.I(\a[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__B (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(\a[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(\a[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__A1 (.I(\a[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(\a[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__I (.I(\b[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__C (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__C (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__C (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__C (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__C (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__C (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__B (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__B (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__B (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__B (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__B (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__D (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__CLK (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__CLK (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__D (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__D (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__D (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(wbs_sel_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(wbs_sel_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(wbs_sel_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(y[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(y[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(y[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(y[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(y[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(y[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(y[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(y[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(wbs_adr_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(wbs_adr_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer6_I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_248 ();
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1463_ (.A1(net27),
    .A2(net5),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1464_ (.I(_0699_),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1465_ (.I(net37),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1466_ (.I(bflip),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1467_ (.A1(\a[1][2] ),
    .A2(net31),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1468_ (.A1(\a[1][1] ),
    .A2(net30),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1469_ (.A1(\a[1][5] ),
    .A2(net34),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1470_ (.A1(\a[1][6] ),
    .A2(net35),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1471_ (.A1(_0702_),
    .A2(_0703_),
    .A3(_0704_),
    .A4(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1472_ (.A1(\a[1][0] ),
    .A2(net29),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1473_ (.A1(\a[1][4] ),
    .A2(net33),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1474_ (.A1(\a[1][7] ),
    .A2(net36),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1475_ (.A1(\a[1][3] ),
    .A2(net32),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1476_ (.A1(_0707_),
    .A2(_0708_),
    .A3(_0709_),
    .A4(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1477_ (.A1(_0701_),
    .A2(_0706_),
    .A3(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1478_ (.I(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1479_ (.A1(\b[1][2] ),
    .A2(net31),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1480_ (.A1(\b[1][1] ),
    .A2(net30),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1481_ (.A1(\b[1][5] ),
    .A2(net34),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1482_ (.A1(\b[1][6] ),
    .A2(net35),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1483_ (.A1(_0714_),
    .A2(_0715_),
    .A3(_0716_),
    .A4(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1484_ (.A1(\b[1][0] ),
    .A2(net29),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1485_ (.A1(\b[1][4] ),
    .A2(net33),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1486_ (.A1(\b[1][7] ),
    .A2(net36),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1487_ (.A1(\b[1][3] ),
    .A2(net32),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1488_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0721_),
    .A4(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1489_ (.A1(_0701_),
    .A2(_0718_),
    .A3(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1490_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1491_ (.A1(_0713_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1492_ (.I(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1493_ (.I(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1494_ (.I(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1495_ (.I(_0701_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1496_ (.A1(_0730_),
    .A2(_0718_),
    .A3(_0723_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1497_ (.A1(_0730_),
    .A2(_0706_),
    .A3(_0711_),
    .B(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1498_ (.A1(_0700_),
    .A2(_0729_),
    .B(_0732_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1499_ (.I(\a[0][0] ),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1500_ (.I(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1501_ (.I(net4),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1502_ (.I(net3),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1503_ (.A1(_0735_),
    .A2(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1504_ (.I(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1505_ (.I(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1506_ (.I(\b[0][0] ),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1507_ (.I(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1508_ (.I(_0741_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1509_ (.I(_0742_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1510_ (.I(net3),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1511_ (.A1(net4),
    .A2(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1512_ (.I(_0745_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1513_ (.I(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1514_ (.A1(_0743_),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1515_ (.I(\c[0][0] ),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1516_ (.I(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1517_ (.I(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1518_ (.I(_0744_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1519_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1520_ (.A1(net4),
    .A2(net3),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1521_ (.I(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1522_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1523_ (.I(\delta_t[0] ),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1524_ (.A1(_0751_),
    .A2(_0753_),
    .B1(_0756_),
    .B2(_0757_),
    .C(_0737_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1525_ (.A1(_0734_),
    .A2(_0739_),
    .B1(_0748_),
    .B2(_0758_),
    .ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1526_ (.I(\a[0][1] ),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1527_ (.I(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1528_ (.I(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1529_ (.I(\b[0][1] ),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1530_ (.I(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1531_ (.I(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1532_ (.A1(_0764_),
    .A2(_0747_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1533_ (.I(\c[0][1] ),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1534_ (.I(_0766_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1535_ (.I(_0767_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1536_ (.I(\delta_t[1] ),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1537_ (.A1(_0768_),
    .A2(_0753_),
    .B1(_0756_),
    .B2(_0769_),
    .C(_0737_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1538_ (.A1(_0761_),
    .A2(_0739_),
    .B1(_0765_),
    .B2(_0770_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1539_ (.I(\c[0][2] ),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1540_ (.I(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1541_ (.I(_0752_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1542_ (.I(\b[0][2] ),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1543_ (.I(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1544_ (.I(_0775_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1545_ (.I(\delta_t[2] ),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1546_ (.A1(_0772_),
    .A2(_0773_),
    .B1(_0746_),
    .B2(_0776_),
    .C1(_0755_),
    .C2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1547_ (.I(\a[0][2] ),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1548_ (.I(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1549_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1550_ (.I(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1551_ (.A1(_0782_),
    .A2(_0738_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1552_ (.A1(_0739_),
    .A2(_0778_),
    .B(_0783_),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1553_ (.I(\c[0][3] ),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1554_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1555_ (.I(\b[0][3] ),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1556_ (.I(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1557_ (.I(\delta_t[3] ),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1558_ (.A1(_0785_),
    .A2(_0773_),
    .B1(_0746_),
    .B2(_0787_),
    .C1(_0755_),
    .C2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1559_ (.I(\a[0][3] ),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1560_ (.I(_0790_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1561_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1562_ (.A1(_0792_),
    .A2(_0738_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1563_ (.A1(_0738_),
    .A2(_0789_),
    .B(_0793_),
    .ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1564_ (.I(\a[0][4] ),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1565_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1566_ (.I(_0795_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _1567_ (.I(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1568_ (.I(\b[0][4] ),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1569_ (.I(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1570_ (.A1(_0799_),
    .A2(_0747_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1571_ (.I(\c[0][4] ),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1572_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1573_ (.A1(_0802_),
    .A2(_0753_),
    .B1(_0756_),
    .B2(\delta_t[4] ),
    .C(_0737_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1574_ (.A1(_0797_),
    .A2(_0739_),
    .B1(_0800_),
    .B2(_0803_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1575_ (.I(\a[0][5] ),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1576_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1577_ (.A1(net4),
    .A2(net3),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1578_ (.I(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1579_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1580_ (.A1(_0805_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1581_ (.I(\b[0][5] ),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1582_ (.I(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1583_ (.I(\c[0][5] ),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1584_ (.I(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1585_ (.I(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1586_ (.I(_0735_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1587_ (.I(_0736_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1588_ (.A1(_0814_),
    .A2(_0815_),
    .B(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1589_ (.A1(_0811_),
    .A2(_0747_),
    .B1(_0756_),
    .B2(\delta_t[5] ),
    .C(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1590_ (.A1(_0809_),
    .A2(_0818_),
    .ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1591_ (.I(\a[0][6] ),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1592_ (.I(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1593_ (.I(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1594_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1595_ (.I(\b[0][6] ),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1596_ (.I(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1597_ (.I(\c[0][6] ),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1598_ (.I(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1599_ (.I(\delta_t[6] ),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1600_ (.I(_0735_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1601_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _1602_ (.I0(_0822_),
    .I1(_0824_),
    .I2(_0826_),
    .I3(_0827_),
    .S0(_0816_),
    .S1(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1603_ (.I(_0830_),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1604_ (.I(\a[0][7] ),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1605_ (.I(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1606_ (.I(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1607_ (.I(\b[0][7] ),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1608_ (.I(\c[0][7] ),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _1609_ (.I0(_0833_),
    .I1(_0834_),
    .I2(_0835_),
    .I3(\delta_t[7] ),
    .S0(_0816_),
    .S1(_0815_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1610_ (.I(_0836_),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1611_ (.I(\delta_t[8] ),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1612_ (.A1(_0828_),
    .A2(_0736_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1613_ (.A1(_0837_),
    .A2(_0838_),
    .ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1614_ (.I(\delta_t[9] ),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1615_ (.A1(_0839_),
    .A2(_0838_),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _1616_ (.I0(\a[1][0] ),
    .I1(\b[1][0] ),
    .I2(\c[1][0] ),
    .I3(_0701_),
    .S0(_0816_),
    .S1(_0815_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1617_ (.I(_0840_),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1618_ (.I(\b[1][1] ),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1619_ (.I(_0736_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1620_ (.I(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1621_ (.A1(\c[1][1] ),
    .A2(_0753_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1622_ (.I(_0815_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1623_ (.A1(\a[1][1] ),
    .A2(_0808_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1624_ (.A1(_0841_),
    .A2(_0843_),
    .B1(_0844_),
    .B2(_0845_),
    .C(_0846_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1625_ (.I(\b[1][2] ),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1626_ (.I(_0752_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1627_ (.A1(\c[1][2] ),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1628_ (.A1(\a[1][2] ),
    .A2(_0808_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1629_ (.A1(_0847_),
    .A2(_0843_),
    .B1(_0849_),
    .B2(_0845_),
    .C(_0850_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1630_ (.I(\b[1][3] ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1631_ (.A1(\c[1][3] ),
    .A2(_0848_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1632_ (.A1(\a[1][3] ),
    .A2(_0808_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1633_ (.A1(_0851_),
    .A2(_0843_),
    .B1(_0852_),
    .B2(_0845_),
    .C(_0853_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1634_ (.I(\b[1][4] ),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1635_ (.A1(\c[1][4] ),
    .A2(_0848_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1636_ (.I(_0807_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1637_ (.A1(\a[1][4] ),
    .A2(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1638_ (.A1(_0854_),
    .A2(_0843_),
    .B1(_0855_),
    .B2(_0845_),
    .C(_0857_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1639_ (.I(\b[1][5] ),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1640_ (.A1(\c[1][5] ),
    .A2(_0848_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1641_ (.A1(\a[1][5] ),
    .A2(_0856_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1642_ (.A1(_0858_),
    .A2(_0842_),
    .B1(_0859_),
    .B2(_0829_),
    .C(_0860_),
    .ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1643_ (.I(\b[1][6] ),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1644_ (.A1(\c[1][6] ),
    .A2(_0773_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1645_ (.A1(\a[1][6] ),
    .A2(_0856_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1646_ (.A1(_0861_),
    .A2(_0842_),
    .B1(_0862_),
    .B2(_0829_),
    .C(_0863_),
    .ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1647_ (.I(\b[1][7] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1648_ (.A1(\c[1][7] ),
    .A2(_0773_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1649_ (.A1(\a[1][7] ),
    .A2(_0856_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1650_ (.A1(_0864_),
    .A2(_0842_),
    .B1(_0865_),
    .B2(_0829_),
    .C(_0866_),
    .ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1651_ (.I(\a[0][0] ),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1652_ (.I(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1653_ (.I(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _1654_ (.A1(bflip),
    .A2(_0706_),
    .A3(_0711_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1655_ (.I(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1656_ (.A1(bflip),
    .A2(_0718_),
    .A3(_0723_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1657_ (.I(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1658_ (.A1(_0827_),
    .A2(\t_reg[5] ),
    .A3(_0871_),
    .A4(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1659_ (.I(\t_reg[5] ),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1660_ (.I(\delta_t[6] ),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1661_ (.A1(_0875_),
    .A2(_0712_),
    .A3(_0724_),
    .B(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1662_ (.A1(_0874_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1663_ (.I(\delta_t[2] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1664_ (.I(\t_reg[1] ),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1665_ (.A1(_0879_),
    .A2(_0880_),
    .A3(_0713_),
    .A4(_0725_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _1666_ (.A1(\delta_t[1] ),
    .A2(\t_reg[0] ),
    .A3(_0871_),
    .A4(_0873_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _1667_ (.I(_0870_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1668_ (.I(_0872_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _1669_ (.A1(\t_reg[2] ),
    .A2(_0883_),
    .A3(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1670_ (.A1(_0880_),
    .A2(_0713_),
    .A3(_0725_),
    .B(_0879_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1671_ (.A1(_0881_),
    .A2(_0882_),
    .B1(_0885_),
    .B2(\delta_t[3] ),
    .C(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _1672_ (.A1(\t_reg[3] ),
    .A2(_0883_),
    .A3(_0884_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1673_ (.I(_0885_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1674_ (.A1(\delta_t[4] ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\delta_t[3] ),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1675_ (.I(_0888_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1676_ (.A1(\delta_t[4] ),
    .A2(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1677_ (.A1(_0887_),
    .A2(_0890_),
    .B(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1678_ (.A1(\delta_t[5] ),
    .A2(\t_reg[4] ),
    .A3(_0871_),
    .A4(_0873_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1679_ (.I(\t_reg[4] ),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1680_ (.I(\delta_t[5] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1681_ (.A1(_0895_),
    .A2(_0713_),
    .A3(_0725_),
    .B(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1682_ (.A1(_0894_),
    .A2(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1683_ (.I(_0896_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1684_ (.A1(\t_reg[4] ),
    .A2(_0726_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1685_ (.A1(_0899_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1686_ (.A1(_0893_),
    .A2(_0898_),
    .B(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1687_ (.A1(_0878_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1688_ (.I(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1689_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1690_ (.I(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(_0869_),
    .A2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1692_ (.I(_0759_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1693_ (.I(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1694_ (.I(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1695_ (.A1(_0893_),
    .A2(_0898_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1696_ (.I(_0911_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1697_ (.I(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1698_ (.A1(_0910_),
    .A2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1699_ (.A1(_0907_),
    .A2(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1700_ (.A1(_0780_),
    .A2(_0912_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1701_ (.A1(_0874_),
    .A2(_0894_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1702_ (.A1(_0877_),
    .A2(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1703_ (.A1(_0874_),
    .A2(_0877_),
    .A3(_0894_),
    .A4(_0897_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1704_ (.A1(_0887_),
    .A2(_0890_),
    .B(_0919_),
    .C(_0892_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1705_ (.I(\delta_t[7] ),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1706_ (.A1(\t_reg[6] ),
    .A2(_0883_),
    .A3(_0884_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1707_ (.A1(_0922_),
    .A2(_0921_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1708_ (.A1(_0918_),
    .A2(_0920_),
    .B(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1709_ (.A1(_0923_),
    .A2(_0918_),
    .A3(_0920_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1710_ (.A1(_0925_),
    .A2(net118),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1711_ (.I(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1712_ (.I(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1713_ (.A1(_0869_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1714_ (.A1(_0909_),
    .A2(_0905_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1715_ (.A1(_0916_),
    .A2(_0929_),
    .A3(_0930_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1716_ (.A1(_0915_),
    .A2(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1717_ (.I(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1718_ (.I(_0913_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1719_ (.I(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1720_ (.A1(_0774_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1721_ (.I(_0906_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_0763_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1723_ (.I(_0928_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1724_ (.I(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1725_ (.I(_0940_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1726_ (.A1(_0741_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1727_ (.A1(_0936_),
    .A2(_0938_),
    .A3(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1728_ (.I(_0934_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1729_ (.I(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1730_ (.I(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1731_ (.I(_0937_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1732_ (.I(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1733_ (.A1(_0742_),
    .A2(_0948_),
    .B1(_0945_),
    .B2(_0764_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1734_ (.I(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1735_ (.A1(_0742_),
    .A2(_0946_),
    .A3(_0938_),
    .A4(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1736_ (.I(_0948_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1737_ (.A1(_0764_),
    .A2(_0742_),
    .A3(_0952_),
    .A4(_0945_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1738_ (.A1(_0951_),
    .A2(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1739_ (.A1(_0943_),
    .A2(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1740_ (.A1(_0933_),
    .A2(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1741_ (.A1(_0943_),
    .A2(_0951_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1742_ (.A1(_0915_),
    .A2(_0931_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1743_ (.A1(_0791_),
    .A2(_0913_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1744_ (.A1(_0909_),
    .A2(_0905_),
    .B1(_0928_),
    .B2(_0869_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1745_ (.A1(_0909_),
    .A2(_0868_),
    .A3(_0904_),
    .A4(_0928_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1746_ (.A1(_0916_),
    .A2(_0960_),
    .B(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1747_ (.A1(\a[0][2] ),
    .A2(_0903_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1748_ (.A1(\delta_t[7] ),
    .A2(\t_reg[6] ),
    .A3(_0727_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1749_ (.A1(\t_reg[7] ),
    .A2(_0883_),
    .A3(_0884_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1750_ (.A1(_0965_),
    .A2(_0837_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1751_ (.A1(_0964_),
    .A2(_0924_),
    .A3(net128),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1752_ (.A1(_0964_),
    .A2(_0924_),
    .B(net121),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1753_ (.I(_0867_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1754_ (.A1(_0967_),
    .A2(_0968_),
    .B(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1755_ (.A1(_0908_),
    .A2(_0927_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1756_ (.A1(_0963_),
    .A2(_0970_),
    .A3(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1757_ (.A1(_0959_),
    .A2(_0962_),
    .A3(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1758_ (.A1(_0958_),
    .A2(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1759_ (.A1(_0943_),
    .A2(_0953_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1760_ (.A1(_0786_),
    .A2(_0944_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1761_ (.A1(_0938_),
    .A2(_0942_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1762_ (.A1(_0938_),
    .A2(_0942_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1763_ (.A1(_0936_),
    .A2(_0977_),
    .B(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1764_ (.I(_0906_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1765_ (.A1(\b[0][2] ),
    .A2(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1766_ (.A1(_0967_),
    .A2(_0968_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1767_ (.I(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1768_ (.I(_0983_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1769_ (.I(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1770_ (.I(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1771_ (.A1(_0740_),
    .A2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1772_ (.A1(_0763_),
    .A2(_0941_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1773_ (.A1(_0981_),
    .A2(_0987_),
    .A3(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1774_ (.A1(_0976_),
    .A2(_0979_),
    .A3(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1775_ (.A1(_0974_),
    .A2(_0975_),
    .A3(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1776_ (.A1(_0956_),
    .A2(_0957_),
    .A3(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1777_ (.I(_0946_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1778_ (.A1(_0743_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(_0949_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1780_ (.A1(_0907_),
    .A2(_0914_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1781_ (.I(_0869_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1782_ (.A1(_0743_),
    .A2(_0997_),
    .B(_0993_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1783_ (.A1(_0951_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1784_ (.A1(_0996_),
    .A2(_0998_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1785_ (.A1(_0933_),
    .A2(_0955_),
    .B(_0999_),
    .C(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1786_ (.A1(_0933_),
    .A2(_0955_),
    .B(_0992_),
    .C(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1787_ (.A1(_0956_),
    .A2(_0957_),
    .B(_0991_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1788_ (.A1(_0958_),
    .A2(_0973_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1789_ (.A1(_0790_),
    .A2(_0903_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1790_ (.A1(_0795_),
    .A2(_0911_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1791_ (.A1(_1005_),
    .A2(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1792_ (.A1(_0970_),
    .A2(_0971_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1793_ (.A1(_0970_),
    .A2(_0971_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1794_ (.A1(_0963_),
    .A2(_1008_),
    .B(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1795_ (.A1(\a[0][2] ),
    .A2(_0926_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1796_ (.A1(_0759_),
    .A2(_0982_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1797_ (.A1(_0923_),
    .A2(_0966_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _1798_ (.A1(_0878_),
    .A2(_0898_),
    .A3(_0923_),
    .A4(_0966_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1799_ (.I(_0965_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1800_ (.A1(\delta_t[8] ),
    .A2(\t_reg[7] ),
    .B(\t_reg[6] ),
    .C(_0726_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1801_ (.A1(_0837_),
    .A2(_1015_),
    .B1(_1016_),
    .B2(_0921_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1802_ (.A1(_0918_),
    .A2(_1013_),
    .B1(_1014_),
    .B2(_0893_),
    .C(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1803_ (.A1(\t_reg[8] ),
    .A2(_0871_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1804_ (.A1(_0873_),
    .A2(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1805_ (.A1(_0839_),
    .A2(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1806_ (.A1(_1018_),
    .A2(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1807_ (.I(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1808_ (.A1(_0868_),
    .A2(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1809_ (.A1(_1011_),
    .A2(_1012_),
    .A3(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1810_ (.A1(_1007_),
    .A2(_1010_),
    .A3(net120),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1811_ (.A1(_0962_),
    .A2(_0972_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1812_ (.A1(_0962_),
    .A2(_0972_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1813_ (.A1(_0959_),
    .A2(_1027_),
    .B(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _1814_ (.A1(_1004_),
    .A2(_1026_),
    .A3(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1815_ (.A1(_0979_),
    .A2(_0989_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1816_ (.A1(_0979_),
    .A2(_0989_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1817_ (.A1(_0976_),
    .A2(_1031_),
    .B(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(\b[0][3] ),
    .A2(_0980_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1819_ (.A1(\b[0][4] ),
    .A2(_0934_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1820_ (.A1(_1034_),
    .A2(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1821_ (.I(_0985_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1822_ (.A1(_0762_),
    .A2(_0940_),
    .B1(_1037_),
    .B2(_0740_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1823_ (.A1(_0762_),
    .A2(_0740_),
    .A3(_0940_),
    .A4(_1037_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1824_ (.A1(_0981_),
    .A2(_1038_),
    .B(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1825_ (.A1(\b[0][2] ),
    .A2(_0939_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1826_ (.I(net131),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1827_ (.I(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1828_ (.I(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1829_ (.A1(\b[0][0] ),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1830_ (.A1(\b[0][1] ),
    .A2(_0986_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1831_ (.A1(_1041_),
    .A2(_1045_),
    .A3(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1832_ (.A1(_1040_),
    .A2(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1833_ (.A1(_1036_),
    .A2(_1048_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1834_ (.A1(_1033_),
    .A2(_1049_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1835_ (.I(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1836_ (.A1(_1030_),
    .A2(_1051_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1837_ (.A1(_0975_),
    .A2(_0990_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1838_ (.A1(_0975_),
    .A2(_0990_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1839_ (.A1(_0974_),
    .A2(_1053_),
    .B(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1840_ (.A1(_1052_),
    .A2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1841_ (.A1(_1003_),
    .A2(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1842_ (.A1(_1002_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1843_ (.A1(_0734_),
    .A2(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1844_ (.I(_1003_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1845_ (.A1(_1060_),
    .A2(_1056_),
    .B1(_1057_),
    .B2(_1002_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1846_ (.A1(_1052_),
    .A2(_1055_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1847_ (.A1(_1034_),
    .A2(_1035_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1848_ (.A1(_1026_),
    .A2(_1029_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1849_ (.A1(_1026_),
    .A2(_1029_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1850_ (.A1(_1004_),
    .A2(_1064_),
    .B(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1851_ (.A1(_1005_),
    .A2(_1006_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1852_ (.A1(_1010_),
    .A2(_1025_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1853_ (.A1(_1010_),
    .A2(_1025_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1854_ (.A1(_1007_),
    .A2(_1068_),
    .B(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1855_ (.A1(\a[0][5] ),
    .A2(_0911_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1856_ (.A1(\a[0][4] ),
    .A2(_0903_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1857_ (.A1(\a[0][3] ),
    .A2(_0926_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1858_ (.A1(_1072_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1859_ (.A1(_1071_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1860_ (.I(_0759_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1861_ (.A1(_1076_),
    .A2(_0983_),
    .B1(_1023_),
    .B2(_0969_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1862_ (.A1(_1076_),
    .A2(_0867_),
    .A3(_0983_),
    .A4(net132),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1863_ (.A1(_1011_),
    .A2(_1077_),
    .B(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1864_ (.A1(\a[0][2] ),
    .A2(_0982_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1865_ (.A1(_1022_),
    .A2(\a[0][1] ),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1866_ (.A1(\t_reg[9] ),
    .A2(_0727_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1867_ (.A1(\delta_t[9] ),
    .A2(_1020_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1868_ (.A1(_1018_),
    .A2(_1021_),
    .B(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1869_ (.A1(_1082_),
    .A2(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1870_ (.A1(_0733_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1871_ (.A1(_1080_),
    .A2(_1081_),
    .A3(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1872_ (.A1(_1079_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1873_ (.A1(_1075_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1874_ (.A1(_1067_),
    .A2(_1070_),
    .A3(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1875_ (.A1(_1066_),
    .A2(net112),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1876_ (.A1(_1063_),
    .A2(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1877_ (.A1(_1040_),
    .A2(_1047_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1878_ (.A1(_1036_),
    .A2(_1048_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1879_ (.A1(_1093_),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1880_ (.A1(_1045_),
    .A2(_1046_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1881_ (.A1(_1045_),
    .A2(_1046_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1882_ (.A1(_1041_),
    .A2(_1096_),
    .B(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1883_ (.A1(_0774_),
    .A2(_1037_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1884_ (.A1(\b[0][1] ),
    .A2(_1044_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1885_ (.A1(_1084_),
    .A2(_1082_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1886_ (.I(net136),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1887_ (.I(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1888_ (.A1(\b[0][0] ),
    .A2(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1889_ (.A1(_1100_),
    .A2(_1104_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1890_ (.A1(_1099_),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1891_ (.A1(_1098_),
    .A2(_1106_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1892_ (.A1(\b[0][5] ),
    .A2(_0935_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1893_ (.A1(\b[0][4] ),
    .A2(_0980_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1894_ (.I(_0939_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1895_ (.A1(\b[0][3] ),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1896_ (.A1(_1109_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1897_ (.A1(_1108_),
    .A2(_1112_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1898_ (.A1(_1107_),
    .A2(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1899_ (.A1(_1095_),
    .A2(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1900_ (.A1(_1092_),
    .A2(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1901_ (.A1(_1030_),
    .A2(_1051_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1902_ (.A1(_1033_),
    .A2(_1049_),
    .B(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1903_ (.A1(_1116_),
    .A2(_1118_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1904_ (.A1(_1062_),
    .A2(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1905_ (.A1(_1061_),
    .A2(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1906_ (.A1(_0910_),
    .A2(_1121_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1907_ (.A1(_1059_),
    .A2(_1122_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1908_ (.I(_1123_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1909_ (.A1(_0910_),
    .A2(_1121_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1910_ (.A1(_1059_),
    .A2(_1122_),
    .B(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1911_ (.I(_1116_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1912_ (.A1(_1126_),
    .A2(_1118_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1913_ (.A1(_1062_),
    .A2(_1119_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1914_ (.A1(_1061_),
    .A2(_1120_),
    .B(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1915_ (.I(_1091_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1916_ (.A1(_1063_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1917_ (.A1(_1095_),
    .A2(_1114_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1918_ (.A1(_1092_),
    .A2(_1115_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1919_ (.A1(_1132_),
    .A2(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1920_ (.A1(_1109_),
    .A2(_1111_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1921_ (.A1(_1108_),
    .A2(_1112_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1922_ (.A1(_1135_),
    .A2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1923_ (.A1(_0823_),
    .A2(_0945_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1924_ (.A1(_1004_),
    .A2(_1064_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1925_ (.A1(_1139_),
    .A2(net111),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1926_ (.I(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1927_ (.A1(_1026_),
    .A2(_1029_),
    .A3(_1090_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1928_ (.A1(_1070_),
    .A2(_1089_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1929_ (.A1(_1089_),
    .A2(_1070_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1930_ (.A1(_1067_),
    .A2(_1143_),
    .B(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1931_ (.I(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1932_ (.A1(_1071_),
    .A2(_1074_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1933_ (.A1(_1072_),
    .A2(_1073_),
    .B(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1934_ (.A1(\a[0][6] ),
    .A2(_0912_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1935_ (.A1(_1148_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1936_ (.A1(_1079_),
    .A2(net130),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1937_ (.A1(_1075_),
    .A2(net125),
    .B(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1938_ (.A1(_0804_),
    .A2(_0904_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1939_ (.A1(_0794_),
    .A2(_0926_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1940_ (.A1(\a[0][3] ),
    .A2(_0983_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1941_ (.A1(_1154_),
    .A2(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1942_ (.A1(_1153_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1943_ (.I(_1101_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1944_ (.A1(_0908_),
    .A2(_1023_),
    .B1(_1158_),
    .B2(_0969_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1945_ (.A1(_1076_),
    .A2(_0969_),
    .A3(_1023_),
    .A4(_1158_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1946_ (.A1(_1080_),
    .A2(_1159_),
    .B(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1947_ (.A1(_1076_),
    .A2(_0867_),
    .B(_1158_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1948_ (.A1(_0760_),
    .A2(_0733_),
    .A3(_1085_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1949_ (.A1(_1162_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1950_ (.A1(_0779_),
    .A2(_1042_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1951_ (.A1(_1161_),
    .A2(_1164_),
    .A3(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1952_ (.A1(_1157_),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1953_ (.A1(_1150_),
    .A2(_1152_),
    .A3(net133),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1954_ (.A1(_1142_),
    .A2(_1146_),
    .A3(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _1955_ (.A1(_1138_),
    .A2(_1141_),
    .A3(net129),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1956_ (.A1(_1098_),
    .A2(_1106_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1957_ (.A1(_1107_),
    .A2(_1113_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1958_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1959_ (.I(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1960_ (.A1(_1100_),
    .A2(_1104_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1961_ (.I(_1037_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1962_ (.I(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1963_ (.A1(_0775_),
    .A2(_1177_),
    .A3(_1105_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1964_ (.A1(_1175_),
    .A2(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1965_ (.I(_1103_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1966_ (.A1(_0763_),
    .A2(_0741_),
    .B(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1967_ (.A1(_0762_),
    .A2(_0741_),
    .A3(_1180_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1968_ (.A1(_1181_),
    .A2(_1182_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1969_ (.I(_1044_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1970_ (.A1(_0774_),
    .A2(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1971_ (.A1(_1183_),
    .A2(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1972_ (.A1(_1179_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1973_ (.A1(\b[0][5] ),
    .A2(_0947_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1974_ (.A1(\b[0][4] ),
    .A2(_0941_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1975_ (.A1(_0786_),
    .A2(_1176_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1976_ (.A1(_1189_),
    .A2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1977_ (.A1(_1188_),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1978_ (.A1(_1187_),
    .A2(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1979_ (.A1(_1187_),
    .A2(_1192_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1980_ (.A1(_1193_),
    .A2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1981_ (.A1(_1174_),
    .A2(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1982_ (.A1(_1137_),
    .A2(_1170_),
    .A3(_1196_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1983_ (.A1(_1131_),
    .A2(_1134_),
    .A3(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1984_ (.A1(_1127_),
    .A2(_1129_),
    .A3(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1985_ (.A1(_0781_),
    .A2(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1986_ (.A1(_1125_),
    .A2(_1200_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1987_ (.I(_1201_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1988_ (.A1(_0782_),
    .A2(_1199_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1989_ (.A1(_1125_),
    .A2(_1200_),
    .B(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1990_ (.A1(_1127_),
    .A2(_1198_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1991_ (.A1(_1127_),
    .A2(_1198_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1992_ (.A1(_1129_),
    .A2(_1204_),
    .B(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1993_ (.A1(_1137_),
    .A2(_1170_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1994_ (.A1(_1134_),
    .A2(_1197_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1995_ (.A1(_1134_),
    .A2(_1197_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1996_ (.A1(_1131_),
    .A2(_1208_),
    .B(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1997_ (.A1(_1137_),
    .A2(_1170_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1998_ (.A1(_1174_),
    .A2(_1195_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1999_ (.A1(_1211_),
    .A2(_1196_),
    .B(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2000_ (.A1(_1179_),
    .A2(_1186_),
    .B(_1193_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2001_ (.I(_1182_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2002_ (.A1(_1183_),
    .A2(_1185_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2003_ (.I(_1180_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2004_ (.A1(_0775_),
    .A2(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2005_ (.A1(_1183_),
    .A2(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2006_ (.A1(_0775_),
    .A2(_1215_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2007_ (.A1(_1215_),
    .A2(_1216_),
    .A3(_1219_),
    .B(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2008_ (.I(_1110_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2009_ (.I(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2010_ (.A1(_0798_),
    .A2(_1176_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2011_ (.A1(_0786_),
    .A2(_1184_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2012_ (.A1(_1224_),
    .A2(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2013_ (.A1(_0810_),
    .A2(_1223_),
    .A3(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2014_ (.A1(_0810_),
    .A2(_1223_),
    .B(_1226_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2015_ (.A1(_1227_),
    .A2(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2016_ (.I(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2017_ (.A1(_1221_),
    .A2(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2018_ (.A1(_1214_),
    .A2(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2019_ (.A1(_1140_),
    .A2(net129),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2020_ (.A1(_1138_),
    .A2(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2021_ (.A1(_1189_),
    .A2(_1190_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2022_ (.A1(_1188_),
    .A2(_1191_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2023_ (.A1(_1235_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _2024_ (.I(_1168_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2025_ (.A1(_1146_),
    .A2(_1238_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2026_ (.A1(_1146_),
    .A2(_1238_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2027_ (.A1(_1142_),
    .A2(net119),
    .A3(_1238_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2028_ (.A1(net122),
    .A2(_1239_),
    .A3(_1240_),
    .B1(_1241_),
    .B2(_1140_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2029_ (.I(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2030_ (.A1(_0819_),
    .A2(_0913_),
    .A3(_1148_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2031_ (.A1(_1152_),
    .A2(_1167_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2032_ (.A1(_1152_),
    .A2(_1167_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2033_ (.A1(_1150_),
    .A2(_1245_),
    .B(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2034_ (.A1(_1154_),
    .A2(_1155_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2035_ (.A1(_1153_),
    .A2(_1156_),
    .B(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2036_ (.A1(\a[0][6] ),
    .A2(_0904_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2037_ (.A1(_1249_),
    .A2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2038_ (.A1(_0831_),
    .A2(_0912_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2039_ (.A1(_1251_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2040_ (.I(_1085_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2041_ (.A1(_0761_),
    .A2(_0733_),
    .B(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2042_ (.A1(_0908_),
    .A2(_0868_),
    .A3(_1102_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2043_ (.A1(_0780_),
    .A2(_1043_),
    .A3(_1255_),
    .A4(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2044_ (.I(_1163_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2045_ (.A1(_1162_),
    .A2(_1258_),
    .B(_1165_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2046_ (.A1(net137),
    .A2(_1257_),
    .A3(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2047_ (.A1(_1157_),
    .A2(_1166_),
    .B(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2048_ (.A1(\a[0][5] ),
    .A2(_0927_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2049_ (.A1(_0794_),
    .A2(_0984_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2050_ (.A1(_0790_),
    .A2(_1042_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2051_ (.A1(_1262_),
    .A2(_1263_),
    .A3(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2052_ (.A1(_0779_),
    .A2(_1102_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2053_ (.A1(_1255_),
    .A2(_1256_),
    .A3(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2054_ (.A1(_1255_),
    .A2(_1256_),
    .B(_1266_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2055_ (.A1(_1162_),
    .A2(_1165_),
    .B(_1256_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2056_ (.A1(_0779_),
    .A2(_1258_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2057_ (.A1(_1267_),
    .A2(_1268_),
    .A3(_1269_),
    .B(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2058_ (.A1(_1265_),
    .A2(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2059_ (.A1(_1261_),
    .A2(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2060_ (.A1(_1253_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2061_ (.A1(_1244_),
    .A2(_1247_),
    .A3(_1274_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2062_ (.A1(_1239_),
    .A2(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2063_ (.A1(\b[0][6] ),
    .A2(_0948_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2064_ (.I(_0944_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2065_ (.A1(\b[0][7] ),
    .A2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2066_ (.A1(_1277_),
    .A2(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2067_ (.A1(_1243_),
    .A2(_1276_),
    .A3(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2068_ (.A1(_1234_),
    .A2(_1237_),
    .A3(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2069_ (.A1(_1213_),
    .A2(_1232_),
    .A3(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2070_ (.A1(_1207_),
    .A2(_1210_),
    .A3(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2071_ (.A1(_1206_),
    .A2(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2072_ (.A1(_0791_),
    .A2(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2073_ (.A1(_1203_),
    .A2(_1286_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2074_ (.I(_1287_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2075_ (.A1(_0792_),
    .A2(_1285_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2076_ (.A1(_1203_),
    .A2(_1286_),
    .B(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2077_ (.A1(_1207_),
    .A2(_1283_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2078_ (.A1(_1206_),
    .A2(_1284_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2079_ (.A1(_1210_),
    .A2(_1290_),
    .B(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2080_ (.I(_1232_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2081_ (.A1(_1293_),
    .A2(_1282_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2082_ (.A1(_1137_),
    .A2(_1170_),
    .A3(_1283_),
    .B1(_1294_),
    .B2(_1213_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2083_ (.I(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2084_ (.I(_1237_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2085_ (.A1(_1297_),
    .A2(_1281_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2086_ (.A1(_1297_),
    .A2(_1281_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2087_ (.A1(_1234_),
    .A2(_1298_),
    .B(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2088_ (.A1(_1234_),
    .A2(_1297_),
    .A3(_1281_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2089_ (.A1(_1214_),
    .A2(_1231_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2090_ (.A1(_1293_),
    .A2(_1301_),
    .B(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2091_ (.A1(_1221_),
    .A2(_1230_),
    .B(_1220_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2092_ (.A1(_1181_),
    .A2(_1218_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2093_ (.A1(_1220_),
    .A2(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2094_ (.I(_1177_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2095_ (.A1(_0810_),
    .A2(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2096_ (.I(_1184_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2097_ (.I(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2098_ (.A1(_0798_),
    .A2(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2099_ (.I(_1217_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2100_ (.A1(_0787_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2101_ (.A1(_1308_),
    .A2(_1311_),
    .A3(_1313_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2102_ (.A1(_1306_),
    .A2(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2103_ (.A1(_1304_),
    .A2(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2104_ (.A1(_1243_),
    .A2(_1276_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2105_ (.A1(_1277_),
    .A2(_1279_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2106_ (.A1(_1317_),
    .A2(_1280_),
    .B(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2107_ (.A1(_1224_),
    .A2(_1225_),
    .B(_1227_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2108_ (.A1(_1146_),
    .A2(_1238_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2109_ (.A1(_1321_),
    .A2(_1275_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2110_ (.A1(_1321_),
    .A2(_1275_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2111_ (.A1(_1242_),
    .A2(_1322_),
    .B(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2112_ (.I(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2113_ (.A1(net124),
    .A2(_1274_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2114_ (.A1(_1247_),
    .A2(_1274_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2115_ (.A1(_1244_),
    .A2(_1326_),
    .B(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2116_ (.A1(_0820_),
    .A2(_0947_),
    .A3(_1249_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2117_ (.A1(_0832_),
    .A2(_0935_),
    .A3(_1251_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2118_ (.A1(_1329_),
    .A2(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2119_ (.A1(_1261_),
    .A2(_1272_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2120_ (.A1(_1253_),
    .A2(_1273_),
    .B(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2121_ (.A1(_1265_),
    .A2(_1271_),
    .B(_1270_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2122_ (.A1(_1162_),
    .A2(_1266_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2123_ (.A1(_1270_),
    .A2(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2124_ (.A1(\a[0][5] ),
    .A2(_0984_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2125_ (.A1(_0795_),
    .A2(_1042_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2126_ (.A1(\a[0][3] ),
    .A2(net134),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2127_ (.A1(_1337_),
    .A2(_1338_),
    .A3(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2128_ (.A1(_1336_),
    .A2(_1340_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2129_ (.A1(_1334_),
    .A2(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2130_ (.A1(_1263_),
    .A2(_1264_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2131_ (.A1(_1263_),
    .A2(_1264_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2132_ (.A1(_1262_),
    .A2(_1343_),
    .B(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2133_ (.A1(\a[0][6] ),
    .A2(_0927_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2134_ (.A1(_1345_),
    .A2(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2135_ (.A1(\a[0][7] ),
    .A2(_0905_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2136_ (.A1(_1347_),
    .A2(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2137_ (.A1(_1342_),
    .A2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2138_ (.A1(_1333_),
    .A2(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2139_ (.A1(_1331_),
    .A2(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2140_ (.A1(_1328_),
    .A2(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2141_ (.A1(\b[0][7] ),
    .A2(_0952_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2142_ (.I(_1223_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2143_ (.A1(_0823_),
    .A2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2144_ (.A1(_1354_),
    .A2(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2145_ (.A1(_1325_),
    .A2(_1353_),
    .A3(_1357_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2146_ (.A1(_1319_),
    .A2(_1320_),
    .A3(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2147_ (.A1(_1303_),
    .A2(_1316_),
    .A3(_1359_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2148_ (.A1(_1360_),
    .A2(_1300_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2149_ (.A1(_1296_),
    .A2(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2150_ (.A1(_0797_),
    .A2(_1292_),
    .A3(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2151_ (.A1(_1289_),
    .A2(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2152_ (.I(_1364_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2153_ (.A1(_1292_),
    .A2(_1362_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2154_ (.A1(_0796_),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2155_ (.A1(_1289_),
    .A2(_1363_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2156_ (.A1(_1296_),
    .A2(_1361_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2157_ (.A1(_1292_),
    .A2(_1362_),
    .B(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2158_ (.A1(_1316_),
    .A2(_1359_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2159_ (.A1(_1303_),
    .A2(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2160_ (.A1(_1300_),
    .A2(_1360_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2161_ (.A1(_1371_),
    .A2(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2162_ (.A1(_1325_),
    .A2(_1353_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2163_ (.A1(_1374_),
    .A2(_1357_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2164_ (.A1(_1320_),
    .A2(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2165_ (.A1(_1320_),
    .A2(_1358_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2166_ (.A1(_1319_),
    .A2(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2167_ (.A1(_1376_),
    .A2(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2168_ (.A1(_1304_),
    .A2(_1315_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2169_ (.A1(_1316_),
    .A2(_1359_),
    .B(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2170_ (.A1(_0776_),
    .A2(_1215_),
    .B1(_1305_),
    .B2(_1314_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2171_ (.I(_1313_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2172_ (.A1(_0798_),
    .A2(_0787_),
    .B(_1312_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2173_ (.A1(_0799_),
    .A2(_1383_),
    .B(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2174_ (.A1(_0811_),
    .A2(_1310_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2175_ (.A1(_1385_),
    .A2(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2176_ (.A1(_1306_),
    .A2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2177_ (.A1(_1382_),
    .A2(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2178_ (.A1(_1354_),
    .A2(_1356_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2179_ (.A1(_1354_),
    .A2(_1356_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2180_ (.A1(_1374_),
    .A2(_1390_),
    .B(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2181_ (.A1(_1311_),
    .A2(_1313_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2182_ (.A1(_1311_),
    .A2(_1313_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2183_ (.A1(_1308_),
    .A2(_1393_),
    .B(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2184_ (.A1(_1328_),
    .A2(_1352_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(_1328_),
    .A2(_1352_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2186_ (.A1(_1324_),
    .A2(_1396_),
    .B(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2187_ (.A1(_1333_),
    .A2(_1350_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2188_ (.A1(_1331_),
    .A2(_1351_),
    .B(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2189_ (.A1(_0820_),
    .A2(_1222_),
    .A3(_1345_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2190_ (.A1(_1347_),
    .A2(_1348_),
    .B(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2191_ (.A1(_1334_),
    .A2(_1341_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2192_ (.A1(_1342_),
    .A2(_1349_),
    .B(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2193_ (.A1(_0781_),
    .A2(_1258_),
    .B1(_1335_),
    .B2(_1340_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2194_ (.I(_1339_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2195_ (.A1(_0794_),
    .A2(_0790_),
    .B(_1102_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2196_ (.A1(_0795_),
    .A2(_1406_),
    .B(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2197_ (.A1(_0804_),
    .A2(_1043_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2198_ (.A1(_1408_),
    .A2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2199_ (.A1(_1336_),
    .A2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2200_ (.A1(_1405_),
    .A2(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2201_ (.A1(_1338_),
    .A2(_1339_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2202_ (.A1(_1338_),
    .A2(_1339_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2203_ (.A1(_1337_),
    .A2(_1413_),
    .B(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2204_ (.A1(_0819_),
    .A2(_0984_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2205_ (.A1(_1415_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2206_ (.A1(_0831_),
    .A2(_0939_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2207_ (.A1(_1417_),
    .A2(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2208_ (.A1(_1417_),
    .A2(_1418_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2209_ (.A1(_1419_),
    .A2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2210_ (.A1(_1412_),
    .A2(_1421_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2211_ (.A1(_1404_),
    .A2(_1422_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2212_ (.A1(_1402_),
    .A2(_1423_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2213_ (.A1(_1400_),
    .A2(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2214_ (.A1(\b[0][7] ),
    .A2(_1355_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2215_ (.I(_1307_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2216_ (.A1(_0823_),
    .A2(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2217_ (.A1(_1426_),
    .A2(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2218_ (.A1(_1398_),
    .A2(_1425_),
    .A3(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2219_ (.A1(_1392_),
    .A2(_1395_),
    .A3(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2220_ (.A1(_1381_),
    .A2(_1389_),
    .A3(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2221_ (.A1(_1379_),
    .A2(_1432_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2222_ (.A1(_1373_),
    .A2(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2223_ (.A1(_0805_),
    .A2(_1369_),
    .A3(_1434_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2224_ (.A1(_1366_),
    .A2(_1367_),
    .B(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2225_ (.A1(_1366_),
    .A2(_1367_),
    .A3(_1435_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2226_ (.A1(_1436_),
    .A2(_1437_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2227_ (.A1(_1369_),
    .A2(_1434_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2228_ (.A1(_0805_),
    .A2(_1438_),
    .B(_1436_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2229_ (.A1(_1373_),
    .A2(_1433_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2230_ (.A1(_1373_),
    .A2(_1433_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2231_ (.A1(_1369_),
    .A2(_1440_),
    .B(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2232_ (.A1(_1389_),
    .A2(_1431_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2233_ (.A1(_1389_),
    .A2(_1431_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2234_ (.A1(_1381_),
    .A2(_1443_),
    .A3(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2235_ (.A1(_1379_),
    .A2(_1432_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2236_ (.A1(_1445_),
    .A2(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2237_ (.I(_1395_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2238_ (.A1(_1448_),
    .A2(_1430_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2239_ (.A1(_1448_),
    .A2(_1430_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2240_ (.A1(_1392_),
    .A2(_1449_),
    .B(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2241_ (.A1(_1382_),
    .A2(_1388_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2242_ (.A1(_1452_),
    .A2(_1443_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2243_ (.A1(_1398_),
    .A2(_1425_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2244_ (.A1(_1426_),
    .A2(_1428_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2245_ (.A1(_1454_),
    .A2(_1429_),
    .B(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2246_ (.A1(_0799_),
    .A2(_1383_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2247_ (.A1(_1384_),
    .A2(_1386_),
    .B(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2248_ (.A1(_1400_),
    .A2(_1424_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2249_ (.A1(_1400_),
    .A2(_1424_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2250_ (.A1(_1398_),
    .A2(_1459_),
    .B(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2251_ (.A1(_1404_),
    .A2(_1422_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2252_ (.A1(_1402_),
    .A2(_1423_),
    .B(_1462_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2253_ (.A1(_1415_),
    .A2(_1416_),
    .B(_1419_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2254_ (.A1(_1405_),
    .A2(_1411_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2255_ (.A1(_1412_),
    .A2(_1421_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2256_ (.A1(_0780_),
    .A2(_1258_),
    .B1(_1336_),
    .B2(_1410_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2257_ (.A1(_0804_),
    .A2(_1103_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2258_ (.A1(_1408_),
    .A2(_0091_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2259_ (.A1(_1336_),
    .A2(_0092_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2260_ (.A1(_0090_),
    .A2(_0093_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2261_ (.A1(_0796_),
    .A2(_1406_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2262_ (.A1(_1407_),
    .A2(_1409_),
    .B(_0095_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2263_ (.A1(_0819_),
    .A2(_1043_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2264_ (.A1(_0096_),
    .A2(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2265_ (.A1(_0831_),
    .A2(_0985_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2266_ (.A1(_0098_),
    .A2(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2267_ (.A1(_0094_),
    .A2(_0100_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2268_ (.A1(_0088_),
    .A2(_0089_),
    .B(_0101_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2269_ (.A1(_0088_),
    .A2(_0089_),
    .A3(_0101_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2270_ (.A1(_0102_),
    .A2(_0103_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2271_ (.A1(_0087_),
    .A2(_0104_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2272_ (.A1(_0086_),
    .A2(_0105_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2273_ (.A1(_0834_),
    .A2(_1427_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2274_ (.I(_1310_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2275_ (.I(_0108_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2276_ (.A1(_0824_),
    .A2(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2277_ (.A1(_0107_),
    .A2(_0110_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2278_ (.A1(_1461_),
    .A2(_0106_),
    .A3(_0111_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2279_ (.A1(_1456_),
    .A2(_1458_),
    .A3(_0112_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2280_ (.A1(_0776_),
    .A2(_1215_),
    .B1(_1306_),
    .B2(_1387_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2281_ (.I(_1312_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2282_ (.A1(_0811_),
    .A2(_0115_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2283_ (.A1(_1385_),
    .A2(_0116_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2284_ (.A1(_1306_),
    .A2(_0117_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2285_ (.A1(_0114_),
    .A2(_0118_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2286_ (.A1(_0113_),
    .A2(_0119_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2287_ (.A1(_1451_),
    .A2(_1453_),
    .A3(_0120_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2288_ (.A1(_1447_),
    .A2(_0121_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2289_ (.A1(_1442_),
    .A2(_0122_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2290_ (.A1(_0822_),
    .A2(_0123_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2291_ (.A1(net123),
    .A2(_0124_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2292_ (.I(_0125_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2293_ (.A1(_1442_),
    .A2(_0122_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2294_ (.A1(_1447_),
    .A2(_0121_),
    .B(_0126_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2295_ (.A1(_0833_),
    .A2(_0127_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2296_ (.A1(_1452_),
    .A2(_1443_),
    .A3(_0120_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2297_ (.A1(_1452_),
    .A2(_1443_),
    .B(_0120_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2298_ (.A1(_1451_),
    .A2(_0129_),
    .B(_0130_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2299_ (.A1(_0086_),
    .A2(_0105_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2300_ (.A1(_1461_),
    .A2(_0106_),
    .B(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2301_ (.A1(_0087_),
    .A2(_0104_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(_0102_),
    .A2(_0134_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2303_ (.A1(_0832_),
    .A2(_0109_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2304_ (.A1(_0135_),
    .A2(_0136_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2305_ (.A1(_1407_),
    .A2(_0091_),
    .B(_0095_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2306_ (.A1(_0821_),
    .A2(_0115_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2307_ (.A1(_0820_),
    .A2(_0108_),
    .A3(_0096_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2308_ (.A1(_0832_),
    .A2(_1427_),
    .A3(_0098_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2309_ (.A1(_0140_),
    .A2(_0141_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2310_ (.A1(_0139_),
    .A2(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2311_ (.A1(_0138_),
    .A2(_0143_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2312_ (.A1(_0094_),
    .A2(_0100_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2313_ (.A1(_0090_),
    .A2(_0093_),
    .B(_0145_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2314_ (.I0(_1270_),
    .I1(_1335_),
    .S(_0092_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2315_ (.A1(_0144_),
    .A2(_0146_),
    .A3(_0147_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2316_ (.A1(_0133_),
    .A2(_0137_),
    .A3(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2317_ (.A1(_1461_),
    .A2(_0106_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2318_ (.A1(_0107_),
    .A2(_0110_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2319_ (.A1(_0107_),
    .A2(_0110_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2320_ (.A1(_0150_),
    .A2(_0151_),
    .B(_0152_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2321_ (.A1(_0113_),
    .A2(_0119_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2322_ (.A1(_0114_),
    .A2(_0118_),
    .B(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2323_ (.A1(_0824_),
    .A2(_0115_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2324_ (.A1(_0834_),
    .A2(_0109_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2325_ (.A1(_1384_),
    .A2(_0116_),
    .B(_1457_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2326_ (.I(_0112_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2327_ (.A1(_1458_),
    .A2(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2328_ (.A1(_1458_),
    .A2(_0159_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2329_ (.A1(_1456_),
    .A2(_0160_),
    .B(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2330_ (.A1(_0157_),
    .A2(_0158_),
    .A3(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2331_ (.I0(_1220_),
    .I1(_1305_),
    .S(_0117_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2332_ (.A1(_0156_),
    .A2(_0163_),
    .A3(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2333_ (.A1(_0153_),
    .A2(_0155_),
    .A3(_0165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2334_ (.A1(_0131_),
    .A2(_0149_),
    .A3(_0166_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2335_ (.A1(_0822_),
    .A2(_0123_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2336_ (.A1(_1439_),
    .A2(_0124_),
    .B(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2337_ (.A1(_0128_),
    .A2(_0167_),
    .A3(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2338_ (.I(_0170_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2339_ (.A1(_0734_),
    .A2(_1058_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2340_ (.I(_0171_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2341_ (.A1(_0757_),
    .A2(\t_reg[0] ),
    .A3(_0729_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2342_ (.A1(\t_reg[1] ),
    .A2(_0727_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2343_ (.A1(_0769_),
    .A2(_0173_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2344_ (.A1(_0172_),
    .A2(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2345_ (.I(_0175_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2346_ (.A1(_0769_),
    .A2(\t_reg[1] ),
    .A3(_0728_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2347_ (.A1(\delta_t[0] ),
    .A2(\t_reg[0] ),
    .A3(_0728_),
    .A4(_0174_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2348_ (.A1(_0176_),
    .A2(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2349_ (.A1(_0777_),
    .A2(_0889_),
    .A3(_0178_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2350_ (.I(_0179_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2351_ (.A1(_0777_),
    .A2(_0889_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2352_ (.A1(_0176_),
    .A2(_0177_),
    .B(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2353_ (.A1(_0777_),
    .A2(_0889_),
    .B(_0181_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2354_ (.A1(_0788_),
    .A2(_0891_),
    .A3(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2355_ (.I(_0183_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2356_ (.I(\delta_t[4] ),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2357_ (.A1(\delta_t[3] ),
    .A2(_0891_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2358_ (.A1(_0788_),
    .A2(_0891_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2359_ (.A1(_0182_),
    .A2(_0185_),
    .B(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2360_ (.A1(_0184_),
    .A2(_0900_),
    .A3(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2361_ (.I(_0188_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2362_ (.A1(\t_reg[5] ),
    .A2(_0728_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2363_ (.A1(_0184_),
    .A2(_0900_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2364_ (.A1(_0184_),
    .A2(_0900_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2365_ (.A1(_0187_),
    .A2(_0190_),
    .B(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2366_ (.A1(\delta_t[5] ),
    .A2(_0189_),
    .A3(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2367_ (.I(_0193_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2368_ (.A1(_0899_),
    .A2(_0189_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2369_ (.A1(_0899_),
    .A2(_0189_),
    .B(_0192_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2370_ (.A1(_0194_),
    .A2(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2371_ (.A1(_0827_),
    .A2(_0922_),
    .A3(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2372_ (.I(_0197_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2373_ (.I(_0921_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2374_ (.A1(_0876_),
    .A2(_0922_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2375_ (.A1(_0827_),
    .A2(\t_reg[6] ),
    .A3(_0729_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2376_ (.A1(_0196_),
    .A2(_0199_),
    .B(_0200_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2377_ (.A1(_0198_),
    .A2(_1015_),
    .A3(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2378_ (.I(_0202_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2379_ (.A1(\delta_t[8] ),
    .A2(_1020_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2380_ (.A1(_0198_),
    .A2(_1015_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2381_ (.A1(_0201_),
    .A2(_0204_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2382_ (.A1(_0198_),
    .A2(_1015_),
    .B(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2383_ (.A1(_0203_),
    .A2(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2384_ (.I(_0207_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2385_ (.A1(\delta_t[8] ),
    .A2(_1020_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2386_ (.A1(_0203_),
    .A2(_0206_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2387_ (.A1(_0208_),
    .A2(_0209_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2388_ (.A1(_0839_),
    .A2(_1082_),
    .A3(_0210_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2389_ (.I(_0211_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2390_ (.A1(\t_reg[0] ),
    .A2(_0729_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2391_ (.A1(_0757_),
    .A2(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2392_ (.I(_0213_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2393_ (.A1(_0749_),
    .A2(_1223_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2394_ (.A1(_0766_),
    .A2(_0937_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2395_ (.A1(_0772_),
    .A2(_0935_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2396_ (.A1(_0215_),
    .A2(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2397_ (.A1(_0214_),
    .A2(_0217_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2398_ (.A1(_0768_),
    .A2(_0946_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2399_ (.A1(_0750_),
    .A2(_0952_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2400_ (.A1(_0219_),
    .A2(_0220_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2401_ (.A1(_0218_),
    .A2(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2402_ (.A1(_0218_),
    .A2(_0221_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2403_ (.A1(_0933_),
    .A2(_0222_),
    .B(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2404_ (.A1(_0214_),
    .A2(_0217_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2405_ (.A1(_0749_),
    .A2(_1307_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2406_ (.A1(_0215_),
    .A2(_0216_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2407_ (.A1(_0766_),
    .A2(_1110_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2408_ (.A1(_0771_),
    .A2(_0980_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2409_ (.A1(_0784_),
    .A2(_0934_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2410_ (.A1(_0228_),
    .A2(_0229_),
    .A3(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2411_ (.A1(_0227_),
    .A2(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2412_ (.A1(_0226_),
    .A2(_0232_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2413_ (.A1(_0225_),
    .A2(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2414_ (.A1(_0974_),
    .A2(_0234_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2415_ (.A1(_0932_),
    .A2(_0222_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2416_ (.A1(_0219_),
    .A2(_0220_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2417_ (.A1(_0751_),
    .A2(_0993_),
    .A3(_0215_),
    .A4(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2418_ (.A1(_0750_),
    .A2(_0997_),
    .B(_0946_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2419_ (.A1(_0996_),
    .A2(_0239_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2420_ (.A1(_0751_),
    .A2(_0993_),
    .B1(_0996_),
    .B2(_0239_),
    .C(_0237_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2421_ (.A1(_0238_),
    .A2(_0240_),
    .B(_0241_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2422_ (.A1(_0236_),
    .A2(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2423_ (.A1(_0224_),
    .A2(_0235_),
    .B(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2424_ (.A1(_0224_),
    .A2(_0235_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2425_ (.I(_0974_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2426_ (.A1(_0225_),
    .A2(_0233_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2427_ (.A1(_0246_),
    .A2(_0234_),
    .B(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2428_ (.A1(_0227_),
    .A2(_0231_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2429_ (.A1(_0226_),
    .A2(_0232_),
    .B(_0249_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2430_ (.I(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2431_ (.A1(_0749_),
    .A2(_1309_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2432_ (.A1(_0801_),
    .A2(_1278_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2433_ (.A1(_0252_),
    .A2(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2434_ (.A1(_0229_),
    .A2(_0230_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2435_ (.A1(_0229_),
    .A2(_0230_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2436_ (.A1(_0228_),
    .A2(_0255_),
    .B(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2437_ (.A1(_0767_),
    .A2(_1176_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2438_ (.A1(\c[0][3] ),
    .A2(_0906_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2439_ (.A1(_0772_),
    .A2(_1110_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2440_ (.A1(_0259_),
    .A2(_0260_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2441_ (.A1(_0258_),
    .A2(_0261_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2442_ (.A1(_0257_),
    .A2(_0262_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2443_ (.A1(_0254_),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2444_ (.A1(_1030_),
    .A2(_0251_),
    .A3(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2445_ (.A1(_0248_),
    .A2(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2446_ (.A1(_0244_),
    .A2(_0245_),
    .B(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2447_ (.A1(_0244_),
    .A2(_0245_),
    .A3(_0266_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2448_ (.A1(_0267_),
    .A2(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2449_ (.A1(_0997_),
    .A2(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2450_ (.A1(_0248_),
    .A2(_0265_),
    .B(_0267_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2451_ (.A1(_0250_),
    .A2(_0264_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2452_ (.A1(_1030_),
    .A2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2453_ (.A1(_0251_),
    .A2(_0264_),
    .B(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2454_ (.A1(_0252_),
    .A2(_0253_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2455_ (.A1(_0257_),
    .A2(_0262_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2456_ (.A1(_0254_),
    .A2(_0263_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2457_ (.A1(_0276_),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2458_ (.A1(_0259_),
    .A2(_0260_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2459_ (.A1(_0767_),
    .A2(_1177_),
    .A3(_0261_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2460_ (.A1(_0279_),
    .A2(_0280_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2461_ (.A1(\c[0][3] ),
    .A2(_0940_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2462_ (.A1(_0771_),
    .A2(_0986_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2463_ (.A1(_0282_),
    .A2(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2464_ (.A1(_0766_),
    .A2(_1309_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2465_ (.A1(_0284_),
    .A2(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2466_ (.A1(_0281_),
    .A2(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2467_ (.A1(\c[0][0] ),
    .A2(_1217_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2468_ (.A1(\c[0][4] ),
    .A2(_0937_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2469_ (.A1(_0288_),
    .A2(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2470_ (.A1(_0812_),
    .A2(_0944_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2471_ (.A1(_0290_),
    .A2(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2472_ (.A1(_0287_),
    .A2(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2473_ (.A1(_0278_),
    .A2(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2474_ (.A1(_1130_),
    .A2(_0275_),
    .A3(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2475_ (.A1(_0274_),
    .A2(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2476_ (.A1(_0761_),
    .A2(_0271_),
    .A3(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2477_ (.A1(_0270_),
    .A2(_0297_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2478_ (.I(_0298_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2479_ (.A1(_0271_),
    .A2(_0296_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2480_ (.A1(_0270_),
    .A2(_0297_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2481_ (.A1(_0910_),
    .A2(_0299_),
    .B(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2482_ (.A1(_1130_),
    .A2(_0252_),
    .A3(_0253_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2483_ (.A1(_1130_),
    .A2(_0275_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2484_ (.A1(_0278_),
    .A2(_0293_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2485_ (.A1(_0303_),
    .A2(_0294_),
    .B(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(\c[0][0] ),
    .A2(_1180_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2487_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2488_ (.A1(_0307_),
    .A2(_0289_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2489_ (.A1(_0290_),
    .A2(_0291_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2490_ (.A1(_0308_),
    .A2(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2491_ (.A1(_0825_),
    .A2(_1278_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2492_ (.I(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2493_ (.A1(_1141_),
    .A2(_1169_),
    .A3(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(_0287_),
    .A2(_0292_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2495_ (.A1(_0281_),
    .A2(_0286_),
    .B(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2496_ (.A1(_0767_),
    .A2(_1309_),
    .A3(_0284_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2497_ (.A1(_0282_),
    .A2(_0283_),
    .B(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2498_ (.A1(\c[0][1] ),
    .A2(_1103_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2499_ (.A1(\c[0][3] ),
    .A2(_0985_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(\c[0][2] ),
    .A2(_1044_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2501_ (.A1(_0319_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2502_ (.A1(_0318_),
    .A2(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2503_ (.A1(_0317_),
    .A2(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2504_ (.A1(\c[0][4] ),
    .A2(_1222_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2505_ (.A1(_0306_),
    .A2(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2506_ (.A1(_0801_),
    .A2(_1222_),
    .A3(_0288_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_0325_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2508_ (.A1(_0812_),
    .A2(_0947_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2509_ (.A1(_0327_),
    .A2(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2510_ (.A1(_0323_),
    .A2(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2511_ (.A1(_0315_),
    .A2(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2512_ (.A1(_0310_),
    .A2(_0313_),
    .A3(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2513_ (.A1(_0302_),
    .A2(_0305_),
    .A3(net117),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2514_ (.A1(_0274_),
    .A2(_0295_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2515_ (.A1(_0271_),
    .A2(_0296_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2516_ (.A1(_0781_),
    .A2(_0333_),
    .A3(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2517_ (.A1(_0301_),
    .A2(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2518_ (.I(_0337_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2519_ (.A1(_0333_),
    .A2(_0335_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2520_ (.A1(_0301_),
    .A2(_0336_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2521_ (.A1(_0782_),
    .A2(_0338_),
    .B(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2522_ (.A1(_0333_),
    .A2(_0335_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2523_ (.A1(_0310_),
    .A2(_0313_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2524_ (.A1(_0305_),
    .A2(_0332_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2525_ (.A1(_0305_),
    .A2(_0332_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2526_ (.A1(_0302_),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2527_ (.A1(_0313_),
    .A2(_0310_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2528_ (.A1(_0315_),
    .A2(_0330_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2529_ (.A1(_0346_),
    .A2(_0331_),
    .B(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2530_ (.A1(_0317_),
    .A2(_0322_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2531_ (.A1(_0323_),
    .A2(_0329_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2532_ (.A1(_0349_),
    .A2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2533_ (.A1(_0319_),
    .A2(_0320_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2534_ (.A1(_0318_),
    .A2(_0321_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2535_ (.A1(_0352_),
    .A2(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2536_ (.A1(_0784_),
    .A2(_1184_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2537_ (.I(_0771_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2538_ (.A1(_0356_),
    .A2(_1254_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2539_ (.A1(_0355_),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2540_ (.A1(_0318_),
    .A2(_0354_),
    .A3(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(\c[0][5] ),
    .A2(_0941_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2542_ (.A1(\c[0][4] ),
    .A2(_0986_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2543_ (.A1(_0306_),
    .A2(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2544_ (.A1(_0360_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2545_ (.A1(_0359_),
    .A2(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2546_ (.I(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2547_ (.A1(_0351_),
    .A2(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2548_ (.I(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2549_ (.A1(_1233_),
    .A2(_0312_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2550_ (.A1(_0327_),
    .A2(_0328_),
    .B(_0326_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2551_ (.A1(\c[0][6] ),
    .A2(_0948_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2552_ (.A1(\c[0][7] ),
    .A2(_1278_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2553_ (.A1(_0370_),
    .A2(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2554_ (.A1(_1243_),
    .A2(_1276_),
    .A3(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2555_ (.A1(_0368_),
    .A2(_0369_),
    .A3(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2556_ (.A1(_0348_),
    .A2(_0367_),
    .A3(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2557_ (.A1(_0342_),
    .A2(_0345_),
    .A3(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2558_ (.A1(_0791_),
    .A2(_0341_),
    .A3(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2559_ (.A1(_0340_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2560_ (.I(_0378_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2561_ (.A1(_0341_),
    .A2(net116),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2562_ (.A1(_0792_),
    .A2(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2563_ (.A1(_0340_),
    .A2(_0377_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2564_ (.A1(_0342_),
    .A2(_0375_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2565_ (.A1(_0333_),
    .A2(_0335_),
    .A3(_0376_),
    .B1(_0382_),
    .B2(net114),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2566_ (.A1(_0366_),
    .A2(_0374_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2567_ (.A1(_0310_),
    .A2(net135),
    .A3(_0375_),
    .B1(_0384_),
    .B2(net113),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2568_ (.A1(_0369_),
    .A2(_0373_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2569_ (.A1(_0369_),
    .A2(_0373_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2570_ (.A1(_0368_),
    .A2(_0386_),
    .B(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2571_ (.A1(_0351_),
    .A2(_0365_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2572_ (.A1(_0367_),
    .A2(_0374_),
    .B(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2573_ (.I(_0318_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2574_ (.A1(_0391_),
    .A2(_0358_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2575_ (.A1(_0391_),
    .A2(_0358_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2576_ (.A1(_0354_),
    .A2(_0392_),
    .A3(_0393_),
    .B1(_0359_),
    .B2(_0363_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2577_ (.A1(_0356_),
    .A2(_1254_),
    .A3(_0355_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2578_ (.A1(_0784_),
    .A2(_0772_),
    .B(_1217_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2579_ (.A1(_0785_),
    .A2(_0357_),
    .B(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2580_ (.A1(_0391_),
    .A2(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2581_ (.A1(_0785_),
    .A2(_0768_),
    .A3(_0357_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2582_ (.A1(_0395_),
    .A2(_0392_),
    .A3(_0398_),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2583_ (.A1(\c[0][5] ),
    .A2(_1177_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2584_ (.A1(_0801_),
    .A2(_1310_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2585_ (.A1(_0307_),
    .A2(_0401_),
    .A3(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2586_ (.I(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2587_ (.A1(_0400_),
    .A2(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2588_ (.A1(_0394_),
    .A2(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2589_ (.I(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2590_ (.A1(_1243_),
    .A2(_1276_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2591_ (.A1(_0370_),
    .A2(_0371_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2592_ (.A1(_0370_),
    .A2(_0371_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2593_ (.A1(_0408_),
    .A2(_0409_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2594_ (.A1(_0288_),
    .A2(_0361_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2595_ (.A1(_0360_),
    .A2(_0362_),
    .B(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2596_ (.A1(\c[0][7] ),
    .A2(_0952_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2597_ (.A1(_0825_),
    .A2(_1355_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2598_ (.A1(_0414_),
    .A2(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2599_ (.A1(_1325_),
    .A2(_1353_),
    .A3(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2600_ (.A1(_0411_),
    .A2(_0413_),
    .A3(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2601_ (.A1(_0390_),
    .A2(_0407_),
    .A3(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2602_ (.A1(_0385_),
    .A2(_0388_),
    .A3(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2603_ (.A1(_0796_),
    .A2(_0383_),
    .A3(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2604_ (.A1(_0380_),
    .A2(_0381_),
    .B(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2605_ (.A1(_0380_),
    .A2(_0381_),
    .A3(_0421_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2606_ (.A1(_0422_),
    .A2(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2607_ (.I(_0424_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2608_ (.A1(_0420_),
    .A2(_0383_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2609_ (.A1(_0383_),
    .A2(_0420_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2610_ (.A1(_0797_),
    .A2(_0425_),
    .A3(_0426_),
    .B(_0422_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2611_ (.I(_0805_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2612_ (.A1(_0388_),
    .A2(_0419_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2613_ (.A1(net115),
    .A2(_0429_),
    .B(_0425_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2614_ (.A1(_0407_),
    .A2(_0418_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2615_ (.A1(_0390_),
    .A2(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2616_ (.A1(_0388_),
    .A2(_0419_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2617_ (.A1(_0432_),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2618_ (.A1(_0413_),
    .A2(_0417_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2619_ (.A1(_0413_),
    .A2(_0417_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2620_ (.A1(_0411_),
    .A2(_0435_),
    .B(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(_0394_),
    .A2(_0405_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2622_ (.A1(_0407_),
    .A2(_0418_),
    .B(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2623_ (.I(_0399_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2624_ (.A1(_0400_),
    .A2(_0404_),
    .B(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2625_ (.A1(_0391_),
    .A2(_0396_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2626_ (.A1(_0440_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2627_ (.A1(_0812_),
    .A2(_0108_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2628_ (.A1(_0802_),
    .A2(_0288_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2629_ (.A1(_0802_),
    .A2(_0750_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2630_ (.A1(_1312_),
    .A2(_0445_),
    .A3(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2631_ (.A1(_0444_),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2632_ (.A1(_0443_),
    .A2(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2633_ (.A1(_0441_),
    .A2(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2634_ (.A1(_1325_),
    .A2(_1353_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2635_ (.A1(_0414_),
    .A2(_0415_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2636_ (.A1(_0451_),
    .A2(_0416_),
    .B(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2637_ (.A1(_0307_),
    .A2(_0402_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2638_ (.A1(_0307_),
    .A2(_0402_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2639_ (.A1(_0401_),
    .A2(_0454_),
    .B(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2640_ (.A1(\c[0][7] ),
    .A2(_1355_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2641_ (.A1(_0825_),
    .A2(_1307_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2642_ (.A1(_0457_),
    .A2(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2643_ (.A1(_1398_),
    .A2(_1425_),
    .A3(_0459_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2644_ (.A1(_0453_),
    .A2(_0456_),
    .A3(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2645_ (.A1(_0450_),
    .A2(_0461_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2646_ (.A1(_0437_),
    .A2(_0439_),
    .A3(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2647_ (.A1(_0434_),
    .A2(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2648_ (.A1(_0428_),
    .A2(_0430_),
    .A3(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2649_ (.A1(_0427_),
    .A2(_0465_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2650_ (.I(_0466_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2651_ (.A1(_0430_),
    .A2(_0464_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2652_ (.A1(_0427_),
    .A2(_0465_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2653_ (.A1(_0428_),
    .A2(_0467_),
    .B(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2654_ (.A1(_0434_),
    .A2(_0463_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2655_ (.A1(_0434_),
    .A2(_0463_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2656_ (.A1(_0430_),
    .A2(_0470_),
    .B(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2657_ (.A1(_0439_),
    .A2(_0462_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2658_ (.A1(_0439_),
    .A2(_0462_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2659_ (.A1(_0437_),
    .A2(_0473_),
    .B(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2660_ (.A1(_1454_),
    .A2(_0459_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2661_ (.A1(_0456_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2662_ (.A1(_0456_),
    .A2(_0460_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2663_ (.A1(_0453_),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2664_ (.A1(_0477_),
    .A2(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2665_ (.A1(_0441_),
    .A2(_0449_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2666_ (.A1(_0450_),
    .A2(_0461_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2667_ (.A1(_0481_),
    .A2(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2668_ (.A1(_0457_),
    .A2(_0458_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2669_ (.A1(_1454_),
    .A2(_0459_),
    .B(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2670_ (.I(_0447_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2671_ (.A1(_0444_),
    .A2(_0486_),
    .B(_0445_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2672_ (.A1(_0835_),
    .A2(_1427_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(_0826_),
    .A2(_0108_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2674_ (.A1(_0488_),
    .A2(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2675_ (.A1(_1461_),
    .A2(_0106_),
    .A3(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2676_ (.A1(_0485_),
    .A2(_0487_),
    .A3(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2677_ (.A1(_0443_),
    .A2(_0448_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2678_ (.A1(_0440_),
    .A2(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2679_ (.A1(_0813_),
    .A2(_1254_),
    .B(_0486_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2680_ (.A1(_0814_),
    .A2(_0486_),
    .B(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2681_ (.A1(_0443_),
    .A2(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2682_ (.I(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2683_ (.A1(_0494_),
    .A2(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2684_ (.A1(_0492_),
    .A2(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2685_ (.A1(_0480_),
    .A2(_0483_),
    .A3(_0500_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2686_ (.A1(_0475_),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2687_ (.A1(_0472_),
    .A2(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2688_ (.A1(_0821_),
    .A2(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2689_ (.A1(_0469_),
    .A2(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2690_ (.I(_0505_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2691_ (.A1(_0821_),
    .A2(_0503_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2692_ (.A1(_0469_),
    .A2(_0504_),
    .B(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2693_ (.I(_0501_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2694_ (.A1(_0475_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2695_ (.A1(_0472_),
    .A2(_0502_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2696_ (.A1(_0509_),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2697_ (.A1(_0483_),
    .A2(_0500_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2698_ (.A1(_0483_),
    .A2(_0500_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2699_ (.A1(_0480_),
    .A2(_0512_),
    .B(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2700_ (.A1(_0835_),
    .A2(_0109_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2701_ (.A1(_0488_),
    .A2(_0489_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2702_ (.A1(_0488_),
    .A2(_0489_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2703_ (.A1(_0150_),
    .A2(_0516_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2704_ (.A1(_0515_),
    .A2(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2705_ (.A1(_0826_),
    .A2(_0115_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2706_ (.A1(_0492_),
    .A2(_0499_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2707_ (.A1(_0494_),
    .A2(_0498_),
    .B(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2708_ (.I(_0491_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2709_ (.A1(_0487_),
    .A2(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2710_ (.A1(_0487_),
    .A2(_0523_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2711_ (.A1(_0485_),
    .A2(_0524_),
    .B(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2712_ (.A1(_0814_),
    .A2(_0486_),
    .B(_0445_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2713_ (.I0(_0440_),
    .I1(_0442_),
    .S(_0496_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2714_ (.A1(_0527_),
    .A2(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2715_ (.A1(_0149_),
    .A2(_0526_),
    .A3(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2716_ (.A1(_0520_),
    .A2(_0522_),
    .A3(_0530_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2717_ (.A1(_0514_),
    .A2(_0519_),
    .A3(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2718_ (.A1(_0511_),
    .A2(_0532_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2719_ (.A1(_0833_),
    .A2(_0507_),
    .A3(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2720_ (.I(_0534_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2721_ (.A1(_0997_),
    .A2(_0269_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2722_ (.I(_0535_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2723_ (.A1(net28),
    .A2(net38),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2724_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2725_ (.A1(net25),
    .A2(_0754_),
    .A3(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2726_ (.A1(net22),
    .A2(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2727_ (.I(net2),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2728_ (.I(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2729_ (.A1(_0837_),
    .A2(_0538_),
    .B(_0539_),
    .C(_0541_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2730_ (.A1(net23),
    .A2(_0538_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2731_ (.A1(_0839_),
    .A2(_0538_),
    .B(_0542_),
    .C(_0541_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2732_ (.A1(net24),
    .A2(_0536_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2733_ (.A1(_0754_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2734_ (.I(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2735_ (.A1(_0757_),
    .A2(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2736_ (.A1(net24),
    .A2(_0537_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2737_ (.A1(_0838_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2738_ (.A1(net6),
    .A2(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2739_ (.I(_0540_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2740_ (.I(_0550_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2741_ (.A1(_0546_),
    .A2(_0549_),
    .B(_0551_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2742_ (.A1(_0769_),
    .A2(_0545_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2743_ (.A1(net11),
    .A2(_0548_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2744_ (.A1(_0552_),
    .A2(_0553_),
    .B(_0551_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2745_ (.I(_0544_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2746_ (.I(_0544_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2747_ (.A1(net16),
    .A2(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2748_ (.A1(_0879_),
    .A2(_0554_),
    .B(_0556_),
    .C(_0541_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2749_ (.A1(_0788_),
    .A2(_0545_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2750_ (.A1(net17),
    .A2(_0548_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2751_ (.A1(_0557_),
    .A2(_0558_),
    .B(_0551_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2752_ (.A1(net18),
    .A2(_0555_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2753_ (.I(net2),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2754_ (.I(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2755_ (.A1(_0184_),
    .A2(_0554_),
    .B(_0559_),
    .C(_0561_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2756_ (.A1(net19),
    .A2(_0555_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2757_ (.A1(_0899_),
    .A2(_0554_),
    .B(_0562_),
    .C(_0561_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2758_ (.A1(net20),
    .A2(_0555_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2759_ (.A1(_0876_),
    .A2(_0554_),
    .B(_0563_),
    .C(_0561_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2760_ (.A1(net21),
    .A2(_0544_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2761_ (.A1(_0198_),
    .A2(_0545_),
    .B(_0564_),
    .C(_0561_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2762_ (.A1(net26),
    .A2(_0537_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2763_ (.A1(_0755_),
    .A2(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2764_ (.A1(net7),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2765_ (.I(_0560_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2766_ (.A1(_0730_),
    .A2(_0566_),
    .B(_0567_),
    .C(_0568_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2767_ (.A1(_0806_),
    .A2(_0547_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2768_ (.I(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2769_ (.I(_0569_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2770_ (.A1(net6),
    .A2(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2771_ (.A1(_0734_),
    .A2(_0570_),
    .B(_0572_),
    .C(_0568_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(net11),
    .A2(_0571_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2773_ (.A1(_0761_),
    .A2(_0570_),
    .B(_0573_),
    .C(_0568_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2774_ (.I(_0569_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2775_ (.A1(_0782_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2776_ (.A1(_0807_),
    .A2(_0547_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2777_ (.A1(net16),
    .A2(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2778_ (.A1(_0575_),
    .A2(_0577_),
    .B(_0551_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2779_ (.A1(_0792_),
    .A2(_0574_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(net17),
    .A2(_0576_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2781_ (.I(_0540_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2782_ (.I(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2783_ (.A1(_0578_),
    .A2(_0579_),
    .B(_0581_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2784_ (.A1(net18),
    .A2(_0571_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2785_ (.A1(_0797_),
    .A2(_0570_),
    .B(_0582_),
    .C(_0568_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2786_ (.A1(net19),
    .A2(_0571_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2787_ (.I(_0560_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2788_ (.A1(_0428_),
    .A2(_0570_),
    .B(_0583_),
    .C(_0584_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2789_ (.A1(_0822_),
    .A2(_0574_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2790_ (.A1(net20),
    .A2(_0576_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2791_ (.A1(_0585_),
    .A2(_0586_),
    .B(_0581_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2792_ (.A1(_0833_),
    .A2(_0574_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2793_ (.A1(net21),
    .A2(_0576_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2794_ (.A1(_0587_),
    .A2(_0588_),
    .B(_0581_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2795_ (.A1(net26),
    .A2(_0537_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2796_ (.A1(_0806_),
    .A2(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2797_ (.I(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2798_ (.A1(\a[1][0] ),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(_0807_),
    .A2(_0589_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2800_ (.I(_0593_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(net7),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2802_ (.A1(_0592_),
    .A2(_0595_),
    .B(_0581_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2803_ (.A1(\a[1][1] ),
    .A2(_0591_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2804_ (.A1(net8),
    .A2(_0594_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2805_ (.I(_0580_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2806_ (.A1(_0596_),
    .A2(_0597_),
    .B(_0598_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2807_ (.A1(\a[1][2] ),
    .A2(_0591_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2808_ (.A1(net9),
    .A2(_0594_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2809_ (.A1(_0599_),
    .A2(_0600_),
    .B(_0598_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2810_ (.A1(\a[1][3] ),
    .A2(_0591_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2811_ (.A1(net10),
    .A2(_0594_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2812_ (.A1(_0601_),
    .A2(_0602_),
    .B(_0598_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2813_ (.I(_0590_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2814_ (.A1(\a[1][4] ),
    .A2(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2815_ (.I(_0593_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2816_ (.A1(net12),
    .A2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2817_ (.A1(_0604_),
    .A2(_0606_),
    .B(_0598_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2818_ (.A1(\a[1][5] ),
    .A2(_0603_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2819_ (.A1(net13),
    .A2(_0605_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2820_ (.I(_0580_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2821_ (.A1(_0607_),
    .A2(_0608_),
    .B(_0609_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(\a[1][6] ),
    .A2(_0603_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2823_ (.A1(net14),
    .A2(_0605_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2824_ (.A1(_0610_),
    .A2(_0611_),
    .B(_0609_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2825_ (.A1(\a[1][7] ),
    .A2(_0603_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2826_ (.A1(net15),
    .A2(_0605_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2827_ (.A1(_0612_),
    .A2(_0613_),
    .B(_0609_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2828_ (.A1(_0746_),
    .A2(_0543_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2829_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2830_ (.A1(_0743_),
    .A2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2831_ (.A1(_0745_),
    .A2(_0543_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2832_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2833_ (.A1(net6),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2834_ (.A1(_0616_),
    .A2(_0619_),
    .B(_0609_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2835_ (.A1(_0764_),
    .A2(_0615_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2836_ (.A1(net11),
    .A2(_0618_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2837_ (.I(_0580_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2838_ (.A1(_0620_),
    .A2(_0621_),
    .B(_0622_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2839_ (.A1(_0776_),
    .A2(_0615_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2840_ (.A1(net16),
    .A2(_0618_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2841_ (.A1(_0623_),
    .A2(_0624_),
    .B(_0622_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2842_ (.A1(_0787_),
    .A2(_0615_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2843_ (.A1(net17),
    .A2(_0618_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2844_ (.A1(_0625_),
    .A2(_0626_),
    .B(_0622_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2845_ (.I(_0614_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2846_ (.A1(_0799_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2847_ (.I(_0617_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2848_ (.A1(net18),
    .A2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2849_ (.A1(_0628_),
    .A2(_0630_),
    .B(_0622_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2850_ (.A1(_0811_),
    .A2(_0627_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2851_ (.A1(net19),
    .A2(_0629_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2852_ (.I(_0540_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2853_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2854_ (.A1(_0631_),
    .A2(_0632_),
    .B(_0634_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2855_ (.A1(_0824_),
    .A2(_0627_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2856_ (.A1(net20),
    .A2(_0629_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2857_ (.A1(_0635_),
    .A2(_0636_),
    .B(_0634_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2858_ (.A1(_0834_),
    .A2(_0627_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2859_ (.A1(net21),
    .A2(_0629_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2860_ (.A1(_0637_),
    .A2(_0638_),
    .B(_0634_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2861_ (.I(\b[1][0] ),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2862_ (.A1(_0745_),
    .A2(_0565_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2863_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2864_ (.I(_0640_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2865_ (.A1(net7),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2866_ (.A1(_0639_),
    .A2(_0641_),
    .B(_0643_),
    .C(_0584_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2867_ (.A1(net8),
    .A2(_0642_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2868_ (.A1(_0841_),
    .A2(_0641_),
    .B(_0644_),
    .C(_0584_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2869_ (.A1(net9),
    .A2(_0642_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2870_ (.A1(_0847_),
    .A2(_0641_),
    .B(_0645_),
    .C(_0584_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2871_ (.A1(net10),
    .A2(_0642_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2872_ (.I(_0560_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2873_ (.A1(_0851_),
    .A2(_0641_),
    .B(_0646_),
    .C(_0647_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2874_ (.I(_0640_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2875_ (.I(_0640_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2876_ (.A1(net12),
    .A2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2877_ (.A1(_0854_),
    .A2(_0648_),
    .B(_0650_),
    .C(_0647_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2878_ (.A1(net13),
    .A2(_0649_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2879_ (.A1(_0858_),
    .A2(_0648_),
    .B(_0651_),
    .C(_0647_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2880_ (.A1(net14),
    .A2(_0649_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2881_ (.A1(_0861_),
    .A2(_0648_),
    .B(_0652_),
    .C(_0647_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2882_ (.A1(net15),
    .A2(_0649_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2883_ (.A1(_0864_),
    .A2(_0648_),
    .B(_0653_),
    .C(_0550_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2884_ (.A1(_0828_),
    .A2(_0744_),
    .A3(_0543_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2885_ (.I(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2886_ (.A1(_0751_),
    .A2(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2887_ (.A1(_0735_),
    .A2(_0744_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2888_ (.A1(_0547_),
    .A2(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2889_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2890_ (.A1(net6),
    .A2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2891_ (.A1(_0656_),
    .A2(_0660_),
    .B(_0634_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2892_ (.A1(_0768_),
    .A2(_0655_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2893_ (.A1(net11),
    .A2(_0659_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2894_ (.I(_0633_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2895_ (.A1(_0661_),
    .A2(_0662_),
    .B(_0663_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2896_ (.A1(net16),
    .A2(_0654_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2897_ (.A1(_0356_),
    .A2(_0655_),
    .B(_0664_),
    .C(_0550_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2898_ (.I(_0654_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2899_ (.A1(_0785_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2900_ (.A1(net17),
    .A2(_0659_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2901_ (.A1(_0666_),
    .A2(_0667_),
    .B(_0663_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2902_ (.A1(_0802_),
    .A2(_0665_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2903_ (.A1(net18),
    .A2(_0659_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2904_ (.A1(_0668_),
    .A2(_0669_),
    .B(_0663_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2905_ (.A1(net19),
    .A2(_0654_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2906_ (.A1(_0814_),
    .A2(_0655_),
    .B(_0670_),
    .C(_0550_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(_0826_),
    .A2(_0665_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2908_ (.A1(net20),
    .A2(_0658_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2909_ (.A1(_0671_),
    .A2(_0672_),
    .B(_0663_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2910_ (.A1(_0835_),
    .A2(_0665_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2911_ (.A1(net21),
    .A2(_0658_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2912_ (.I(_0633_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2913_ (.A1(_0673_),
    .A2(_0674_),
    .B(_0675_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2914_ (.A1(_0828_),
    .A2(_0752_),
    .A3(_0565_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2915_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2916_ (.A1(\c[1][0] ),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2917_ (.A1(_0589_),
    .A2(_0657_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2918_ (.I(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2919_ (.A1(net7),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2920_ (.A1(_0678_),
    .A2(_0681_),
    .B(_0675_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2921_ (.A1(\c[1][1] ),
    .A2(_0677_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2922_ (.A1(net8),
    .A2(_0680_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2923_ (.A1(_0682_),
    .A2(_0683_),
    .B(_0675_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2924_ (.A1(\c[1][2] ),
    .A2(_0677_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2925_ (.A1(net9),
    .A2(_0680_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2926_ (.A1(_0684_),
    .A2(_0685_),
    .B(_0675_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2927_ (.A1(\c[1][3] ),
    .A2(_0677_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2928_ (.A1(net10),
    .A2(_0680_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2929_ (.I(_0633_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2930_ (.A1(_0686_),
    .A2(_0687_),
    .B(_0688_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2931_ (.I(_0676_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2932_ (.A1(\c[1][4] ),
    .A2(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2933_ (.I(_0679_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2934_ (.A1(net12),
    .A2(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2935_ (.A1(_0690_),
    .A2(_0692_),
    .B(_0688_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2936_ (.A1(\c[1][5] ),
    .A2(_0689_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2937_ (.A1(net13),
    .A2(_0691_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2938_ (.A1(_0693_),
    .A2(_0694_),
    .B(_0688_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(\c[1][6] ),
    .A2(_0689_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2940_ (.A1(net14),
    .A2(_0691_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2941_ (.A1(_0695_),
    .A2(_0696_),
    .B(_0688_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2942_ (.A1(\c[1][7] ),
    .A2(_0689_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2943_ (.A1(net15),
    .A2(_0691_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2944_ (.A1(_0697_),
    .A2(_0698_),
    .B(_0541_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2945_ (.D(_0027_),
    .CLK(net73),
    .Q(\delta_t[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2946_ (.D(_0028_),
    .CLK(net73),
    .Q(\delta_t[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2947_ (.D(_0001_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2948_ (.D(_0002_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2949_ (.D(_0003_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2950_ (.D(_0004_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2951_ (.D(_0005_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2952_ (.D(_0006_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2953_ (.D(_0007_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2954_ (.D(_0008_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2955_ (.D(_0009_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2956_ (.D(_0010_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2957_ (.D(_0011_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2958_ (.D(_0012_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2959_ (.D(_0013_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2960_ (.D(_0014_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2961_ (.D(_0015_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2962_ (.D(_0016_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2963_ (.D(_0000_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2964_ (.D(_0017_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2965_ (.D(_0018_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2966_ (.D(_0019_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2967_ (.D(_0020_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2968_ (.D(_0021_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2969_ (.D(_0022_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2970_ (.D(_0023_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2971_ (.D(_0024_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2972_ (.D(_0025_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2973_ (.D(_0026_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\t_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2974_ (.D(_0029_),
    .CLK(net90),
    .Q(\delta_t[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2975_ (.D(_0030_),
    .CLK(net90),
    .Q(\delta_t[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2976_ (.D(_0031_),
    .CLK(net82),
    .Q(\delta_t[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2977_ (.D(_0032_),
    .CLK(net82),
    .Q(\delta_t[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2978_ (.D(_0033_),
    .CLK(net83),
    .Q(\delta_t[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _2979_ (.D(_0034_),
    .CLK(net74),
    .Q(\delta_t[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2980_ (.D(_0035_),
    .CLK(net74),
    .Q(\delta_t[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2981_ (.D(_0036_),
    .CLK(net75),
    .Q(\delta_t[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2982_ (.D(_0037_),
    .CLK(net89),
    .Q(bflip));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2983_ (.D(_0038_),
    .CLK(net75),
    .Q(\a[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2984_ (.D(_0039_),
    .CLK(net74),
    .Q(\a[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2985_ (.D(_0040_),
    .CLK(net83),
    .Q(\a[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2986_ (.D(_0041_),
    .CLK(net74),
    .Q(\a[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2987_ (.D(_0042_),
    .CLK(net75),
    .Q(\a[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2988_ (.D(_0043_),
    .CLK(net78),
    .Q(\a[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2989_ (.D(_0044_),
    .CLK(net76),
    .Q(\a[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2990_ (.D(_0045_),
    .CLK(net76),
    .Q(\a[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2991_ (.D(_0046_),
    .CLK(net90),
    .Q(\a[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2992_ (.D(_0047_),
    .CLK(net87),
    .Q(\a[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2993_ (.D(_0048_),
    .CLK(net87),
    .Q(\a[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2994_ (.D(_0049_),
    .CLK(net88),
    .Q(\a[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2995_ (.D(_0050_),
    .CLK(net91),
    .Q(\a[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2996_ (.D(_0051_),
    .CLK(net91),
    .Q(\a[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2997_ (.D(_0052_),
    .CLK(net91),
    .Q(\a[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2998_ (.D(_0053_),
    .CLK(net91),
    .Q(\a[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2999_ (.D(_0054_),
    .CLK(net92),
    .Q(\b[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3000_ (.D(_0055_),
    .CLK(net85),
    .Q(\b[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3001_ (.D(_0056_),
    .CLK(net85),
    .Q(\b[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3002_ (.D(_0057_),
    .CLK(net85),
    .Q(\b[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3003_ (.D(_0058_),
    .CLK(net85),
    .Q(\b[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3004_ (.D(_0059_),
    .CLK(net84),
    .Q(\b[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3005_ (.D(_0060_),
    .CLK(net77),
    .Q(\b[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3006_ (.D(_0061_),
    .CLK(net73),
    .Q(\b[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3007_ (.D(_0062_),
    .CLK(net87),
    .Q(\b[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3008_ (.D(_0063_),
    .CLK(net87),
    .Q(\b[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3009_ (.D(_0064_),
    .CLK(net88),
    .Q(\b[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3010_ (.D(_0065_),
    .CLK(net88),
    .Q(\b[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3011_ (.D(_0066_),
    .CLK(net92),
    .Q(\b[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3012_ (.D(_0067_),
    .CLK(net92),
    .Q(\b[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3013_ (.D(_0068_),
    .CLK(net93),
    .Q(\b[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3014_ (.D(_0069_),
    .CLK(net93),
    .Q(\b[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3015_ (.D(_0070_),
    .CLK(net84),
    .Q(\c[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3016_ (.D(_0071_),
    .CLK(net84),
    .Q(\c[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3017_ (.D(_0072_),
    .CLK(net84),
    .Q(\c[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3018_ (.D(_0073_),
    .CLK(net76),
    .Q(\c[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3019_ (.D(_0074_),
    .CLK(net76),
    .Q(\c[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3020_ (.D(_0075_),
    .CLK(net77),
    .Q(\c[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3021_ (.D(_0076_),
    .CLK(net73),
    .Q(\c[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3022_ (.D(_0077_),
    .CLK(net79),
    .Q(\c[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3023_ (.D(_0078_),
    .CLK(net83),
    .Q(\c[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3024_ (.D(_0079_),
    .CLK(net80),
    .Q(\c[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3025_ (.D(_0080_),
    .CLK(net80),
    .Q(\c[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3026_ (.D(_0081_),
    .CLK(net80),
    .Q(\c[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3027_ (.D(_0082_),
    .CLK(net81),
    .Q(\c[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3028_ (.D(_0083_),
    .CLK(net81),
    .Q(\c[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3029_ (.D(_0084_),
    .CLK(net80),
    .Q(\c[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3030_ (.D(_0085_),
    .CLK(net83),
    .Q(\c[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout73 (.I(net79),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout75 (.I(net78),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout78 (.I(net79),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout79 (.I(net96),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout80 (.I(net82),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout81 (.I(net82),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout82 (.I(net86),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout83 (.I(net86),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout84 (.I(net86),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout86 (.I(net95),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout90 (.I(net94),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout91 (.I(net92),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout92 (.I(net94),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout95 (.I(net96),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout96 (.I(net1),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(wb_clk_i),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(wbs_dat_i[19]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(wbs_dat_i[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(wbs_dat_i[20]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input13 (.I(wbs_dat_i[21]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(wbs_dat_i[22]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input15 (.I(wbs_dat_i[23]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(wbs_dat_i[2]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(wbs_dat_i[3]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(wbs_dat_i[4]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input19 (.I(wbs_dat_i[5]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(wb_rst_i),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input20 (.I(wbs_dat_i[6]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input21 (.I(wbs_dat_i[7]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(wbs_dat_i[8]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(wbs_dat_i[9]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input24 (.I(wbs_sel_i[0]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input25 (.I(wbs_sel_i[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input26 (.I(wbs_sel_i[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(wbs_stb_i),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(wbs_we_i),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input29 (.I(y[0]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(wbs_adr_i[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(y[1]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input31 (.I(y[2]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input32 (.I(y[3]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(y[4]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(y[5]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input35 (.I(y[6]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input36 (.I(y[7]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(wbs_adr_i[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(wbs_cyc_i),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(wbs_dat_i[0]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input7 (.I(wbs_dat_i[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input8 (.I(wbs_dat_i[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(wbs_dat_i[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel interp_tri_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(active));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output39 (.I(net39),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output41 (.I(net41),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output43 (.I(net43),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output51 (.I(net51),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output53 (.I(net53),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(x_end[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output58 (.I(net58),
    .Z(x_end[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output59 (.I(net59),
    .Z(x_end[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output60 (.I(net60),
    .Z(x_end[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output61 (.I(net61),
    .Z(x_end[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output62 (.I(net62),
    .Z(x_end[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output63 (.I(net63),
    .Z(x_end[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(x_end[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output65 (.I(net65),
    .Z(x_start[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output66 (.I(net66),
    .Z(x_start[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output67 (.I(net67),
    .Z(x_start[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output68 (.I(net68),
    .Z(x_start[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output69 (.I(net69),
    .Z(x_start[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output70 (.I(net70),
    .Z(x_start[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output71 (.I(net71),
    .Z(x_start[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output72 (.I(net72),
    .Z(x_start[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer1 (.I(_1090_),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(net139),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_0966_),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(_1142_),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(_1439_),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer14 (.I(_1247_),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer15 (.I(net127),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(_1145_),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer17 (.I(_1088_),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer18 (.I(_0966_),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer19 (.I(_1169_),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(_1090_),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer20 (.I(_1087_),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer21 (.I(_1022_),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer22 (.I(_1022_),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer23 (.I(_1167_),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer24 (.I(net138),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer25 (.I(_0313_),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer26 (.I(_1101_),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer27 (.I(_1161_),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer28 (.I(_1158_),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer29 (.I(_1025_),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(_0348_),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_0345_),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_0385_),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(_0376_),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(_0332_),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer8 (.I(_0924_),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(net126),
    .Z(net119));
 assign wbs_dat_o[10] = net97;
 assign wbs_dat_o[11] = net98;
 assign wbs_dat_o[12] = net99;
 assign wbs_dat_o[13] = net100;
 assign wbs_dat_o[14] = net101;
 assign wbs_dat_o[15] = net102;
 assign wbs_dat_o[24] = net103;
 assign wbs_dat_o[25] = net104;
 assign wbs_dat_o[26] = net105;
 assign wbs_dat_o[27] = net106;
 assign wbs_dat_o[28] = net107;
 assign wbs_dat_o[29] = net108;
 assign wbs_dat_o[30] = net109;
 assign wbs_dat_o[31] = net110;
endmodule

