// SPDX-FileCopyrightText: 2022 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module gf180_ram_64x8_wrapper (
	CLK,
	CEN,
	GWEN,
	WEN,
	A,
	D,
	Q
);

input           CLK;
input           CEN;    //Chip Enable
input           GWEN;   //Global Write Enable
input   [7:0]  	WEN;    //Write Enable
input   [5:0]   A;
input   [7:0]  	D;
output	[7:0]	Q;

gf180mcu_fd_ip_sram__sram64x8m8wm1 RAM (
    .CLK(CLK), 
    .CEN(CEN), 
    .GWEN(GWEN), 
    .WEN(WEN), 
    .A(A), 
    .D(D), 
    .Q(Q), 
    .VDD(), 
    .VSS());

endmodule