magic
tech gf180mcuD
magscale 1 5
timestamp 1700139237
<< obsm1 >>
rect 500 500 43686 23788
<< metal2 >>
rect 1872 23988 1928 24388
rect 2222 23988 2278 24388
rect 2672 23988 2728 24388
rect 6722 23988 6778 24388
rect 7072 23988 7128 24388
rect 7272 23988 7328 24388
rect 7497 23988 7553 24388
rect 7722 23988 7778 24388
rect 8022 23988 8078 24388
rect 12122 23988 12178 24388
rect 12522 23988 12578 24388
rect 12872 23988 12928 24388
rect 15472 23988 15528 24388
rect 15972 23988 16028 24388
rect 16372 23988 16428 24388
rect 18422 23988 18478 24388
rect 23284 23988 23340 24388
rect 26472 23988 26528 24388
rect 27322 23988 27378 24388
rect 28172 23988 28228 24388
rect 29622 23988 29678 24388
rect 31672 23988 31728 24388
rect 31872 23988 31928 24388
rect 32472 23988 32528 24388
rect 36522 23988 36578 24388
rect 36872 23988 36928 24388
rect 37072 23988 37128 24388
rect 37272 23988 37328 24388
rect 37472 23988 37528 24388
rect 37822 23988 37878 24388
rect 41922 23988 41978 24388
rect 42322 23988 42378 24388
rect 42672 23988 42728 24388
<< obsm2 >>
rect 500 23958 1842 24052
rect 1958 23958 2192 24052
rect 2308 23958 2642 24052
rect 2758 23958 6692 24052
rect 6808 23958 7042 24052
rect 7158 23958 7242 24052
rect 7358 23958 7467 24052
rect 7583 23958 7692 24052
rect 7808 23958 7992 24052
rect 8108 23958 12092 24052
rect 12208 23958 12492 24052
rect 12608 23958 12842 24052
rect 12958 23958 15442 24052
rect 15558 23958 15942 24052
rect 16058 23958 16342 24052
rect 16458 23958 18392 24052
rect 18508 23958 23254 24052
rect 23370 23958 26442 24052
rect 26558 23958 27292 24052
rect 27408 23958 28142 24052
rect 28258 23958 29592 24052
rect 29708 23958 31642 24052
rect 31758 23958 31842 24052
rect 31958 23958 32442 24052
rect 32558 23958 36492 24052
rect 36608 23958 36842 24052
rect 36958 23958 37042 24052
rect 37158 23958 37242 24052
rect 37358 23958 37442 24052
rect 37558 23958 37792 24052
rect 37908 23958 41892 24052
rect 42008 23958 42292 24052
rect 42408 23958 42642 24052
rect 42758 23958 43686 24052
rect 500 500 43686 23958
<< obsm3 >>
rect 500 500 43686 23788
<< metal4 >>
rect 522 1568 822 22736
rect 922 1568 1222 22736
rect 42863 1568 43163 22736
rect 43263 1568 43563 22736
<< labels >>
rlabel metal2 s 26472 23988 26528 24388 6 A[0]
port 1 nsew signal input
rlabel metal2 s 27322 23988 27378 24388 6 A[1]
port 2 nsew signal input
rlabel metal2 s 28172 23988 28228 24388 6 A[2]
port 3 nsew signal input
rlabel metal2 s 15472 23988 15528 24388 6 A[3]
port 4 nsew signal input
rlabel metal2 s 15972 23988 16028 24388 6 A[4]
port 5 nsew signal input
rlabel metal2 s 16372 23988 16428 24388 6 A[5]
port 6 nsew signal input
rlabel metal2 s 18422 23988 18478 24388 6 CEN
port 7 nsew signal input
rlabel metal2 s 29622 23988 29678 24388 6 CLK
port 8 nsew signal input
rlabel metal2 s 42672 23988 42728 24388 6 D[0]
port 9 nsew signal input
rlabel metal2 s 37472 23988 37528 24388 6 D[1]
port 10 nsew signal input
rlabel metal2 s 36872 23988 36928 24388 6 D[2]
port 11 nsew signal input
rlabel metal2 s 31672 23988 31728 24388 6 D[3]
port 12 nsew signal input
rlabel metal2 s 12872 23988 12928 24388 6 D[4]
port 13 nsew signal input
rlabel metal2 s 7722 23988 7778 24388 6 D[5]
port 14 nsew signal input
rlabel metal2 s 7072 23988 7128 24388 6 D[6]
port 15 nsew signal input
rlabel metal2 s 1872 23988 1928 24388 6 D[7]
port 16 nsew signal input
rlabel metal2 s 23284 23988 23340 24388 6 GWEN
port 17 nsew signal input
rlabel metal2 s 41922 23988 41978 24388 6 Q[0]
port 18 nsew signal output
rlabel metal2 s 37822 23988 37878 24388 6 Q[1]
port 19 nsew signal output
rlabel metal2 s 36522 23988 36578 24388 6 Q[2]
port 20 nsew signal output
rlabel metal2 s 32472 23988 32528 24388 6 Q[3]
port 21 nsew signal output
rlabel metal2 s 12122 23988 12178 24388 6 Q[4]
port 22 nsew signal output
rlabel metal2 s 8022 23988 8078 24388 6 Q[5]
port 23 nsew signal output
rlabel metal2 s 6722 23988 6778 24388 6 Q[6]
port 24 nsew signal output
rlabel metal2 s 2672 23988 2728 24388 6 Q[7]
port 25 nsew signal output
rlabel metal4 s 522 1568 822 22736 6 VDD
port 26 nsew power bidirectional
rlabel metal4 s 42863 1568 43163 22736 6 VDD
port 26 nsew power bidirectional
rlabel metal4 s 922 1568 1222 22736 6 VSS
port 27 nsew ground bidirectional
rlabel metal4 s 43263 1568 43563 22736 6 VSS
port 27 nsew ground bidirectional
rlabel metal2 s 42322 23988 42378 24388 6 WEN[0]
port 28 nsew signal input
rlabel metal2 s 37272 23988 37328 24388 6 WEN[1]
port 29 nsew signal input
rlabel metal2 s 37072 23988 37128 24388 6 WEN[2]
port 30 nsew signal input
rlabel metal2 s 31872 23988 31928 24388 6 WEN[3]
port 31 nsew signal input
rlabel metal2 s 12522 23988 12578 24388 6 WEN[4]
port 32 nsew signal input
rlabel metal2 s 7497 23988 7553 24388 6 WEN[5]
port 33 nsew signal input
rlabel metal2 s 7272 23988 7328 24388 6 WEN[6]
port 34 nsew signal input
rlabel metal2 s 2222 23988 2278 24388 6 WEN[7]
port 35 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44486 24388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2408122
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/gf180_ram_64x8_wrapper/runs/23_11_16_07_53/results/signoff/gf180_ram_64x8_wrapper.magic.gds
string GDS_START 2322632
<< end >>

