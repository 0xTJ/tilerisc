// This is the unpowered netlist.
module tinyrv (clk,
    alu_out_out,
    inst,
    mem_load_out,
    pc,
    pc_next);
 input clk;
 output [31:0] alu_out_out;
 input [31:0] inst;
 input [31:0] mem_load_out;
 input [31:0] pc;
 output [31:0] pc_next;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \reg_file.reg_storage[10][0] ;
 wire \reg_file.reg_storage[10][10] ;
 wire \reg_file.reg_storage[10][11] ;
 wire \reg_file.reg_storage[10][12] ;
 wire \reg_file.reg_storage[10][13] ;
 wire \reg_file.reg_storage[10][14] ;
 wire \reg_file.reg_storage[10][15] ;
 wire \reg_file.reg_storage[10][16] ;
 wire \reg_file.reg_storage[10][17] ;
 wire \reg_file.reg_storage[10][18] ;
 wire \reg_file.reg_storage[10][19] ;
 wire \reg_file.reg_storage[10][1] ;
 wire \reg_file.reg_storage[10][20] ;
 wire \reg_file.reg_storage[10][21] ;
 wire \reg_file.reg_storage[10][22] ;
 wire \reg_file.reg_storage[10][23] ;
 wire \reg_file.reg_storage[10][24] ;
 wire \reg_file.reg_storage[10][25] ;
 wire \reg_file.reg_storage[10][26] ;
 wire \reg_file.reg_storage[10][27] ;
 wire \reg_file.reg_storage[10][28] ;
 wire \reg_file.reg_storage[10][29] ;
 wire \reg_file.reg_storage[10][2] ;
 wire \reg_file.reg_storage[10][30] ;
 wire \reg_file.reg_storage[10][31] ;
 wire \reg_file.reg_storage[10][3] ;
 wire \reg_file.reg_storage[10][4] ;
 wire \reg_file.reg_storage[10][5] ;
 wire \reg_file.reg_storage[10][6] ;
 wire \reg_file.reg_storage[10][7] ;
 wire \reg_file.reg_storage[10][8] ;
 wire \reg_file.reg_storage[10][9] ;
 wire \reg_file.reg_storage[11][0] ;
 wire \reg_file.reg_storage[11][10] ;
 wire \reg_file.reg_storage[11][11] ;
 wire \reg_file.reg_storage[11][12] ;
 wire \reg_file.reg_storage[11][13] ;
 wire \reg_file.reg_storage[11][14] ;
 wire \reg_file.reg_storage[11][15] ;
 wire \reg_file.reg_storage[11][16] ;
 wire \reg_file.reg_storage[11][17] ;
 wire \reg_file.reg_storage[11][18] ;
 wire \reg_file.reg_storage[11][19] ;
 wire \reg_file.reg_storage[11][1] ;
 wire \reg_file.reg_storage[11][20] ;
 wire \reg_file.reg_storage[11][21] ;
 wire \reg_file.reg_storage[11][22] ;
 wire \reg_file.reg_storage[11][23] ;
 wire \reg_file.reg_storage[11][24] ;
 wire \reg_file.reg_storage[11][25] ;
 wire \reg_file.reg_storage[11][26] ;
 wire \reg_file.reg_storage[11][27] ;
 wire \reg_file.reg_storage[11][28] ;
 wire \reg_file.reg_storage[11][29] ;
 wire \reg_file.reg_storage[11][2] ;
 wire \reg_file.reg_storage[11][30] ;
 wire \reg_file.reg_storage[11][31] ;
 wire \reg_file.reg_storage[11][3] ;
 wire \reg_file.reg_storage[11][4] ;
 wire \reg_file.reg_storage[11][5] ;
 wire \reg_file.reg_storage[11][6] ;
 wire \reg_file.reg_storage[11][7] ;
 wire \reg_file.reg_storage[11][8] ;
 wire \reg_file.reg_storage[11][9] ;
 wire \reg_file.reg_storage[12][0] ;
 wire \reg_file.reg_storage[12][10] ;
 wire \reg_file.reg_storage[12][11] ;
 wire \reg_file.reg_storage[12][12] ;
 wire \reg_file.reg_storage[12][13] ;
 wire \reg_file.reg_storage[12][14] ;
 wire \reg_file.reg_storage[12][15] ;
 wire \reg_file.reg_storage[12][16] ;
 wire \reg_file.reg_storage[12][17] ;
 wire \reg_file.reg_storage[12][18] ;
 wire \reg_file.reg_storage[12][19] ;
 wire \reg_file.reg_storage[12][1] ;
 wire \reg_file.reg_storage[12][20] ;
 wire \reg_file.reg_storage[12][21] ;
 wire \reg_file.reg_storage[12][22] ;
 wire \reg_file.reg_storage[12][23] ;
 wire \reg_file.reg_storage[12][24] ;
 wire \reg_file.reg_storage[12][25] ;
 wire \reg_file.reg_storage[12][26] ;
 wire \reg_file.reg_storage[12][27] ;
 wire \reg_file.reg_storage[12][28] ;
 wire \reg_file.reg_storage[12][29] ;
 wire \reg_file.reg_storage[12][2] ;
 wire \reg_file.reg_storage[12][30] ;
 wire \reg_file.reg_storage[12][31] ;
 wire \reg_file.reg_storage[12][3] ;
 wire \reg_file.reg_storage[12][4] ;
 wire \reg_file.reg_storage[12][5] ;
 wire \reg_file.reg_storage[12][6] ;
 wire \reg_file.reg_storage[12][7] ;
 wire \reg_file.reg_storage[12][8] ;
 wire \reg_file.reg_storage[12][9] ;
 wire \reg_file.reg_storage[13][0] ;
 wire \reg_file.reg_storage[13][10] ;
 wire \reg_file.reg_storage[13][11] ;
 wire \reg_file.reg_storage[13][12] ;
 wire \reg_file.reg_storage[13][13] ;
 wire \reg_file.reg_storage[13][14] ;
 wire \reg_file.reg_storage[13][15] ;
 wire \reg_file.reg_storage[13][16] ;
 wire \reg_file.reg_storage[13][17] ;
 wire \reg_file.reg_storage[13][18] ;
 wire \reg_file.reg_storage[13][19] ;
 wire \reg_file.reg_storage[13][1] ;
 wire \reg_file.reg_storage[13][20] ;
 wire \reg_file.reg_storage[13][21] ;
 wire \reg_file.reg_storage[13][22] ;
 wire \reg_file.reg_storage[13][23] ;
 wire \reg_file.reg_storage[13][24] ;
 wire \reg_file.reg_storage[13][25] ;
 wire \reg_file.reg_storage[13][26] ;
 wire \reg_file.reg_storage[13][27] ;
 wire \reg_file.reg_storage[13][28] ;
 wire \reg_file.reg_storage[13][29] ;
 wire \reg_file.reg_storage[13][2] ;
 wire \reg_file.reg_storage[13][30] ;
 wire \reg_file.reg_storage[13][31] ;
 wire \reg_file.reg_storage[13][3] ;
 wire \reg_file.reg_storage[13][4] ;
 wire \reg_file.reg_storage[13][5] ;
 wire \reg_file.reg_storage[13][6] ;
 wire \reg_file.reg_storage[13][7] ;
 wire \reg_file.reg_storage[13][8] ;
 wire \reg_file.reg_storage[13][9] ;
 wire \reg_file.reg_storage[14][0] ;
 wire \reg_file.reg_storage[14][10] ;
 wire \reg_file.reg_storage[14][11] ;
 wire \reg_file.reg_storage[14][12] ;
 wire \reg_file.reg_storage[14][13] ;
 wire \reg_file.reg_storage[14][14] ;
 wire \reg_file.reg_storage[14][15] ;
 wire \reg_file.reg_storage[14][16] ;
 wire \reg_file.reg_storage[14][17] ;
 wire \reg_file.reg_storage[14][18] ;
 wire \reg_file.reg_storage[14][19] ;
 wire \reg_file.reg_storage[14][1] ;
 wire \reg_file.reg_storage[14][20] ;
 wire \reg_file.reg_storage[14][21] ;
 wire \reg_file.reg_storage[14][22] ;
 wire \reg_file.reg_storage[14][23] ;
 wire \reg_file.reg_storage[14][24] ;
 wire \reg_file.reg_storage[14][25] ;
 wire \reg_file.reg_storage[14][26] ;
 wire \reg_file.reg_storage[14][27] ;
 wire \reg_file.reg_storage[14][28] ;
 wire \reg_file.reg_storage[14][29] ;
 wire \reg_file.reg_storage[14][2] ;
 wire \reg_file.reg_storage[14][30] ;
 wire \reg_file.reg_storage[14][31] ;
 wire \reg_file.reg_storage[14][3] ;
 wire \reg_file.reg_storage[14][4] ;
 wire \reg_file.reg_storage[14][5] ;
 wire \reg_file.reg_storage[14][6] ;
 wire \reg_file.reg_storage[14][7] ;
 wire \reg_file.reg_storage[14][8] ;
 wire \reg_file.reg_storage[14][9] ;
 wire \reg_file.reg_storage[15][0] ;
 wire \reg_file.reg_storage[15][10] ;
 wire \reg_file.reg_storage[15][11] ;
 wire \reg_file.reg_storage[15][12] ;
 wire \reg_file.reg_storage[15][13] ;
 wire \reg_file.reg_storage[15][14] ;
 wire \reg_file.reg_storage[15][15] ;
 wire \reg_file.reg_storage[15][16] ;
 wire \reg_file.reg_storage[15][17] ;
 wire \reg_file.reg_storage[15][18] ;
 wire \reg_file.reg_storage[15][19] ;
 wire \reg_file.reg_storage[15][1] ;
 wire \reg_file.reg_storage[15][20] ;
 wire \reg_file.reg_storage[15][21] ;
 wire \reg_file.reg_storage[15][22] ;
 wire \reg_file.reg_storage[15][23] ;
 wire \reg_file.reg_storage[15][24] ;
 wire \reg_file.reg_storage[15][25] ;
 wire \reg_file.reg_storage[15][26] ;
 wire \reg_file.reg_storage[15][27] ;
 wire \reg_file.reg_storage[15][28] ;
 wire \reg_file.reg_storage[15][29] ;
 wire \reg_file.reg_storage[15][2] ;
 wire \reg_file.reg_storage[15][30] ;
 wire \reg_file.reg_storage[15][31] ;
 wire \reg_file.reg_storage[15][3] ;
 wire \reg_file.reg_storage[15][4] ;
 wire \reg_file.reg_storage[15][5] ;
 wire \reg_file.reg_storage[15][6] ;
 wire \reg_file.reg_storage[15][7] ;
 wire \reg_file.reg_storage[15][8] ;
 wire \reg_file.reg_storage[15][9] ;
 wire \reg_file.reg_storage[1][0] ;
 wire \reg_file.reg_storage[1][10] ;
 wire \reg_file.reg_storage[1][11] ;
 wire \reg_file.reg_storage[1][12] ;
 wire \reg_file.reg_storage[1][13] ;
 wire \reg_file.reg_storage[1][14] ;
 wire \reg_file.reg_storage[1][15] ;
 wire \reg_file.reg_storage[1][16] ;
 wire \reg_file.reg_storage[1][17] ;
 wire \reg_file.reg_storage[1][18] ;
 wire \reg_file.reg_storage[1][19] ;
 wire \reg_file.reg_storage[1][1] ;
 wire \reg_file.reg_storage[1][20] ;
 wire \reg_file.reg_storage[1][21] ;
 wire \reg_file.reg_storage[1][22] ;
 wire \reg_file.reg_storage[1][23] ;
 wire \reg_file.reg_storage[1][24] ;
 wire \reg_file.reg_storage[1][25] ;
 wire \reg_file.reg_storage[1][26] ;
 wire \reg_file.reg_storage[1][27] ;
 wire \reg_file.reg_storage[1][28] ;
 wire \reg_file.reg_storage[1][29] ;
 wire \reg_file.reg_storage[1][2] ;
 wire \reg_file.reg_storage[1][30] ;
 wire \reg_file.reg_storage[1][31] ;
 wire \reg_file.reg_storage[1][3] ;
 wire \reg_file.reg_storage[1][4] ;
 wire \reg_file.reg_storage[1][5] ;
 wire \reg_file.reg_storage[1][6] ;
 wire \reg_file.reg_storage[1][7] ;
 wire \reg_file.reg_storage[1][8] ;
 wire \reg_file.reg_storage[1][9] ;
 wire \reg_file.reg_storage[2][0] ;
 wire \reg_file.reg_storage[2][10] ;
 wire \reg_file.reg_storage[2][11] ;
 wire \reg_file.reg_storage[2][12] ;
 wire \reg_file.reg_storage[2][13] ;
 wire \reg_file.reg_storage[2][14] ;
 wire \reg_file.reg_storage[2][15] ;
 wire \reg_file.reg_storage[2][16] ;
 wire \reg_file.reg_storage[2][17] ;
 wire \reg_file.reg_storage[2][18] ;
 wire \reg_file.reg_storage[2][19] ;
 wire \reg_file.reg_storage[2][1] ;
 wire \reg_file.reg_storage[2][20] ;
 wire \reg_file.reg_storage[2][21] ;
 wire \reg_file.reg_storage[2][22] ;
 wire \reg_file.reg_storage[2][23] ;
 wire \reg_file.reg_storage[2][24] ;
 wire \reg_file.reg_storage[2][25] ;
 wire \reg_file.reg_storage[2][26] ;
 wire \reg_file.reg_storage[2][27] ;
 wire \reg_file.reg_storage[2][28] ;
 wire \reg_file.reg_storage[2][29] ;
 wire \reg_file.reg_storage[2][2] ;
 wire \reg_file.reg_storage[2][30] ;
 wire \reg_file.reg_storage[2][31] ;
 wire \reg_file.reg_storage[2][3] ;
 wire \reg_file.reg_storage[2][4] ;
 wire \reg_file.reg_storage[2][5] ;
 wire \reg_file.reg_storage[2][6] ;
 wire \reg_file.reg_storage[2][7] ;
 wire \reg_file.reg_storage[2][8] ;
 wire \reg_file.reg_storage[2][9] ;
 wire \reg_file.reg_storage[3][0] ;
 wire \reg_file.reg_storage[3][10] ;
 wire \reg_file.reg_storage[3][11] ;
 wire \reg_file.reg_storage[3][12] ;
 wire \reg_file.reg_storage[3][13] ;
 wire \reg_file.reg_storage[3][14] ;
 wire \reg_file.reg_storage[3][15] ;
 wire \reg_file.reg_storage[3][16] ;
 wire \reg_file.reg_storage[3][17] ;
 wire \reg_file.reg_storage[3][18] ;
 wire \reg_file.reg_storage[3][19] ;
 wire \reg_file.reg_storage[3][1] ;
 wire \reg_file.reg_storage[3][20] ;
 wire \reg_file.reg_storage[3][21] ;
 wire \reg_file.reg_storage[3][22] ;
 wire \reg_file.reg_storage[3][23] ;
 wire \reg_file.reg_storage[3][24] ;
 wire \reg_file.reg_storage[3][25] ;
 wire \reg_file.reg_storage[3][26] ;
 wire \reg_file.reg_storage[3][27] ;
 wire \reg_file.reg_storage[3][28] ;
 wire \reg_file.reg_storage[3][29] ;
 wire \reg_file.reg_storage[3][2] ;
 wire \reg_file.reg_storage[3][30] ;
 wire \reg_file.reg_storage[3][31] ;
 wire \reg_file.reg_storage[3][3] ;
 wire \reg_file.reg_storage[3][4] ;
 wire \reg_file.reg_storage[3][5] ;
 wire \reg_file.reg_storage[3][6] ;
 wire \reg_file.reg_storage[3][7] ;
 wire \reg_file.reg_storage[3][8] ;
 wire \reg_file.reg_storage[3][9] ;
 wire \reg_file.reg_storage[4][0] ;
 wire \reg_file.reg_storage[4][10] ;
 wire \reg_file.reg_storage[4][11] ;
 wire \reg_file.reg_storage[4][12] ;
 wire \reg_file.reg_storage[4][13] ;
 wire \reg_file.reg_storage[4][14] ;
 wire \reg_file.reg_storage[4][15] ;
 wire \reg_file.reg_storage[4][16] ;
 wire \reg_file.reg_storage[4][17] ;
 wire \reg_file.reg_storage[4][18] ;
 wire \reg_file.reg_storage[4][19] ;
 wire \reg_file.reg_storage[4][1] ;
 wire \reg_file.reg_storage[4][20] ;
 wire \reg_file.reg_storage[4][21] ;
 wire \reg_file.reg_storage[4][22] ;
 wire \reg_file.reg_storage[4][23] ;
 wire \reg_file.reg_storage[4][24] ;
 wire \reg_file.reg_storage[4][25] ;
 wire \reg_file.reg_storage[4][26] ;
 wire \reg_file.reg_storage[4][27] ;
 wire \reg_file.reg_storage[4][28] ;
 wire \reg_file.reg_storage[4][29] ;
 wire \reg_file.reg_storage[4][2] ;
 wire \reg_file.reg_storage[4][30] ;
 wire \reg_file.reg_storage[4][31] ;
 wire \reg_file.reg_storage[4][3] ;
 wire \reg_file.reg_storage[4][4] ;
 wire \reg_file.reg_storage[4][5] ;
 wire \reg_file.reg_storage[4][6] ;
 wire \reg_file.reg_storage[4][7] ;
 wire \reg_file.reg_storage[4][8] ;
 wire \reg_file.reg_storage[4][9] ;
 wire \reg_file.reg_storage[5][0] ;
 wire \reg_file.reg_storage[5][10] ;
 wire \reg_file.reg_storage[5][11] ;
 wire \reg_file.reg_storage[5][12] ;
 wire \reg_file.reg_storage[5][13] ;
 wire \reg_file.reg_storage[5][14] ;
 wire \reg_file.reg_storage[5][15] ;
 wire \reg_file.reg_storage[5][16] ;
 wire \reg_file.reg_storage[5][17] ;
 wire \reg_file.reg_storage[5][18] ;
 wire \reg_file.reg_storage[5][19] ;
 wire \reg_file.reg_storage[5][1] ;
 wire \reg_file.reg_storage[5][20] ;
 wire \reg_file.reg_storage[5][21] ;
 wire \reg_file.reg_storage[5][22] ;
 wire \reg_file.reg_storage[5][23] ;
 wire \reg_file.reg_storage[5][24] ;
 wire \reg_file.reg_storage[5][25] ;
 wire \reg_file.reg_storage[5][26] ;
 wire \reg_file.reg_storage[5][27] ;
 wire \reg_file.reg_storage[5][28] ;
 wire \reg_file.reg_storage[5][29] ;
 wire \reg_file.reg_storage[5][2] ;
 wire \reg_file.reg_storage[5][30] ;
 wire \reg_file.reg_storage[5][31] ;
 wire \reg_file.reg_storage[5][3] ;
 wire \reg_file.reg_storage[5][4] ;
 wire \reg_file.reg_storage[5][5] ;
 wire \reg_file.reg_storage[5][6] ;
 wire \reg_file.reg_storage[5][7] ;
 wire \reg_file.reg_storage[5][8] ;
 wire \reg_file.reg_storage[5][9] ;
 wire \reg_file.reg_storage[6][0] ;
 wire \reg_file.reg_storage[6][10] ;
 wire \reg_file.reg_storage[6][11] ;
 wire \reg_file.reg_storage[6][12] ;
 wire \reg_file.reg_storage[6][13] ;
 wire \reg_file.reg_storage[6][14] ;
 wire \reg_file.reg_storage[6][15] ;
 wire \reg_file.reg_storage[6][16] ;
 wire \reg_file.reg_storage[6][17] ;
 wire \reg_file.reg_storage[6][18] ;
 wire \reg_file.reg_storage[6][19] ;
 wire \reg_file.reg_storage[6][1] ;
 wire \reg_file.reg_storage[6][20] ;
 wire \reg_file.reg_storage[6][21] ;
 wire \reg_file.reg_storage[6][22] ;
 wire \reg_file.reg_storage[6][23] ;
 wire \reg_file.reg_storage[6][24] ;
 wire \reg_file.reg_storage[6][25] ;
 wire \reg_file.reg_storage[6][26] ;
 wire \reg_file.reg_storage[6][27] ;
 wire \reg_file.reg_storage[6][28] ;
 wire \reg_file.reg_storage[6][29] ;
 wire \reg_file.reg_storage[6][2] ;
 wire \reg_file.reg_storage[6][30] ;
 wire \reg_file.reg_storage[6][31] ;
 wire \reg_file.reg_storage[6][3] ;
 wire \reg_file.reg_storage[6][4] ;
 wire \reg_file.reg_storage[6][5] ;
 wire \reg_file.reg_storage[6][6] ;
 wire \reg_file.reg_storage[6][7] ;
 wire \reg_file.reg_storage[6][8] ;
 wire \reg_file.reg_storage[6][9] ;
 wire \reg_file.reg_storage[7][0] ;
 wire \reg_file.reg_storage[7][10] ;
 wire \reg_file.reg_storage[7][11] ;
 wire \reg_file.reg_storage[7][12] ;
 wire \reg_file.reg_storage[7][13] ;
 wire \reg_file.reg_storage[7][14] ;
 wire \reg_file.reg_storage[7][15] ;
 wire \reg_file.reg_storage[7][16] ;
 wire \reg_file.reg_storage[7][17] ;
 wire \reg_file.reg_storage[7][18] ;
 wire \reg_file.reg_storage[7][19] ;
 wire \reg_file.reg_storage[7][1] ;
 wire \reg_file.reg_storage[7][20] ;
 wire \reg_file.reg_storage[7][21] ;
 wire \reg_file.reg_storage[7][22] ;
 wire \reg_file.reg_storage[7][23] ;
 wire \reg_file.reg_storage[7][24] ;
 wire \reg_file.reg_storage[7][25] ;
 wire \reg_file.reg_storage[7][26] ;
 wire \reg_file.reg_storage[7][27] ;
 wire \reg_file.reg_storage[7][28] ;
 wire \reg_file.reg_storage[7][29] ;
 wire \reg_file.reg_storage[7][2] ;
 wire \reg_file.reg_storage[7][30] ;
 wire \reg_file.reg_storage[7][31] ;
 wire \reg_file.reg_storage[7][3] ;
 wire \reg_file.reg_storage[7][4] ;
 wire \reg_file.reg_storage[7][5] ;
 wire \reg_file.reg_storage[7][6] ;
 wire \reg_file.reg_storage[7][7] ;
 wire \reg_file.reg_storage[7][8] ;
 wire \reg_file.reg_storage[7][9] ;
 wire \reg_file.reg_storage[8][0] ;
 wire \reg_file.reg_storage[8][10] ;
 wire \reg_file.reg_storage[8][11] ;
 wire \reg_file.reg_storage[8][12] ;
 wire \reg_file.reg_storage[8][13] ;
 wire \reg_file.reg_storage[8][14] ;
 wire \reg_file.reg_storage[8][15] ;
 wire \reg_file.reg_storage[8][16] ;
 wire \reg_file.reg_storage[8][17] ;
 wire \reg_file.reg_storage[8][18] ;
 wire \reg_file.reg_storage[8][19] ;
 wire \reg_file.reg_storage[8][1] ;
 wire \reg_file.reg_storage[8][20] ;
 wire \reg_file.reg_storage[8][21] ;
 wire \reg_file.reg_storage[8][22] ;
 wire \reg_file.reg_storage[8][23] ;
 wire \reg_file.reg_storage[8][24] ;
 wire \reg_file.reg_storage[8][25] ;
 wire \reg_file.reg_storage[8][26] ;
 wire \reg_file.reg_storage[8][27] ;
 wire \reg_file.reg_storage[8][28] ;
 wire \reg_file.reg_storage[8][29] ;
 wire \reg_file.reg_storage[8][2] ;
 wire \reg_file.reg_storage[8][30] ;
 wire \reg_file.reg_storage[8][31] ;
 wire \reg_file.reg_storage[8][3] ;
 wire \reg_file.reg_storage[8][4] ;
 wire \reg_file.reg_storage[8][5] ;
 wire \reg_file.reg_storage[8][6] ;
 wire \reg_file.reg_storage[8][7] ;
 wire \reg_file.reg_storage[8][8] ;
 wire \reg_file.reg_storage[8][9] ;
 wire \reg_file.reg_storage[9][0] ;
 wire \reg_file.reg_storage[9][10] ;
 wire \reg_file.reg_storage[9][11] ;
 wire \reg_file.reg_storage[9][12] ;
 wire \reg_file.reg_storage[9][13] ;
 wire \reg_file.reg_storage[9][14] ;
 wire \reg_file.reg_storage[9][15] ;
 wire \reg_file.reg_storage[9][16] ;
 wire \reg_file.reg_storage[9][17] ;
 wire \reg_file.reg_storage[9][18] ;
 wire \reg_file.reg_storage[9][19] ;
 wire \reg_file.reg_storage[9][1] ;
 wire \reg_file.reg_storage[9][20] ;
 wire \reg_file.reg_storage[9][21] ;
 wire \reg_file.reg_storage[9][22] ;
 wire \reg_file.reg_storage[9][23] ;
 wire \reg_file.reg_storage[9][24] ;
 wire \reg_file.reg_storage[9][25] ;
 wire \reg_file.reg_storage[9][26] ;
 wire \reg_file.reg_storage[9][27] ;
 wire \reg_file.reg_storage[9][28] ;
 wire \reg_file.reg_storage[9][29] ;
 wire \reg_file.reg_storage[9][2] ;
 wire \reg_file.reg_storage[9][30] ;
 wire \reg_file.reg_storage[9][31] ;
 wire \reg_file.reg_storage[9][3] ;
 wire \reg_file.reg_storage[9][4] ;
 wire \reg_file.reg_storage[9][5] ;
 wire \reg_file.reg_storage[9][6] ;
 wire \reg_file.reg_storage[9][7] ;
 wire \reg_file.reg_storage[9][8] ;
 wire \reg_file.reg_storage[9][9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A3 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__S0 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__S1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__I (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__B (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__I (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__I1 (.I(\reg_file.reg_storage[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__I2 (.I(\reg_file.reg_storage[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__S0 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__S1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I0 (.I(\reg_file.reg_storage[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I3 (.I(\reg_file.reg_storage[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__S0 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__S1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__S0 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__S1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__B2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A3 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A3 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A4 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__S0 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__S1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I1 (.I(\reg_file.reg_storage[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I2 (.I(\reg_file.reg_storage[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__S0 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__S1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__I0 (.I(\reg_file.reg_storage[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__I3 (.I(\reg_file.reg_storage[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__S0 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__S1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__S0 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__S1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__B2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I0 (.I(\reg_file.reg_storage[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I1 (.I(\reg_file.reg_storage[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__S (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I0 (.I(\reg_file.reg_storage[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__S (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I2 (.I(\reg_file.reg_storage[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I3 (.I(\reg_file.reg_storage[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__S0 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__S1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__C (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__S0 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__S1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I1 (.I(\reg_file.reg_storage[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__S0 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__S1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__C (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__I2 (.I(\reg_file.reg_storage[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__I3 (.I(\reg_file.reg_storage[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__S0 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__S1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(\reg_file.reg_storage[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(\reg_file.reg_storage[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(\reg_file.reg_storage[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__B (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__I (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__S1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I1 (.I(\reg_file.reg_storage[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__S0 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__S1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__S0 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__S1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__B1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I0 (.I(\reg_file.reg_storage[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__S (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__S (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__S0 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__S1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__C (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I0 (.I(\reg_file.reg_storage[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I1 (.I(\reg_file.reg_storage[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I2 (.I(\reg_file.reg_storage[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I3 (.I(\reg_file.reg_storage[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__S0 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__S1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I0 (.I(\reg_file.reg_storage[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I3 (.I(\reg_file.reg_storage[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__S0 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__S1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__C (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__B1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__S0 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__S1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(\reg_file.reg_storage[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__B (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I0 (.I(\reg_file.reg_storage[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I1 (.I(\reg_file.reg_storage[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I2 (.I(\reg_file.reg_storage[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I3 (.I(\reg_file.reg_storage[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__S0 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__S1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I0 (.I(\reg_file.reg_storage[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I3 (.I(\reg_file.reg_storage[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__S0 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__S1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__S0 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__S1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__S0 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__S1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__B (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__S0 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__S1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__S0 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__S1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__S0 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__S1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__S0 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__S1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__B (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S0 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__S0 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__S1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__S0 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__S1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I2 (.I(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I3 (.I(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__S1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__B (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__S0 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__S1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__S0 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__S1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__S0 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__S1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__B2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I2 (.I(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I3 (.I(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__S0 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__S1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__I (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__S0 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__S1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__S0 (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__S1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__S0 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__S1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__B1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__S (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__S (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I2 (.I(\reg_file.reg_storage[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I3 (.I(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__S0 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__S1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__C (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__S0 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__S1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__I1 (.I(\reg_file.reg_storage[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__S0 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__C (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__I (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I2 (.I(\reg_file.reg_storage[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I3 (.I(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__S0 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__S1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__B (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__S0 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__S1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__I1 (.I(\reg_file.reg_storage[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__S0 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__S1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__S0 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__S1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__B1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__I0 (.I(\reg_file.reg_storage[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__S (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__S (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I2 (.I(\reg_file.reg_storage[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I3 (.I(\reg_file.reg_storage[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__S0 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__S1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__C (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I1 (.I(\reg_file.reg_storage[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__S0 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__S1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__I0 (.I(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__I1 (.I(\reg_file.reg_storage[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__I3 (.I(\reg_file.reg_storage[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__S0 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__S1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__C (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__B1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I2 (.I(\reg_file.reg_storage[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I3 (.I(\reg_file.reg_storage[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__S0 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__S1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(\reg_file.reg_storage[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__B (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__I1 (.I(\reg_file.reg_storage[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__S0 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__S1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I0 (.I(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I1 (.I(\reg_file.reg_storage[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I3 (.I(\reg_file.reg_storage[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__S0 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__S1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__S0 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__S1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__I2 (.I(\reg_file.reg_storage[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__S0 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(\reg_file.reg_storage[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(\reg_file.reg_storage[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__S0 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I1 (.I(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I2 (.I(\reg_file.reg_storage[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__S0 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I0 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I3 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__S0 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__S1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__B1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I2 (.I(\reg_file.reg_storage[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__S0 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(\reg_file.reg_storage[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(\reg_file.reg_storage[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__S0 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__S1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I1 (.I(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I2 (.I(\reg_file.reg_storage[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__S0 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__S1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__S0 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__S1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__B2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I0 (.I(\reg_file.reg_storage[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I1 (.I(\reg_file.reg_storage[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I0 (.I(\reg_file.reg_storage[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__S (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__I2 (.I(\reg_file.reg_storage[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__S0 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__S1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__C (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__S0 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__S1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I1 (.I(\reg_file.reg_storage[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__S0 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__C (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I2 (.I(\reg_file.reg_storage[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__S0 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__S1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(\reg_file.reg_storage[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__I (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(\reg_file.reg_storage[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(\reg_file.reg_storage[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__B (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__S0 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I1 (.I(\reg_file.reg_storage[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__S0 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__S1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__S0 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__S1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__B1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__B2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A3 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__I1 (.I(\reg_file.reg_storage[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__C (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I3 (.I(\reg_file.reg_storage[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__S0 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__C (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__B1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I1 (.I(\reg_file.reg_storage[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__S0 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__S1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I3 (.I(\reg_file.reg_storage[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__S0 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__S1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__S0 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__S1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__S0 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__S1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__S0 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__S1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__B (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__S0 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__S1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__S0 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__S1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__S0 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__S1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__B1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__S (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__S0 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__S1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__S0 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__S1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__S0 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__S1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A4 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__S (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I0 (.I(\reg_file.reg_storage[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I1 (.I(\reg_file.reg_storage[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__S1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__S0 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__S1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__S0 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__S (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I0 (.I(\reg_file.reg_storage[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I1 (.I(\reg_file.reg_storage[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__S0 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__S1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__B (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__S0 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__S0 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I3 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__S0 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__S1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__B2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I2 (.I(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I3 (.I(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__S0 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__S1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(\reg_file.reg_storage[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(\reg_file.reg_storage[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__B (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__S0 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__S1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I1 (.I(\reg_file.reg_storage[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I2 (.I(\reg_file.reg_storage[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__S0 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__S1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__S1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__B2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I2 (.I(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I3 (.I(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__S0 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__S1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A2 (.I(\reg_file.reg_storage[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(\reg_file.reg_storage[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__B (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__S1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I1 (.I(\reg_file.reg_storage[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I2 (.I(\reg_file.reg_storage[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__S1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__S0 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__S1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__B1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I0 (.I(\reg_file.reg_storage[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I1 (.I(\reg_file.reg_storage[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I0 (.I(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__S (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I2 (.I(\reg_file.reg_storage[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I3 (.I(\reg_file.reg_storage[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__S1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__C (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__S0 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__S1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I1 (.I(\reg_file.reg_storage[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I2 (.I(\reg_file.reg_storage[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__S1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__C (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I2 (.I(\reg_file.reg_storage[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I3 (.I(\reg_file.reg_storage[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__S1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__I (.I(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(\reg_file.reg_storage[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(\reg_file.reg_storage[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__B (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__S0 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__S1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I1 (.I(\reg_file.reg_storage[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I2 (.I(\reg_file.reg_storage[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__S1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__S0 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__S1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__S0 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__S1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__I (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__B (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__S0 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__S1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__S0 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__S1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__S0 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__S1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__B2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__S0 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__S1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__B (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__S0 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__S1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__S0 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__S1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__S0 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__S1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__B1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__B1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__I (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__B2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__I (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__I (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__I (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__S0 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__S1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(\reg_file.reg_storage[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__B (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__S0 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__S1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__S0 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__S1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__I (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__S0 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__S1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__I (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__S0 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__S1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__I (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__S0 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__S1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__S0 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__S1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I3 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__S0 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__S1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__B2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__I (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__I1 (.I(\reg_file.reg_storage[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__S1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__B (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__S (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__S0 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__S1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__S0 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__S1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__S (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__S0 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__S1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__B (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__S0 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__S0 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__S0 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__S1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__S0 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__S1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__B (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__S0 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__S1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I0 (.I(\reg_file.reg_storage[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__S0 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__S1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__S0 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__S1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__S0 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__S1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__B (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__I0 (.I(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__I2 (.I(\reg_file.reg_storage[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__I3 (.I(\reg_file.reg_storage[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__S0 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__S1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__I0 (.I(\reg_file.reg_storage[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__I3 (.I(\reg_file.reg_storage[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__S0 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__S1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__S0 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__S1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__B2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__I (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__B (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I0 (.I(\reg_file.reg_storage[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I1 (.I(\reg_file.reg_storage[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__S0 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__S1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__B (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I0 (.I(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I1 (.I(\reg_file.reg_storage[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I2 (.I(\reg_file.reg_storage[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I3 (.I(\reg_file.reg_storage[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__S0 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__S1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I0 (.I(\reg_file.reg_storage[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I3 (.I(\reg_file.reg_storage[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__S0 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__S1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__S0 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__S1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__B2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__S0 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__S1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(\reg_file.reg_storage[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__B (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__S1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__S0 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__S1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__S0 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__S1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__B2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__S (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I0 (.I(\reg_file.reg_storage[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I1 (.I(\reg_file.reg_storage[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__S0 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__S1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__I2 (.I(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__S0 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__S1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I0 (.I(\reg_file.reg_storage[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I3 (.I(\reg_file.reg_storage[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S0 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__S (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__S (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__S0 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__S1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I2 (.I(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__S0 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__S1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I0 (.I(\reg_file.reg_storage[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I3 (.I(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__S0 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__S1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__S (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__S (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__S0 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__S1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__B (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__I1 (.I(\reg_file.reg_storage[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__I2 (.I(\reg_file.reg_storage[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__S0 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__S1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I0 (.I(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I3 (.I(\reg_file.reg_storage[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__S0 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__S1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__S0 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__S1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__B2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I0 (.I(\reg_file.reg_storage[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I1 (.I(\reg_file.reg_storage[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__S0 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__S1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__C (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__B (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__B (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I0 (.I(\reg_file.reg_storage[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I1 (.I(\reg_file.reg_storage[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I2 (.I(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I3 (.I(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__S0 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__S1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I0 (.I(\reg_file.reg_storage[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I1 (.I(\reg_file.reg_storage[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I3 (.I(\reg_file.reg_storage[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__S0 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__S1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__B (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__B (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__I0 (.I(\reg_file.reg_storage[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__S (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I0 (.I(\reg_file.reg_storage[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I1 (.I(\reg_file.reg_storage[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__S0 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__S1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__S0 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__S0 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__S1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__S (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A2 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__S (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I0 (.I(\reg_file.reg_storage[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__S0 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__S1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__B (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I2 (.I(\reg_file.reg_storage[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__S0 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__S1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I0 (.I(\reg_file.reg_storage[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__S0 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__S1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__S0 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__S1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__B2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__S0 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__S1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__B (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I2 (.I(\reg_file.reg_storage[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__S0 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__S1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I0 (.I(\reg_file.reg_storage[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I3 (.I(\reg_file.reg_storage[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__S0 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__S1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__S0 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__S1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I0 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__S0 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__S1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__B (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__S0 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__S1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__S0 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__S1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I3 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__S0 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__S1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I0 (.I(\reg_file.reg_storage[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__S (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__S (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S0 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__C (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I1 (.I(\reg_file.reg_storage[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I2 (.I(\reg_file.reg_storage[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__S0 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__S1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I0 (.I(\reg_file.reg_storage[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I3 (.I(\reg_file.reg_storage[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__S0 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__S1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__C (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I0 (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__S (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I0 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__S (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__S (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__I (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__B2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A3 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__B (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__S0 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__S1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__B (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__I1 (.I(\reg_file.reg_storage[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__I2 (.I(\reg_file.reg_storage[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__S0 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__S1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__I0 (.I(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__I3 (.I(\reg_file.reg_storage[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__S0 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__S1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__S0 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__S1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__B1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__S (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__S (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__S (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__B (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__S (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__S (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__I (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__S (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I0 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__S (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__I (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__I (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__B (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__I (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I0 (.I(\reg_file.reg_storage[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I1 (.I(\reg_file.reg_storage[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__S0 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__S1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__I (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__I (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(\reg_file.reg_storage[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__B (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__S0 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__S1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__S0 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__S1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__I (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I1 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I3 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__S0 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__S1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__B2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__I (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__B (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__C (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__I (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I0 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__S (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__S (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__I1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__S (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I0 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__B2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__I0 (.I(\reg_file.reg_storage[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__I1 (.I(\reg_file.reg_storage[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__S0 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__S1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__B (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I0 (.I(\reg_file.reg_storage[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I1 (.I(\reg_file.reg_storage[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I2 (.I(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I3 (.I(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I0 (.I(\reg_file.reg_storage[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I1 (.I(\reg_file.reg_storage[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I3 (.I(\reg_file.reg_storage[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__S1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__I1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__S0 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__S1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__B1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__B (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__I (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__I (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__B (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__I (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__S (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__S (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__I (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__I (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__S (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__S (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__I (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A4 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__S0 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__S1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__B (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__I2 (.I(\reg_file.reg_storage[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__S0 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__S1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I0 (.I(\reg_file.reg_storage[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I3 (.I(\reg_file.reg_storage[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__S0 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__S1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__I1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__S0 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__S1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__B1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__B (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I0 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__S (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__S (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A3 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__I (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__I (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__C (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I0 (.I(\reg_file.reg_storage[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__S0 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__S1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__I (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__B (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I2 (.I(\reg_file.reg_storage[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__S0 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__S1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__I0 (.I(\reg_file.reg_storage[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__S0 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__S1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__I1 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__S0 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__S1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__B1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__B2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__B (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__I0 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__I1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__C (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__I0 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__S (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__S (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A2 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__B (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(\reg_file.reg_storage[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__B (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__I1 (.I(\reg_file.reg_storage[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__I2 (.I(\reg_file.reg_storage[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__S0 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__I0 (.I(\reg_file.reg_storage[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__I3 (.I(\reg_file.reg_storage[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__S0 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__S1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__S0 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__S1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__B1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__B (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__B (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__I (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__S (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__C (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__S (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I0 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I1 (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I0 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__S0 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__S1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__B (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__S0 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__S1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__S0 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__S1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__S0 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__S1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__B1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__I (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__B (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__I (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__I0 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__S (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__S (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__B1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__S (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__B (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__I (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__I (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__S0 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__S1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(\reg_file.reg_storage[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__B (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__S0 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__S1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__S0 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__S1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__S0 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__S1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__B (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__B2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__B (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__I0 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__I1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__I0 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__I1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A3 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__B (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__I0 (.I(\reg_file.reg_storage[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__I1 (.I(\reg_file.reg_storage[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__S0 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__S1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__B (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__I0 (.I(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__I1 (.I(\reg_file.reg_storage[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__I2 (.I(\reg_file.reg_storage[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__I3 (.I(\reg_file.reg_storage[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__S0 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__S1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__I0 (.I(\reg_file.reg_storage[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__I3 (.I(\reg_file.reg_storage[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__S0 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__S1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__S0 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__S1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__B1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__B2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__B (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__I0 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__I1 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I0 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__S (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__I (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__B (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__S0 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__S1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__I (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__I (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__I (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__B (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I2 (.I(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S0 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__I0 (.I(\reg_file.reg_storage[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__I3 (.I(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__S0 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__S1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__I (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__I1 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__S0 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__S1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__B1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__B2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__B (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__B (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I0 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I0 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__S (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__B (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__B2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I0 (.I(\reg_file.reg_storage[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I1 (.I(\reg_file.reg_storage[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__S0 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__S1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__B (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I2 (.I(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__S0 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__S1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__I0 (.I(\reg_file.reg_storage[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__I3 (.I(\reg_file.reg_storage[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__S0 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__S1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__I2 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__I3 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__S0 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__S1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__B1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__B (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__B (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__B (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__S0 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__S1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__B (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__S0 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__S1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__S0 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__S1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__S0 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__S1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__B1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__B2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__B (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__S (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I1 (.I(\reg_file.reg_storage[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__S0 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__S1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__B (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__S0 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__S1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__S0 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__S1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__I1 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__S0 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__S1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__B1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__B2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__S (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A2 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__B (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__I (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__B2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__B (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__I (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__S0 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__S1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__B (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I0 (.I(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I2 (.I(\reg_file.reg_storage[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I3 (.I(\reg_file.reg_storage[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__S0 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__S1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__I0 (.I(\reg_file.reg_storage[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__I3 (.I(\reg_file.reg_storage[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__S0 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__S1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__S0 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__S1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__B1 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__B2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__I (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__B (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__B (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A1 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__C (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__B (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__B1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__C1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__C2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__S0 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__S1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__B (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__S0 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__S1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__I0 (.I(\reg_file.reg_storage[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__S0 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__S1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__S0 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__S1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__B (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__C (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__B (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__B1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__C2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__I (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__S0 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__S1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A2 (.I(\reg_file.reg_storage[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__B (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__S0 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__S1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__S0 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__S1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__S0 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__S1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__B1 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__B2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__I (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__S0 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__S1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__B (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__S0 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__S1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__S0 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__S1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__S0 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__S1 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__B1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__B2 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A2 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__C (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__B (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__I (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__B (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__I (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__B (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__B (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__B (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__C (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A4 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__I (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__S (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__S (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__I0 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__S (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__C (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__I1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A1 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__B1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__B (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__B (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__I (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__S (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__S (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A1 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__S (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__C (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__B (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__B (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__S (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__C (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__B (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__B1 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A1 (.I(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__I (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__B2 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__B (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__S (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A2 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A2 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__C (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A2 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__B (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__B1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__B (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A2 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__C (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A3 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__C (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__B (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__C (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__B (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__C (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A2 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__B (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__B1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__B (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__B (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__I0 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__I1 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__S (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__C (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A3 (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__B (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A2 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__B (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A2 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A4 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__B (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__B (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__C (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__B1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__B2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__B2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__B (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__B (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__I0 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__I1 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__S (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A2 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__C (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__I (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A2 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__B (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__B1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__B1 (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A2 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__I (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A3 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__A1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__I (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__I (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A2 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A2 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__B1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A3 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A2 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__B1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__I (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__I (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__B1 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A1 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__A2 (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__B1 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__B (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__I (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__B1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__I (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A2 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__B1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__B2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__B (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A2 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__I (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__I (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__B (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__I (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__B2 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__B (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__I (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A2 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A2 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A2 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__I (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__I (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__B2 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__I (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__B (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A3 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__I (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__S (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__B2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__I (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__S (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__I (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__I (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__I (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__I (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__I (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__B (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__B1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__I (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__I (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__I (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__I (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A2 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__C (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A3 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__B2 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A1 (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__I (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__I (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__S (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A2 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__B1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__I (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__I (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__I (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__B1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__B1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__I (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__B1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__I (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__B1 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A1 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__I (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__I (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__B1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__I (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__B1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__I (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__I (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__I0 (.I(\reg_file.reg_storage[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__S (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__I (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__I (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__B1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__I (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B1 (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__I (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__I (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A1 (.I(\reg_file.reg_storage[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__B1 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A2 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(\reg_file.reg_storage[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__B1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__S (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__I (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__B1 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__I (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__I (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__B1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A1 (.I(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__I (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(\reg_file.reg_storage[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__B1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A1 (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__I (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__I (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__A1 (.I(\reg_file.reg_storage[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__B1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__I (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__I0 (.I(\reg_file.reg_storage[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__S (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__A2 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__B1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__S (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__B1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__S (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A2 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__B1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(\reg_file.reg_storage[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__I (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__B1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A1 (.I(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__I (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__I (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__I (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__B1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__I (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A1 (.I(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__B1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__A1 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__I (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__I (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__B1 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__I (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__B1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__I (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__A1 (.I(\reg_file.reg_storage[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A1 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__B1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__I (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__I (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__B1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__B2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A1 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__I (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__S (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__S (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__I (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__I (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A2 (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__S (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__A2 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A2 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__I (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A2 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A1 (.I(\reg_file.reg_storage[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A2 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__I (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A2 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A2 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__I (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A2 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__I (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__I0 (.I(\reg_file.reg_storage[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__A2 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__A2 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__A1 (.I(\reg_file.reg_storage[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A2 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(\reg_file.reg_storage[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A2 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__I (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(\reg_file.reg_storage[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__I0 (.I(\reg_file.reg_storage[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(\reg_file.reg_storage[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__I (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A2 (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__I (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__I (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__I (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__I (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__I (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__I (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A2 (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A2 (.I(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__A2 (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A2 (.I(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A2 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A2 (.I(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A2 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__A2 (.I(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__I (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A2 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A1 (.I(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A2 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A2 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A2 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__A2 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A2 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__I (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A2 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__I0 (.I(\reg_file.reg_storage[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__S (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A2 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__A2 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(\reg_file.reg_storage[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A2 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A1 (.I(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A2 (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__S (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__I (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A1 (.I(\reg_file.reg_storage[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(\reg_file.reg_storage[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A1 (.I(\reg_file.reg_storage[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__I0 (.I(\reg_file.reg_storage[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__S (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__S (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__S (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A1 (.I(\reg_file.reg_storage[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__I (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A1 (.I(\reg_file.reg_storage[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A1 (.I(\reg_file.reg_storage[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__I (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A1 (.I(\reg_file.reg_storage[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A2 (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__I0 (.I(\reg_file.reg_storage[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__S (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__S (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A2 (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__I (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__I (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__S (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__S (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__I (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__I (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__I (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A2 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A2 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__S (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__I (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A2 (.I(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A2 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A2 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__I (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A2 (.I(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A2 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(\reg_file.reg_storage[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A2 (.I(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A2 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__I (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A2 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A2 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__I (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__I (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I0 (.I(\reg_file.reg_storage[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(\reg_file.reg_storage[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(\reg_file.reg_storage[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__I (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(\reg_file.reg_storage[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__A1 (.I(\reg_file.reg_storage[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__I0 (.I(\reg_file.reg_storage[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(\reg_file.reg_storage[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__I (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A1 (.I(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A2 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(\reg_file.reg_storage[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A2 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__I (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A2 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A2 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(\reg_file.reg_storage[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A2 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A2 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__I (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__I (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__I (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__I (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A1 (.I(\reg_file.reg_storage[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A1 (.I(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__I (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__I1 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(\reg_file.reg_storage[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__I (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__A1 (.I(\reg_file.reg_storage[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A2 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__I (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(\reg_file.reg_storage[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A2 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__I (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A1 (.I(\reg_file.reg_storage[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A2 (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__I (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A2 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__I (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A2 (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__I (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__I (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(\reg_file.reg_storage[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__I (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__I (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__I (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A1 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__I1 (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__I (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A1 (.I(\reg_file.reg_storage[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A1 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A2 (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__I (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A1 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A2 (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__I (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__I (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__I (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A2 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A1 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A2 (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__I1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__S (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__S (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A2 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A1 (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A2 (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__I (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__I (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A2 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A2 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__I (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__I (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A1 (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A2 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__I (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__I (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A2 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__I (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__I (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A1 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A2 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__I (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__I (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__I (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__S (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__I (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__I1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__S (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__I (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A2 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__I (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__S (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__S (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__I (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__I (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A1 (.I(\reg_file.reg_storage[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A1 (.I(\reg_file.reg_storage[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__I1 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__S (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__I (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(\reg_file.reg_storage[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A1 (.I(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(\reg_file.reg_storage[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__I (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(\reg_file.reg_storage[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__I (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__S (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A1 (.I(\reg_file.reg_storage[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__I (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A1 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__I1 (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__S (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A1 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__I (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A1 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__I1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__S (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__S (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__S (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A1 (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A1 (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__I (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A2 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__S (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__I1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__S (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__S (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__S (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__I (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A1 (.I(\reg_file.reg_storage[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__I1 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__S (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A1 (.I(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__I (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__I (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__S (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A1 (.I(\reg_file.reg_storage[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__I1 (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__S (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__I (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A1 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A1 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A1 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__I1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__S (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__S (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A1 (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__I (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A1 (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A1 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__I1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A2 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__I (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__S (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__S (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__I (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A1 (.I(\reg_file.reg_storage[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A1 (.I(\reg_file.reg_storage[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__I1 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__S (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__I (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A1 (.I(\reg_file.reg_storage[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A1 (.I(\reg_file.reg_storage[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__I (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__I (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__I (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__I (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__S (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A1 (.I(\reg_file.reg_storage[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A1 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__I1 (.I(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__S (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__I (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A1 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A1 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A1 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__I1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__S (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__S (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A1 (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__I (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__A1 (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A1 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__I1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__I (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__S (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__I (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__I0 (.I(\reg_file.reg_storage[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__S (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__I (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__I (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__I (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__I (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__I (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__S (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__I (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__I (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__I (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A2 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__I (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__A2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A2 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__I (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__I (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A2 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__A2 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__I (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A2 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A2 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__I (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__I (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A2 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__I (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__I (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__I0 (.I(\reg_file.reg_storage[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__S (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__A2 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__I (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__I (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__I (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__S (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__I (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__I (.I(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__I (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__I (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__I (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__S (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__S (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__S (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A1 (.I(\reg_file.reg_storage[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A2 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__I (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__A2 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__I (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A2 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__I (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__I (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__I (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__I (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A1 (.I(\reg_file.reg_storage[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__I (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__S (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__I (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__S (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__I (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__S (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__S (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__I (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__I (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__I (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__I (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__I0 (.I(\reg_file.reg_storage[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__S (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A2 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A2 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__I (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A2 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A2 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__I0 (.I(\reg_file.reg_storage[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A1 (.I(\reg_file.reg_storage[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__I (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A1 (.I(\reg_file.reg_storage[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__S (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__S (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(\reg_file.reg_storage[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A1 (.I(\reg_file.reg_storage[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__I (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__S (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__S (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__I (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__S (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__I0 (.I(\reg_file.reg_storage[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__S (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__I (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__I (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__I0 (.I(\reg_file.reg_storage[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__S (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__I (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__I (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__I (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__I (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__I (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__S (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A2 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__I0 (.I(\reg_file.reg_storage[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__S (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__I (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(\reg_file.reg_storage[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A2 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A2 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__S (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__S (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__S (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A1 (.I(\reg_file.reg_storage[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__I (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(\reg_file.reg_storage[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(\reg_file.reg_storage[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__S (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8454__S (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__I (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__I (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__S (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__S (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__I (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__I (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__I (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__I (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__S (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__I (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__I (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__I (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__I (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__I (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__I0 (.I(\reg_file.reg_storage[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__S (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__S (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__I (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(\reg_file.reg_storage[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__S (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__S (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__S (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__A2 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A2 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__A2 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A2 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A1 (.I(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__S (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__S (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__I (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__I (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__S (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__S (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__I (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__I (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__I (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__I (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__I (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A1 (.I(\reg_file.reg_storage[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__I1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__S (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__I (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A1 (.I(\reg_file.reg_storage[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A1 (.I(\reg_file.reg_storage[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__I (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__I (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__I (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__I (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__I1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__S (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__I (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A1 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__S (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__I (.I(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__I (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__I1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__S (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__S (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__S (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__I (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A1 (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__I (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__A2 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__A2 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A1 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A2 (.I(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__A2 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A1 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__I1 (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__S (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__S (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A2 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A1 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__S (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__S (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__I (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__I (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__I (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__I (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__A1 (.I(\reg_file.reg_storage[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A1 (.I(\reg_file.reg_storage[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__I1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__S (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A1 (.I(\reg_file.reg_storage[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A1 (.I(\reg_file.reg_storage[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__I (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A1 (.I(\reg_file.reg_storage[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A2 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__A2 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__A2 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__I (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__A2 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__I0 (.I(\reg_file.reg_storage[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__I1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__S (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A1 (.I(\reg_file.reg_storage[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A2 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__I (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A1 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__I0 (.I(\reg_file.reg_storage[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__S (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__I (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__I (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__I0 (.I(\reg_file.reg_storage[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__I1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__S (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__S (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__I0 (.I(\reg_file.reg_storage[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__S (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__I (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__A1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__A2 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A1 (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A2 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__I (.I(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A2 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A1 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A2 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A1 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__I1 (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__S (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__I0 (.I(\reg_file.reg_storage[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__S (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A1 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__I (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__I (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__S (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__S (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__I (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__I (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__I (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__A2 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A2 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__I1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__S (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__I (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__A1 (.I(\reg_file.reg_storage[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__A1 (.I(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__I (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A2 (.I(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__A1 (.I(\reg_file.reg_storage[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A2 (.I(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__I (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A1 (.I(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__A2 (.I(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A1 (.I(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__A2 (.I(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__I (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__I (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__I1 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__S (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A1 (.I(\reg_file.reg_storage[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A1 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__S (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__I (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A2 (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A2 (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__A2 (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__I1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__S (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8762__S (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A2 (.I(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__I (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A2 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__A1 (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__A2 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__A2 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__A2 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A2 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A1 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A2 (.I(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A2 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A1 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A2 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__I1 (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A2 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A1 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A2 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9140__CLK (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(inst[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(inst[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(inst[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(inst[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(inst[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(inst[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(inst[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(inst[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(inst[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(inst[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(inst[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(inst[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(inst[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(inst[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(inst[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(inst[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(inst[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(inst[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(inst[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(inst[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(inst[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(inst[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(inst[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(inst[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(inst[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(mem_load_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(mem_load_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(mem_load_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(mem_load_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(mem_load_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(mem_load_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(mem_load_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(inst[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(mem_load_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(mem_load_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(mem_load_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(mem_load_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(mem_load_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(mem_load_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(mem_load_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(mem_load_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(mem_load_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(mem_load_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(inst[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(mem_load_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(mem_load_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(mem_load_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(mem_load_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(mem_load_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(mem_load_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(mem_load_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(mem_load_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(mem_load_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(mem_load_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(inst[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(mem_load_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(mem_load_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(mem_load_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(mem_load_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(mem_load_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(pc[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(pc[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(pc[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(pc[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(pc[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(inst[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(pc[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(pc[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(pc[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(pc[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(pc[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(pc[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(pc[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(pc[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(pc[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(pc[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(inst[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(pc[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(pc[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(pc[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(pc[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(pc[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(pc[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(pc[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(pc[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(pc[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(pc[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(inst[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(pc[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(pc[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(pc[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(pc[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(pc[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(pc[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(pc[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(inst[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap161_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap162_I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap163_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap164_I (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap165_I (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap166_I (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer11_I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer15_I (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer18_I (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer19_I (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer22_I (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer26_I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer2_I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer34_I (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer37_I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer39_I (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer40_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer4_I (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer52_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer55_I (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer58_I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer59_I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer62_I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4361_ (.I(net27),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4362_ (.A1(net29),
    .A2(_0480_),
    .A3(net28),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4363_ (.I(net23),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4364_ (.I(net29),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4365_ (.A1(_0482_),
    .A2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4366_ (.I(net26),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4367_ (.I(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4368_ (.I(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4369_ (.A1(_0481_),
    .A2(_0484_),
    .B(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4370_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4371_ (.I(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4372_ (.I(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4373_ (.I(net8),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4374_ (.I(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4375_ (.I(net7),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4376_ (.I(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4377_ (.I(net11),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4378_ (.A1(net10),
    .A2(net9),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4379_ (.A1(_0493_),
    .A2(_0495_),
    .A3(_0496_),
    .A4(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4380_ (.A1(_0488_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4381_ (.I(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4382_ (.I(_0500_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4383_ (.I(_0494_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4384_ (.I(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4385_ (.I(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4386_ (.I(_0492_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4387_ (.I(_0505_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4388_ (.I(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4389_ (.I0(\reg_file.reg_storage[4][14] ),
    .I1(\reg_file.reg_storage[5][14] ),
    .I2(\reg_file.reg_storage[6][14] ),
    .I3(\reg_file.reg_storage[7][14] ),
    .S0(_0504_),
    .S1(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4390_ (.I(_0493_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4391_ (.I(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4392_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4393_ (.I(\reg_file.reg_storage[1][14] ),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4394_ (.I(_0494_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4395_ (.I(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4396_ (.I(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4397_ (.A1(_0515_),
    .A2(\reg_file.reg_storage[3][14] ),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4398_ (.I(_0495_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4399_ (.I(_0517_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4400_ (.I(_0493_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4401_ (.I(_0519_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4402_ (.A1(_0518_),
    .A2(\reg_file.reg_storage[2][14] ),
    .B(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4403_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0516_),
    .B2(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4404_ (.I(net7),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4405_ (.I(_0523_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4406_ (.I(_0524_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4407_ (.I(_0506_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4408_ (.I0(\reg_file.reg_storage[12][14] ),
    .I1(\reg_file.reg_storage[13][14] ),
    .I2(\reg_file.reg_storage[14][14] ),
    .I3(\reg_file.reg_storage[15][14] ),
    .S0(_0525_),
    .S1(_0526_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4409_ (.I0(\reg_file.reg_storage[8][14] ),
    .I1(\reg_file.reg_storage[9][14] ),
    .I2(\reg_file.reg_storage[10][14] ),
    .I3(\reg_file.reg_storage[11][14] ),
    .S0(_0525_),
    .S1(_0507_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4410_ (.I(net9),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4412_ (.I(_0530_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4413_ (.I(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4414_ (.I(net10),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4415_ (.I(_0533_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4416_ (.I(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4417_ (.I0(_0508_),
    .I1(_0522_),
    .I2(_0527_),
    .I3(_0528_),
    .S0(_0532_),
    .S1(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4418_ (.A1(net70),
    .A2(_0491_),
    .B1(_0501_),
    .B2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4419_ (.A1(net29),
    .A2(net28),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4420_ (.A1(net26),
    .A2(net23),
    .A3(net27),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4421_ (.A1(_0538_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4422_ (.A1(net27),
    .A2(_0538_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4423_ (.A1(_0481_),
    .A2(_0541_),
    .B(_0486_),
    .C(_0482_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4424_ (.A1(_0485_),
    .A2(net23),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4425_ (.A1(net28),
    .A2(_0539_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4426_ (.I(net29),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4427_ (.A1(_0543_),
    .A2(_0541_),
    .B1(_0544_),
    .B2(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4428_ (.A1(_0540_),
    .A2(_0542_),
    .A3(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4429_ (.I(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4430_ (.I(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4431_ (.I(net6),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4432_ (.I(_0483_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4433_ (.I(net27),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4434_ (.A1(_0482_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4435_ (.I(_0485_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4436_ (.A1(_0554_),
    .A2(_0483_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4437_ (.A1(_0551_),
    .A2(_0553_),
    .B1(_0555_),
    .B2(_0552_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4438_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4439_ (.I(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4440_ (.A1(net25),
    .A2(_0556_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4441_ (.I(_0559_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4442_ (.A1(_0550_),
    .A2(_0558_),
    .B(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4443_ (.I(net16),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4444_ (.I(net15),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4445_ (.I(net14),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4446_ (.I(net13),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4447_ (.I(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4448_ (.A1(_0564_),
    .A2(_0566_),
    .A3(net17),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4449_ (.A1(_0562_),
    .A2(_0563_),
    .A3(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4450_ (.A1(_0540_),
    .A2(_0542_),
    .A3(_0546_),
    .A4(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4451_ (.I(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4452_ (.I(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4453_ (.I(net13),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4454_ (.I(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4455_ (.I(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4456_ (.I(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4457_ (.I(net14),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4458_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4459_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4460_ (.I(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4461_ (.I0(\reg_file.reg_storage[4][14] ),
    .I1(\reg_file.reg_storage[5][14] ),
    .I2(\reg_file.reg_storage[6][14] ),
    .I3(\reg_file.reg_storage[7][14] ),
    .S0(_0575_),
    .S1(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4462_ (.I(_0564_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4463_ (.I(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4464_ (.I(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4465_ (.I(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4466_ (.I(_0565_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4467_ (.I(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4468_ (.I(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4469_ (.A1(_0587_),
    .A2(\reg_file.reg_storage[3][14] ),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4470_ (.I(_0566_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4471_ (.I(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4472_ (.I(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4473_ (.I(_0581_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4474_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4475_ (.A1(_0591_),
    .A2(\reg_file.reg_storage[2][14] ),
    .B(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4476_ (.A1(_0584_),
    .A2(_0512_),
    .B1(_0588_),
    .B2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4477_ (.I(_0574_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4478_ (.I(_0578_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4479_ (.I0(\reg_file.reg_storage[12][14] ),
    .I1(\reg_file.reg_storage[13][14] ),
    .I2(\reg_file.reg_storage[14][14] ),
    .I3(\reg_file.reg_storage[15][14] ),
    .S0(_0596_),
    .S1(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4480_ (.I0(\reg_file.reg_storage[8][14] ),
    .I1(\reg_file.reg_storage[9][14] ),
    .I2(\reg_file.reg_storage[10][14] ),
    .I3(\reg_file.reg_storage[11][14] ),
    .S0(_0596_),
    .S1(_0597_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4481_ (.I(_0563_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4482_ (.I(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4483_ (.I(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4484_ (.I(net16),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4485_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4486_ (.I0(_0580_),
    .I1(_0595_),
    .I2(_0598_),
    .I3(_0599_),
    .S0(_0602_),
    .S1(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4487_ (.A1(_0549_),
    .A2(_0561_),
    .B1(_0571_),
    .B2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4488_ (.A1(_0537_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4489_ (.A1(_0537_),
    .A2(_0606_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4490_ (.A1(_0607_),
    .A2(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4491_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4492_ (.I(_0489_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4493_ (.I(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4494_ (.I(_0499_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4495_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4496_ (.I(net9),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4497_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4498_ (.I0(\reg_file.reg_storage[2][13] ),
    .I1(\reg_file.reg_storage[3][13] ),
    .S(_0513_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4499_ (.I(net8),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4500_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4501_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4502_ (.I0(\reg_file.reg_storage[1][13] ),
    .I1(_0617_),
    .S(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4503_ (.I(_0530_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4504_ (.I(net7),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4505_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4506_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(\reg_file.reg_storage[5][13] ),
    .I2(\reg_file.reg_storage[6][13] ),
    .I3(\reg_file.reg_storage[7][13] ),
    .S0(_0624_),
    .S1(_0619_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4507_ (.A1(_0622_),
    .A2(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4508_ (.I(_0533_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4509_ (.A1(_0616_),
    .A2(_0621_),
    .B(_0626_),
    .C(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4510_ (.I(_0622_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4511_ (.I(_0623_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4512_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4513_ (.I(_0505_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4514_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(\reg_file.reg_storage[13][13] ),
    .I2(\reg_file.reg_storage[14][13] ),
    .I3(\reg_file.reg_storage[15][13] ),
    .S0(_0631_),
    .S1(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4515_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(\reg_file.reg_storage[9][13] ),
    .I2(\reg_file.reg_storage[10][13] ),
    .I3(\reg_file.reg_storage[11][13] ),
    .S0(_0624_),
    .S1(_0619_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4516_ (.A1(_0615_),
    .A2(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4517_ (.I(_0534_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4518_ (.A1(_0629_),
    .A2(_0633_),
    .B(_0635_),
    .C(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4519_ (.A1(_0628_),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4520_ (.A1(net69),
    .A2(_0612_),
    .B1(_0614_),
    .B2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4521_ (.I(_0547_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4522_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4523_ (.I(net5),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4524_ (.A1(_0642_),
    .A2(_0558_),
    .B(_0560_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4525_ (.I(_0565_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4526_ (.I(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4527_ (.I(_0564_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4528_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4529_ (.I0(\reg_file.reg_storage[4][13] ),
    .I1(\reg_file.reg_storage[5][13] ),
    .I2(\reg_file.reg_storage[6][13] ),
    .I3(\reg_file.reg_storage[7][13] ),
    .S0(_0645_),
    .S1(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4530_ (.I(_0592_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4531_ (.I(\reg_file.reg_storage[1][13] ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4532_ (.I(_0585_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4533_ (.I(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4534_ (.A1(_0652_),
    .A2(\reg_file.reg_storage[3][13] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4535_ (.I(_0589_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4536_ (.I(_0582_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4537_ (.A1(_0654_),
    .A2(\reg_file.reg_storage[2][13] ),
    .B(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4538_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_0653_),
    .B2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4539_ (.I(_0644_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4540_ (.I0(\reg_file.reg_storage[12][13] ),
    .I1(\reg_file.reg_storage[13][13] ),
    .I2(\reg_file.reg_storage[14][13] ),
    .I3(\reg_file.reg_storage[15][13] ),
    .S0(_0658_),
    .S1(_0647_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4541_ (.I0(\reg_file.reg_storage[8][13] ),
    .I1(\reg_file.reg_storage[9][13] ),
    .I2(\reg_file.reg_storage[10][13] ),
    .I3(\reg_file.reg_storage[11][13] ),
    .S0(_0645_),
    .S1(_0647_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4542_ (.I(_0563_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4543_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4544_ (.I(net16),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4545_ (.I(_0663_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4546_ (.I0(_0648_),
    .I1(_0657_),
    .I2(_0659_),
    .I3(_0660_),
    .S0(_0662_),
    .S1(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4547_ (.I(_0569_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4548_ (.I(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4549_ (.A1(_0641_),
    .A2(_0643_),
    .B1(_0665_),
    .B2(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4550_ (.A1(_0639_),
    .A2(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4551_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4552_ (.I(net68),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4553_ (.I(_0489_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4554_ (.I(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4555_ (.I(_0500_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4556_ (.I(_0615_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4557_ (.I(_0513_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4558_ (.I0(\reg_file.reg_storage[2][12] ),
    .I1(\reg_file.reg_storage[3][12] ),
    .S(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4559_ (.I(_0492_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4560_ (.I(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4561_ (.I0(\reg_file.reg_storage[1][12] ),
    .I1(_0677_),
    .S(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4562_ (.I(_0530_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4563_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4564_ (.I(_0630_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4565_ (.I(_0492_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4566_ (.I(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4567_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(\reg_file.reg_storage[5][12] ),
    .I2(\reg_file.reg_storage[6][12] ),
    .I3(\reg_file.reg_storage[7][12] ),
    .S0(_0683_),
    .S1(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4568_ (.A1(_0682_),
    .A2(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4569_ (.I(_0627_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4570_ (.A1(_0675_),
    .A2(_0680_),
    .B(_0687_),
    .C(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _4571_ (.I(_0682_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4572_ (.I(_0683_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4573_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(\reg_file.reg_storage[13][12] ),
    .I2(\reg_file.reg_storage[14][12] ),
    .I3(\reg_file.reg_storage[15][12] ),
    .S0(_0691_),
    .S1(_0679_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4574_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(\reg_file.reg_storage[9][12] ),
    .I2(\reg_file.reg_storage[10][12] ),
    .I3(\reg_file.reg_storage[11][12] ),
    .S0(_0631_),
    .S1(_0685_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4575_ (.A1(_0616_),
    .A2(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4576_ (.I(_0533_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4577_ (.I(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4578_ (.A1(_0690_),
    .A2(_0692_),
    .B(_0694_),
    .C(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4579_ (.A1(_0689_),
    .A2(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4580_ (.A1(_0671_),
    .A2(_0673_),
    .B1(_0674_),
    .B2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4581_ (.I(net4),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4582_ (.A1(_0700_),
    .A2(_0558_),
    .B(_0560_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4583_ (.I(_0573_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4584_ (.I(_0577_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4585_ (.I(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4586_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(\reg_file.reg_storage[5][12] ),
    .I2(\reg_file.reg_storage[6][12] ),
    .I3(\reg_file.reg_storage[7][12] ),
    .S0(_0702_),
    .S1(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4587_ (.I(_0655_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4588_ (.I(\reg_file.reg_storage[1][12] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4589_ (.I(_0572_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4590_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4591_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4592_ (.I(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4593_ (.A1(_0711_),
    .A2(\reg_file.reg_storage[3][12] ),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4594_ (.A1(_0591_),
    .A2(\reg_file.reg_storage[2][12] ),
    .B(_0649_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4595_ (.A1(_0706_),
    .A2(_0707_),
    .B1(_0712_),
    .B2(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4596_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(\reg_file.reg_storage[13][12] ),
    .I2(\reg_file.reg_storage[14][12] ),
    .I3(\reg_file.reg_storage[15][12] ),
    .S0(_0710_),
    .S1(_0704_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4597_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(\reg_file.reg_storage[9][12] ),
    .I2(\reg_file.reg_storage[10][12] ),
    .I3(\reg_file.reg_storage[11][12] ),
    .S0(_0710_),
    .S1(_0704_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4598_ (.I(_0601_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4599_ (.I(_0603_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4600_ (.I0(_0705_),
    .I1(_0714_),
    .I2(_0715_),
    .I3(_0716_),
    .S0(_0717_),
    .S1(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4601_ (.A1(_0549_),
    .A2(_0701_),
    .B1(_0719_),
    .B2(_0571_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4602_ (.A1(_0699_),
    .A2(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4603_ (.A1(_0699_),
    .A2(_0720_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4604_ (.A1(_0722_),
    .A2(_0721_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4605_ (.I(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4606_ (.I(_0490_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4607_ (.I(_0613_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4608_ (.I(_0523_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4609_ (.I(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4610_ (.I(_0618_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4611_ (.I(_0729_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4612_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(\reg_file.reg_storage[5][11] ),
    .I2(\reg_file.reg_storage[6][11] ),
    .I3(\reg_file.reg_storage[7][11] ),
    .S0(_0728_),
    .S1(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4613_ (.I(_0493_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4614_ (.I(_0732_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4615_ (.I(\reg_file.reg_storage[1][11] ),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4616_ (.I(_0513_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4617_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_0736_),
    .A2(\reg_file.reg_storage[3][11] ),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4619_ (.A1(_0518_),
    .A2(\reg_file.reg_storage[2][11] ),
    .B(_0520_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4620_ (.A1(_0733_),
    .A2(_0734_),
    .B1(_0737_),
    .B2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4621_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(\reg_file.reg_storage[13][11] ),
    .I2(\reg_file.reg_storage[14][11] ),
    .I3(\reg_file.reg_storage[15][11] ),
    .S0(_0514_),
    .S1(_0730_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4622_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(\reg_file.reg_storage[9][11] ),
    .I2(\reg_file.reg_storage[10][11] ),
    .I3(\reg_file.reg_storage[11][11] ),
    .S0(_0728_),
    .S1(_0730_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4623_ (.I(_0681_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4624_ (.I0(_0731_),
    .I1(_0739_),
    .I2(_0740_),
    .I3(_0741_),
    .S0(_0742_),
    .S1(_0535_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4625_ (.A1(net67),
    .A2(_0725_),
    .B1(_0726_),
    .B2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4626_ (.I(_0640_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4627_ (.I(net25),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4628_ (.I(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4629_ (.A1(_0485_),
    .A2(net23),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4630_ (.A1(_0545_),
    .A2(_0552_),
    .A3(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4631_ (.I(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4632_ (.A1(_0747_),
    .A2(_0557_),
    .A3(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4633_ (.I(_0750_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4634_ (.A1(net30),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4635_ (.I(_0566_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4636_ (.I(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4637_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4638_ (.I(_0545_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4639_ (.I(_0552_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4640_ (.A1(_0757_),
    .A2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4641_ (.A1(_0554_),
    .A2(_0756_),
    .A3(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4642_ (.A1(_0751_),
    .A2(_0753_),
    .A3(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4643_ (.I(_0651_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4644_ (.I(_0564_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4645_ (.I(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4646_ (.I0(\reg_file.reg_storage[4][11] ),
    .I1(\reg_file.reg_storage[5][11] ),
    .I2(\reg_file.reg_storage[6][11] ),
    .I3(\reg_file.reg_storage[7][11] ),
    .S0(net185),
    .S1(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4647_ (.I(_0583_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4648_ (.I(_0586_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4649_ (.A1(_0767_),
    .A2(\reg_file.reg_storage[3][11] ),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4650_ (.I(_0590_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4651_ (.I(_0592_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4652_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][11] ),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4653_ (.A1(_0766_),
    .A2(_0734_),
    .B1(_0768_),
    .B2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4654_ (.I0(\reg_file.reg_storage[12][11] ),
    .I1(\reg_file.reg_storage[13][11] ),
    .I2(\reg_file.reg_storage[14][11] ),
    .I3(\reg_file.reg_storage[15][11] ),
    .S0(_0586_),
    .S1(_0764_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4655_ (.I0(\reg_file.reg_storage[8][11] ),
    .I1(\reg_file.reg_storage[9][11] ),
    .I2(\reg_file.reg_storage[10][11] ),
    .I3(\reg_file.reg_storage[11][11] ),
    .S0(net185),
    .S1(_0764_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4656_ (.I(_0663_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4657_ (.I0(_0765_),
    .I1(_0772_),
    .I2(_0773_),
    .I3(_0774_),
    .S0(_0602_),
    .S1(_0775_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4658_ (.I(_0570_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4659_ (.A1(_0745_),
    .A2(_0761_),
    .B1(_0776_),
    .B2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4660_ (.A1(_0744_),
    .A2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4661_ (.A1(_0744_),
    .A2(_0778_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4662_ (.A1(_0779_),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4663_ (.I(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4664_ (.I(_0500_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4665_ (.I(_0523_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4666_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4667_ (.I(net8),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4668_ (.I(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4669_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(\reg_file.reg_storage[5][10] ),
    .I2(\reg_file.reg_storage[6][10] ),
    .I3(\reg_file.reg_storage[7][10] ),
    .S0(_0785_),
    .S1(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4670_ (.I(_0510_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4671_ (.I(\reg_file.reg_storage[1][10] ),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4672_ (.I(_0624_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4673_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_0792_),
    .A2(\reg_file.reg_storage[3][10] ),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4675_ (.I(_0517_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4676_ (.I(_0519_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4677_ (.A1(_0794_),
    .A2(\reg_file.reg_storage[2][10] ),
    .B(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4678_ (.A1(_0789_),
    .A2(_0790_),
    .B1(_0793_),
    .B2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4679_ (.I(_0784_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4680_ (.I(_0505_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4681_ (.I(_0799_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4682_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(\reg_file.reg_storage[13][10] ),
    .I2(\reg_file.reg_storage[14][10] ),
    .I3(\reg_file.reg_storage[15][10] ),
    .S0(_0798_),
    .S1(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4683_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(\reg_file.reg_storage[9][10] ),
    .I2(\reg_file.reg_storage[10][10] ),
    .I3(\reg_file.reg_storage[11][10] ),
    .S0(_0798_),
    .S1(_0800_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4684_ (.I(_0622_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4685_ (.I(_0533_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4686_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4687_ (.I0(_0788_),
    .I1(_0797_),
    .I2(_0801_),
    .I3(_0802_),
    .S0(_0803_),
    .S1(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4688_ (.A1(net66),
    .A2(_0673_),
    .B1(_0783_),
    .B2(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4689_ (.I(_0482_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4690_ (.A1(_0808_),
    .A2(_0757_),
    .A3(_0758_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4691_ (.I(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4692_ (.A1(net24),
    .A2(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4693_ (.I0(\reg_file.reg_storage[4][10] ),
    .I1(\reg_file.reg_storage[5][10] ),
    .I2(\reg_file.reg_storage[6][10] ),
    .I3(\reg_file.reg_storage[7][10] ),
    .S0(_0710_),
    .S1(_0579_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4694_ (.I(_0575_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4695_ (.A1(_0813_),
    .A2(\reg_file.reg_storage[3][10] ),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4696_ (.A1(_0591_),
    .A2(\reg_file.reg_storage[2][10] ),
    .B(_0593_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4697_ (.A1(_0706_),
    .A2(_0790_),
    .B1(_0814_),
    .B2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4698_ (.I0(\reg_file.reg_storage[12][10] ),
    .I1(\reg_file.reg_storage[13][10] ),
    .I2(\reg_file.reg_storage[14][10] ),
    .I3(\reg_file.reg_storage[15][10] ),
    .S0(_0575_),
    .S1(_0579_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4699_ (.I0(\reg_file.reg_storage[8][10] ),
    .I1(\reg_file.reg_storage[9][10] ),
    .I2(\reg_file.reg_storage[10][10] ),
    .I3(\reg_file.reg_storage[11][10] ),
    .S0(_0575_),
    .S1(_0579_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4700_ (.I0(_0812_),
    .I1(_0816_),
    .I2(_0817_),
    .I3(_0818_),
    .S0(_0717_),
    .S1(_0604_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4701_ (.A1(_0549_),
    .A2(_0811_),
    .B1(_0819_),
    .B2(_0571_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4702_ (.A1(_0807_),
    .A2(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4703_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4704_ (.A1(_0807_),
    .A2(_0820_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4705_ (.A1(_0822_),
    .A2(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4706_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4707_ (.I(net96),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4708_ (.I0(\reg_file.reg_storage[2][9] ),
    .I1(\reg_file.reg_storage[3][9] ),
    .S(_0727_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4709_ (.I0(\reg_file.reg_storage[1][9] ),
    .I1(_0827_),
    .S(_0620_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4710_ (.I(_0618_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4711_ (.I0(\reg_file.reg_storage[4][9] ),
    .I1(\reg_file.reg_storage[5][9] ),
    .I2(\reg_file.reg_storage[6][9] ),
    .I3(\reg_file.reg_storage[7][9] ),
    .S0(_0624_),
    .S1(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4712_ (.A1(_0622_),
    .A2(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4713_ (.I(_0627_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4714_ (.A1(_0616_),
    .A2(_0828_),
    .B(_0831_),
    .C(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4715_ (.I0(\reg_file.reg_storage[12][9] ),
    .I1(\reg_file.reg_storage[13][9] ),
    .I2(\reg_file.reg_storage[14][9] ),
    .I3(\reg_file.reg_storage[15][9] ),
    .S0(_0683_),
    .S1(_0620_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4716_ (.I(net9),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4717_ (.I(_0623_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4718_ (.I(_0618_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4719_ (.I0(\reg_file.reg_storage[8][9] ),
    .I1(\reg_file.reg_storage[9][9] ),
    .I2(\reg_file.reg_storage[10][9] ),
    .I3(\reg_file.reg_storage[11][9] ),
    .S0(_0836_),
    .S1(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4720_ (.A1(_0835_),
    .A2(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4721_ (.A1(_0532_),
    .A2(_0834_),
    .B(_0839_),
    .C(_0636_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(_0833_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4723_ (.A1(_0826_),
    .A2(_0725_),
    .B1(_0501_),
    .B2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4724_ (.I(_0640_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4725_ (.I(_0809_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4726_ (.A1(net22),
    .A2(_0844_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4727_ (.I(_0644_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4728_ (.I(_0576_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4729_ (.I(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4730_ (.I0(\reg_file.reg_storage[4][9] ),
    .I1(\reg_file.reg_storage[5][9] ),
    .I2(\reg_file.reg_storage[6][9] ),
    .I3(\reg_file.reg_storage[7][9] ),
    .S0(_0846_),
    .S1(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4731_ (.I(\reg_file.reg_storage[1][9] ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4732_ (.A1(_0702_),
    .A2(\reg_file.reg_storage[3][9] ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4733_ (.I(_0589_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4734_ (.I(_0581_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4735_ (.A1(_0852_),
    .A2(\reg_file.reg_storage[2][9] ),
    .B(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4736_ (.A1(_0593_),
    .A2(_0850_),
    .B1(_0851_),
    .B2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4737_ (.I0(\reg_file.reg_storage[12][9] ),
    .I1(\reg_file.reg_storage[13][9] ),
    .I2(\reg_file.reg_storage[14][9] ),
    .I3(\reg_file.reg_storage[15][9] ),
    .S0(_0709_),
    .S1(_0848_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4738_ (.I0(\reg_file.reg_storage[8][9] ),
    .I1(\reg_file.reg_storage[9][9] ),
    .I2(\reg_file.reg_storage[10][9] ),
    .I3(\reg_file.reg_storage[11][9] ),
    .S0(_0846_),
    .S1(_0848_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4739_ (.I(_0661_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4740_ (.I(_0663_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4741_ (.I0(_0849_),
    .I1(_0855_),
    .I2(_0856_),
    .I3(_0857_),
    .S0(_0858_),
    .S1(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4742_ (.I(_0666_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4743_ (.A1(_0843_),
    .A2(_0845_),
    .B1(_0860_),
    .B2(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4744_ (.A1(_0842_),
    .A2(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4745_ (.I(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4746_ (.I(_0611_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4747_ (.I(_0865_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4748_ (.I0(\reg_file.reg_storage[2][8] ),
    .I1(\reg_file.reg_storage[3][8] ),
    .S(_0798_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4749_ (.I(_0829_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4750_ (.I0(\reg_file.reg_storage[1][8] ),
    .I1(_0867_),
    .S(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4751_ (.I(_0729_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4752_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(\reg_file.reg_storage[5][8] ),
    .I2(\reg_file.reg_storage[6][8] ),
    .I3(\reg_file.reg_storage[7][8] ),
    .S0(_0791_),
    .S1(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4753_ (.A1(_0803_),
    .A2(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4754_ (.A1(_0675_),
    .A2(_0869_),
    .B(_0872_),
    .C(_0688_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4755_ (.I(_0529_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4756_ (.I(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4757_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(\reg_file.reg_storage[13][8] ),
    .I2(\reg_file.reg_storage[14][8] ),
    .I3(\reg_file.reg_storage[15][8] ),
    .S0(_0736_),
    .S1(_0868_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4758_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(\reg_file.reg_storage[9][8] ),
    .I2(\reg_file.reg_storage[10][8] ),
    .I3(\reg_file.reg_storage[11][8] ),
    .S0(_0735_),
    .S1(_0870_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4759_ (.A1(_0675_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4760_ (.A1(_0875_),
    .A2(_0876_),
    .B(_0878_),
    .C(_0696_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4761_ (.A1(_0873_),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4762_ (.A1(net95),
    .A2(_0866_),
    .B1(_0674_),
    .B2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4763_ (.I(_0548_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4764_ (.A1(net21),
    .A2(_0844_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4765_ (.I(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4766_ (.I(_0585_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4767_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4768_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4769_ (.I(_0703_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4770_ (.I0(\reg_file.reg_storage[4][8] ),
    .I1(\reg_file.reg_storage[5][8] ),
    .I2(\reg_file.reg_storage[6][8] ),
    .I3(\reg_file.reg_storage[7][8] ),
    .S0(_0887_),
    .S1(_0888_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4771_ (.I(_0770_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4772_ (.I(\reg_file.reg_storage[1][8] ),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4773_ (.I(_0754_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4774_ (.I(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4775_ (.A1(_0893_),
    .A2(\reg_file.reg_storage[3][8] ),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4776_ (.I(_0590_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4777_ (.A1(_0895_),
    .A2(\reg_file.reg_storage[2][8] ),
    .B(_0766_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4778_ (.A1(_0890_),
    .A2(_0891_),
    .B1(_0894_),
    .B2(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4779_ (.I0(\reg_file.reg_storage[12][8] ),
    .I1(\reg_file.reg_storage[13][8] ),
    .I2(\reg_file.reg_storage[14][8] ),
    .I3(\reg_file.reg_storage[15][8] ),
    .S0(_0755_),
    .S1(_0888_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4780_ (.I0(\reg_file.reg_storage[8][8] ),
    .I1(\reg_file.reg_storage[9][8] ),
    .I2(\reg_file.reg_storage[10][8] ),
    .I3(\reg_file.reg_storage[11][8] ),
    .S0(_0755_),
    .S1(_0888_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4781_ (.I(_0662_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4782_ (.I0(_0889_),
    .I1(_0897_),
    .I2(_0898_),
    .I3(_0899_),
    .S0(_0900_),
    .S1(_0718_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4783_ (.I(_0570_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4784_ (.A1(_0882_),
    .A2(_0884_),
    .B1(_0901_),
    .B2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4785_ (.A1(_0881_),
    .A2(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4786_ (.A1(_0881_),
    .A2(_0903_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4787_ (.A1(_0904_),
    .A2(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4788_ (.I(_0906_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4789_ (.I(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4790_ (.A1(_0483_),
    .A2(_0553_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4791_ (.I(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4792_ (.I(_0749_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4793_ (.A1(net2),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4794_ (.A1(_0562_),
    .A2(_0910_),
    .A3(_0911_),
    .B(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4795_ (.I(_0565_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4796_ (.I(_0576_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4797_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(\reg_file.reg_storage[5][3] ),
    .I2(\reg_file.reg_storage[6][3] ),
    .I3(\reg_file.reg_storage[7][3] ),
    .S0(_0914_),
    .S1(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4798_ (.I(\reg_file.reg_storage[1][3] ),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4799_ (.A1(_0708_),
    .A2(\reg_file.reg_storage[3][3] ),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4800_ (.A1(_0589_),
    .A2(\reg_file.reg_storage[2][3] ),
    .B(_0581_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4801_ (.A1(_0582_),
    .A2(_0917_),
    .B1(_0918_),
    .B2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4802_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(\reg_file.reg_storage[13][3] ),
    .I2(\reg_file.reg_storage[14][3] ),
    .I3(\reg_file.reg_storage[15][3] ),
    .S0(_0566_),
    .S1(_0915_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4803_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(\reg_file.reg_storage[9][3] ),
    .I2(\reg_file.reg_storage[10][3] ),
    .I3(\reg_file.reg_storage[11][3] ),
    .S0(_0914_),
    .S1(_0915_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4804_ (.I0(_0916_),
    .I1(_0920_),
    .I2(_0921_),
    .I3(_0922_),
    .S0(_0600_),
    .S1(_0663_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4805_ (.A1(_0547_),
    .A2(_0913_),
    .B1(_0923_),
    .B2(_0666_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4806_ (.I(_0623_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4807_ (.I0(\reg_file.reg_storage[4][3] ),
    .I1(\reg_file.reg_storage[5][3] ),
    .I2(\reg_file.reg_storage[6][3] ),
    .I3(\reg_file.reg_storage[7][3] ),
    .S0(_0925_),
    .S1(_0837_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4808_ (.A1(_0784_),
    .A2(\reg_file.reg_storage[3][3] ),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4809_ (.I(_0495_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4810_ (.A1(_0928_),
    .A2(\reg_file.reg_storage[2][3] ),
    .B(_0509_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4811_ (.A1(_0732_),
    .A2(_0917_),
    .B1(_0927_),
    .B2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4812_ (.I0(\reg_file.reg_storage[12][3] ),
    .I1(\reg_file.reg_storage[13][3] ),
    .I2(\reg_file.reg_storage[14][3] ),
    .I3(\reg_file.reg_storage[15][3] ),
    .S0(_0836_),
    .S1(_0829_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4813_ (.I0(\reg_file.reg_storage[8][3] ),
    .I1(\reg_file.reg_storage[9][3] ),
    .I2(\reg_file.reg_storage[10][3] ),
    .I3(\reg_file.reg_storage[11][3] ),
    .S0(_0836_),
    .S1(_0829_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4814_ (.I0(_0926_),
    .I1(_0930_),
    .I2(_0931_),
    .I3(_0932_),
    .S0(_0874_),
    .S1(_0534_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4815_ (.A1(net90),
    .A2(_0490_),
    .B1(_0613_),
    .B2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4816_ (.A1(_0934_),
    .A2(_0924_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4817_ (.A1(net32),
    .A2(_0750_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4818_ (.A1(_0661_),
    .A2(_0909_),
    .A3(_0911_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4819_ (.A1(_0936_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4820_ (.I(net15),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4821_ (.I0(\reg_file.reg_storage[2][2] ),
    .I1(\reg_file.reg_storage[3][2] ),
    .S(_0573_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4822_ (.I0(\reg_file.reg_storage[1][2] ),
    .I1(_0940_),
    .S(_0578_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4823_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(\reg_file.reg_storage[5][2] ),
    .I2(\reg_file.reg_storage[6][2] ),
    .I3(\reg_file.reg_storage[7][2] ),
    .S0(_0914_),
    .S1(_0847_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4824_ (.A1(_0661_),
    .A2(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4825_ (.I(_0562_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4826_ (.A1(_0939_),
    .A2(_0941_),
    .B(_0943_),
    .C(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4827_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(\reg_file.reg_storage[13][2] ),
    .I2(\reg_file.reg_storage[14][2] ),
    .I3(\reg_file.reg_storage[15][2] ),
    .S0(_0885_),
    .S1(_0763_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4828_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(\reg_file.reg_storage[9][2] ),
    .I2(\reg_file.reg_storage[10][2] ),
    .I3(\reg_file.reg_storage[11][2] ),
    .S0(_0914_),
    .S1(_0915_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4829_ (.A1(_0939_),
    .A2(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4830_ (.A1(_0601_),
    .A2(_0946_),
    .B(_0948_),
    .C(_0603_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4831_ (.A1(_0945_),
    .A2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4832_ (.A1(_0640_),
    .A2(_0938_),
    .B1(_0950_),
    .B2(_0666_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4833_ (.I0(\reg_file.reg_storage[4][2] ),
    .I1(\reg_file.reg_storage[5][2] ),
    .I2(\reg_file.reg_storage[6][2] ),
    .I3(\reg_file.reg_storage[7][2] ),
    .S0(_0925_),
    .S1(_0506_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4834_ (.I(_0509_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4835_ (.I(\reg_file.reg_storage[1][2] ),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4836_ (.I(_0494_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4837_ (.I(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4838_ (.A1(_0956_),
    .A2(\reg_file.reg_storage[3][2] ),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4839_ (.A1(_0928_),
    .A2(\reg_file.reg_storage[2][2] ),
    .B(_0519_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4840_ (.A1(_0953_),
    .A2(_0954_),
    .B1(_0957_),
    .B2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4841_ (.I0(\reg_file.reg_storage[12][2] ),
    .I1(\reg_file.reg_storage[13][2] ),
    .I2(\reg_file.reg_storage[14][2] ),
    .I3(\reg_file.reg_storage[15][2] ),
    .S0(_0925_),
    .S1(_0837_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4842_ (.I0(\reg_file.reg_storage[8][2] ),
    .I1(\reg_file.reg_storage[9][2] ),
    .I2(\reg_file.reg_storage[10][2] ),
    .I3(\reg_file.reg_storage[11][2] ),
    .S0(_0925_),
    .S1(_0837_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4843_ (.I0(_0952_),
    .I1(_0959_),
    .I2(_0960_),
    .I3(_0961_),
    .S0(_0874_),
    .S1(_0804_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4844_ (.A1(net87),
    .A2(_0490_),
    .B1(_0500_),
    .B2(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4845_ (.A1(_0951_),
    .A2(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4846_ (.A1(net207),
    .A2(net173),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4847_ (.A1(_0551_),
    .A2(_0480_),
    .A3(net31),
    .A4(_0543_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4848_ (.A1(_0853_),
    .A2(_0909_),
    .A3(_0911_),
    .B(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4849_ (.I0(\reg_file.reg_storage[2][1] ),
    .I1(\reg_file.reg_storage[3][1] ),
    .S(_0585_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4850_ (.I(_0576_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4851_ (.I0(\reg_file.reg_storage[1][1] ),
    .I1(_0968_),
    .S(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4852_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(\reg_file.reg_storage[5][1] ),
    .I2(\reg_file.reg_storage[6][1] ),
    .I3(\reg_file.reg_storage[7][1] ),
    .S0(_0572_),
    .S1(_0577_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4853_ (.A1(_0600_),
    .A2(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4854_ (.A1(_0939_),
    .A2(_0970_),
    .B(_0972_),
    .C(_0944_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4855_ (.I(_0600_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4856_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(\reg_file.reg_storage[13][1] ),
    .I2(\reg_file.reg_storage[14][1] ),
    .I3(\reg_file.reg_storage[15][1] ),
    .S0(_0708_),
    .S1(_0969_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4857_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(\reg_file.reg_storage[9][1] ),
    .I2(\reg_file.reg_storage[10][1] ),
    .I3(\reg_file.reg_storage[11][1] ),
    .S0(_0572_),
    .S1(_0577_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4858_ (.A1(_0939_),
    .A2(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4859_ (.A1(_0974_),
    .A2(_0975_),
    .B(_0977_),
    .C(_0603_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4860_ (.A1(_0973_),
    .A2(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4861_ (.A1(_0843_),
    .A2(net209),
    .B1(_0979_),
    .B2(_0861_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4862_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(\reg_file.reg_storage[5][1] ),
    .I2(\reg_file.reg_storage[6][1] ),
    .I3(\reg_file.reg_storage[7][1] ),
    .S0(_0955_),
    .S1(_0729_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4863_ (.I(\reg_file.reg_storage[1][1] ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4864_ (.A1(_0784_),
    .A2(\reg_file.reg_storage[3][1] ),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4865_ (.A1(_0928_),
    .A2(\reg_file.reg_storage[2][1] ),
    .B(_0509_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4866_ (.A1(_0732_),
    .A2(_0982_),
    .B1(_0983_),
    .B2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4867_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(\reg_file.reg_storage[13][1] ),
    .I2(\reg_file.reg_storage[14][1] ),
    .I3(\reg_file.reg_storage[15][1] ),
    .S0(_0955_),
    .S1(_0678_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4868_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(\reg_file.reg_storage[9][1] ),
    .I2(\reg_file.reg_storage[10][1] ),
    .I3(\reg_file.reg_storage[11][1] ),
    .S0(_0955_),
    .S1(_0678_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4869_ (.I0(_0981_),
    .I1(_0985_),
    .I2(_0986_),
    .I3(_0987_),
    .S0(_0874_),
    .S1(_0534_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4870_ (.A1(net76),
    .A2(_0611_),
    .B1(_0613_),
    .B2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4871_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4872_ (.A1(_0980_),
    .A2(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4873_ (.A1(_0895_),
    .A2(_0557_),
    .A3(_0752_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4874_ (.I(_0646_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4875_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(\reg_file.reg_storage[5][0] ),
    .I2(\reg_file.reg_storage[6][0] ),
    .I3(\reg_file.reg_storage[7][0] ),
    .S0(_0709_),
    .S1(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4876_ (.I(\reg_file.reg_storage[1][0] ),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4877_ (.I(_0582_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4878_ (.A1(\reg_file.reg_storage[3][0] ),
    .A2(_0596_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4879_ (.A1(\reg_file.reg_storage[2][0] ),
    .A2(_0852_),
    .B(_0853_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4880_ (.A1(_0995_),
    .A2(_0996_),
    .B1(_0997_),
    .B2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4881_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(\reg_file.reg_storage[13][0] ),
    .I2(\reg_file.reg_storage[14][0] ),
    .I3(\reg_file.reg_storage[15][0] ),
    .S0(_0574_),
    .S1(_0993_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4882_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(\reg_file.reg_storage[9][0] ),
    .I2(\reg_file.reg_storage[10][0] ),
    .I3(\reg_file.reg_storage[11][0] ),
    .S0(_0709_),
    .S1(_0993_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4883_ (.I0(_0994_),
    .I1(_0999_),
    .I2(_1000_),
    .I3(_1001_),
    .S0(_0601_),
    .S1(_0859_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4884_ (.A1(_0548_),
    .A2(_0992_),
    .B1(_1002_),
    .B2(_0861_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4885_ (.I(_1003_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4886_ (.A1(_0489_),
    .A2(_0498_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4887_ (.I(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4888_ (.I(_0732_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4889_ (.I(_0836_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4890_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(\reg_file.reg_storage[3][0] ),
    .S(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4891_ (.I(_0684_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4892_ (.A1(_1010_),
    .A2(\reg_file.reg_storage[1][0] ),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4893_ (.A1(_1007_),
    .A2(_1009_),
    .B(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4894_ (.I(_0530_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4895_ (.I(_0505_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4896_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(\reg_file.reg_storage[5][0] ),
    .I2(\reg_file.reg_storage[6][0] ),
    .I3(\reg_file.reg_storage[7][0] ),
    .S0(_0727_),
    .S1(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4897_ (.A1(_1013_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4898_ (.A1(_0803_),
    .A2(_1012_),
    .B(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4899_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(\reg_file.reg_storage[9][0] ),
    .I2(\reg_file.reg_storage[10][0] ),
    .I3(\reg_file.reg_storage[11][0] ),
    .S0(_0524_),
    .S1(_1014_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4900_ (.A1(_0835_),
    .A2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4901_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(\reg_file.reg_storage[13][0] ),
    .I2(\reg_file.reg_storage[14][0] ),
    .I3(\reg_file.reg_storage[15][0] ),
    .S0(_0727_),
    .S1(_1014_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4902_ (.A1(_1013_),
    .A2(_1020_),
    .B(_0804_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4903_ (.A1(_1019_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4904_ (.A1(_0832_),
    .A2(_1017_),
    .B(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4905_ (.A1(net65),
    .A2(_0672_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4906_ (.A1(_1006_),
    .A2(_1023_),
    .B(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4907_ (.A1(_1004_),
    .A2(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4908_ (.A1(_0540_),
    .A2(_0542_),
    .A3(_0546_),
    .A4(_0568_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4909_ (.A1(_0973_),
    .A2(_0978_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4910_ (.A1(_0538_),
    .A2(_0539_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4911_ (.I(net28),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4912_ (.A1(_0551_),
    .A2(_0480_),
    .A3(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4913_ (.A1(_0758_),
    .A2(_0538_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(_0487_),
    .A2(_0808_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4915_ (.A1(_1031_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4916_ (.A1(_0757_),
    .A2(_1030_),
    .A3(_0539_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4917_ (.A1(_0748_),
    .A2(_1032_),
    .B(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4918_ (.A1(_1029_),
    .A2(_1034_),
    .A3(_1036_),
    .B(_0967_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4919_ (.A1(_1027_),
    .A2(_1028_),
    .B(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4920_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4921_ (.I(_0990_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4922_ (.A1(_1039_),
    .A2(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4923_ (.A1(_0991_),
    .A2(_1026_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4924_ (.A1(_1029_),
    .A2(_1034_),
    .A3(_1036_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4925_ (.A1(_0936_),
    .A2(_0937_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4926_ (.A1(_0945_),
    .A2(_0949_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4927_ (.A1(_1043_),
    .A2(_1044_),
    .B1(_1045_),
    .B2(_1027_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4928_ (.A1(_1046_),
    .A2(net188),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4929_ (.I(_0924_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4930_ (.A1(_0934_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4931_ (.I(_1048_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4932_ (.I(_1050_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4933_ (.I(_0934_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4934_ (.I(_1052_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4935_ (.A1(_1051_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4936_ (.A1(_0965_),
    .A2(_1042_),
    .B1(_1047_),
    .B2(net198),
    .C(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4937_ (.A1(net3),
    .A2(_0752_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4938_ (.A1(_0910_),
    .A2(_0750_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4939_ (.A1(net17),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4940_ (.A1(_1056_),
    .A2(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4941_ (.I0(\reg_file.reg_storage[2][4] ),
    .I1(\reg_file.reg_storage[3][4] ),
    .S(_0885_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4942_ (.A1(_0578_),
    .A2(\reg_file.reg_storage[1][4] ),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4943_ (.A1(_0655_),
    .A2(_1060_),
    .B(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4944_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(\reg_file.reg_storage[5][4] ),
    .I2(\reg_file.reg_storage[6][4] ),
    .I3(\reg_file.reg_storage[7][4] ),
    .S0(_0573_),
    .S1(_0646_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4945_ (.A1(_0974_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4946_ (.A1(_0858_),
    .A2(_1062_),
    .B(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4947_ (.A1(_0664_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4948_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(\reg_file.reg_storage[13][4] ),
    .I2(\reg_file.reg_storage[14][4] ),
    .I3(\reg_file.reg_storage[15][4] ),
    .S0(_0644_),
    .S1(_0763_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4949_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(\reg_file.reg_storage[9][4] ),
    .I2(\reg_file.reg_storage[10][4] ),
    .I3(\reg_file.reg_storage[11][4] ),
    .S0(_0708_),
    .S1(_0969_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4950_ (.I0(_1067_),
    .I1(_1068_),
    .S(_0974_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4951_ (.A1(_0944_),
    .A2(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4952_ (.A1(_1027_),
    .A2(_1066_),
    .A3(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4953_ (.A1(_0641_),
    .A2(_1059_),
    .B(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4954_ (.I(_0630_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4955_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(\reg_file.reg_storage[5][4] ),
    .I2(\reg_file.reg_storage[6][4] ),
    .I3(\reg_file.reg_storage[7][4] ),
    .S0(_1073_),
    .S1(_0632_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4956_ (.I(\reg_file.reg_storage[1][4] ),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4957_ (.I(_0523_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4958_ (.A1(_1076_),
    .A2(\reg_file.reg_storage[3][4] ),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4959_ (.I(_0928_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4960_ (.A1(_1078_),
    .A2(\reg_file.reg_storage[2][4] ),
    .B(_0953_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4961_ (.A1(_0795_),
    .A2(_1075_),
    .B1(_1077_),
    .B2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4962_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(\reg_file.reg_storage[13][4] ),
    .I2(\reg_file.reg_storage[14][4] ),
    .I3(\reg_file.reg_storage[15][4] ),
    .S0(_1008_),
    .S1(_1010_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4963_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(\reg_file.reg_storage[9][4] ),
    .I2(\reg_file.reg_storage[10][4] ),
    .I3(\reg_file.reg_storage[11][4] ),
    .S0(_1008_),
    .S1(_1010_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4964_ (.I0(_1074_),
    .I1(_1080_),
    .I2(_1081_),
    .I3(_1082_),
    .S0(_0531_),
    .S1(_0695_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4965_ (.A1(net91),
    .A2(_0865_),
    .B1(_0614_),
    .B2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4966_ (.A1(_1072_),
    .A2(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4967_ (.I(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4968_ (.I(_0611_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4969_ (.I0(\reg_file.reg_storage[4][6] ),
    .I1(\reg_file.reg_storage[5][6] ),
    .I2(\reg_file.reg_storage[6][6] ),
    .I3(\reg_file.reg_storage[7][6] ),
    .S0(_0631_),
    .S1(_0632_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4970_ (.I(\reg_file.reg_storage[1][6] ),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4971_ (.I(_0502_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4972_ (.A1(_1090_),
    .A2(\reg_file.reg_storage[3][6] ),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4973_ (.A1(_1078_),
    .A2(\reg_file.reg_storage[2][6] ),
    .B(_0953_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4974_ (.A1(_0795_),
    .A2(_1089_),
    .B1(_1091_),
    .B2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4975_ (.I0(\reg_file.reg_storage[12][6] ),
    .I1(\reg_file.reg_storage[13][6] ),
    .I2(\reg_file.reg_storage[14][6] ),
    .I3(\reg_file.reg_storage[15][6] ),
    .S0(_1073_),
    .S1(_1010_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4976_ (.I0(\reg_file.reg_storage[8][6] ),
    .I1(\reg_file.reg_storage[9][6] ),
    .I2(\reg_file.reg_storage[10][6] ),
    .I3(\reg_file.reg_storage[11][6] ),
    .S0(_1073_),
    .S1(_0632_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4977_ (.I0(_1088_),
    .I1(_1093_),
    .I2(_1094_),
    .I3(_1095_),
    .S0(_1013_),
    .S1(_0636_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4978_ (.A1(net93),
    .A2(_1087_),
    .B1(_0726_),
    .B2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4979_ (.A1(net19),
    .A2(_0844_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4980_ (.I0(\reg_file.reg_storage[4][6] ),
    .I1(\reg_file.reg_storage[5][6] ),
    .I2(\reg_file.reg_storage[6][6] ),
    .I3(\reg_file.reg_storage[7][6] ),
    .S0(_0645_),
    .S1(_0647_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4981_ (.A1(_0652_),
    .A2(\reg_file.reg_storage[3][6] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4982_ (.A1(_0654_),
    .A2(\reg_file.reg_storage[2][6] ),
    .B(_0583_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4983_ (.A1(_0649_),
    .A2(_1089_),
    .B1(_1100_),
    .B2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4984_ (.I(_0847_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4985_ (.I0(\reg_file.reg_storage[12][6] ),
    .I1(\reg_file.reg_storage[13][6] ),
    .I2(\reg_file.reg_storage[14][6] ),
    .I3(\reg_file.reg_storage[15][6] ),
    .S0(_0658_),
    .S1(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4986_ (.I0(\reg_file.reg_storage[8][6] ),
    .I1(\reg_file.reg_storage[9][6] ),
    .I2(\reg_file.reg_storage[10][6] ),
    .I3(\reg_file.reg_storage[11][6] ),
    .S0(_0658_),
    .S1(_1103_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4987_ (.I0(_1099_),
    .I1(_1102_),
    .I2(_1104_),
    .I3(_1105_),
    .S0(_0858_),
    .S1(_0664_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4988_ (.A1(_0843_),
    .A2(_1098_),
    .B1(_1106_),
    .B2(_0667_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4989_ (.A1(net192),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4990_ (.A1(net192),
    .A2(_1107_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4991_ (.A1(_1108_),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4992_ (.I(net187),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4993_ (.I0(\reg_file.reg_storage[2][5] ),
    .I1(\reg_file.reg_storage[3][5] ),
    .S(_0630_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4994_ (.I0(\reg_file.reg_storage[1][5] ),
    .I1(_1112_),
    .S(_0786_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4995_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(\reg_file.reg_storage[5][5] ),
    .I2(\reg_file.reg_storage[6][5] ),
    .I3(\reg_file.reg_storage[7][5] ),
    .S0(_0502_),
    .S1(_0684_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4996_ (.A1(_0681_),
    .A2(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4997_ (.A1(_0835_),
    .A2(_1113_),
    .B(_1115_),
    .C(_0627_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4998_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(\reg_file.reg_storage[13][5] ),
    .I2(\reg_file.reg_storage[14][5] ),
    .I3(\reg_file.reg_storage[15][5] ),
    .S0(_0503_),
    .S1(_0786_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4999_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(\reg_file.reg_storage[9][5] ),
    .I2(\reg_file.reg_storage[10][5] ),
    .I3(\reg_file.reg_storage[11][5] ),
    .S0(_0502_),
    .S1(_0678_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5000_ (.A1(_0615_),
    .A2(_1118_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5001_ (.A1(_0742_),
    .A2(_1117_),
    .B(_1119_),
    .C(_0695_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5002_ (.A1(_1116_),
    .A2(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5003_ (.A1(net92),
    .A2(_0612_),
    .B1(_0614_),
    .B2(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5004_ (.A1(net18),
    .A2(_0809_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5005_ (.I(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5006_ (.I(_0847_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5007_ (.I0(\reg_file.reg_storage[4][5] ),
    .I1(\reg_file.reg_storage[5][5] ),
    .I2(\reg_file.reg_storage[6][5] ),
    .I3(\reg_file.reg_storage[7][5] ),
    .S0(_0651_),
    .S1(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5008_ (.I(\reg_file.reg_storage[1][5] ),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5009_ (.A1(_0586_),
    .A2(\reg_file.reg_storage[3][5] ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5010_ (.A1(_0590_),
    .A2(\reg_file.reg_storage[2][5] ),
    .B(_0592_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5011_ (.A1(_0996_),
    .A2(_1127_),
    .B1(_1128_),
    .B2(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5012_ (.I0(\reg_file.reg_storage[12][5] ),
    .I1(\reg_file.reg_storage[13][5] ),
    .I2(\reg_file.reg_storage[14][5] ),
    .I3(\reg_file.reg_storage[15][5] ),
    .S0(_0885_),
    .S1(_0703_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5013_ (.I0(\reg_file.reg_storage[8][5] ),
    .I1(\reg_file.reg_storage[9][5] ),
    .I2(\reg_file.reg_storage[10][5] ),
    .I3(\reg_file.reg_storage[11][5] ),
    .S0(_0651_),
    .S1(_1125_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5014_ (.I0(_1126_),
    .I1(_1130_),
    .I2(_1131_),
    .I3(_1132_),
    .S0(_0974_),
    .S1(_0859_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5015_ (.A1(_0548_),
    .A2(_1124_),
    .B1(_1133_),
    .B2(_0570_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5016_ (.A1(_1122_),
    .A2(_1134_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5017_ (.I(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5018_ (.I(_0684_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5019_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(\reg_file.reg_storage[5][7] ),
    .I2(\reg_file.reg_storage[6][7] ),
    .I3(\reg_file.reg_storage[7][7] ),
    .S0(_1008_),
    .S1(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5020_ (.I(_0519_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5021_ (.I(\reg_file.reg_storage[1][7] ),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5022_ (.A1(_1076_),
    .A2(\reg_file.reg_storage[3][7] ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5023_ (.A1(_0517_),
    .A2(\reg_file.reg_storage[2][7] ),
    .B(_0953_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5024_ (.A1(_1139_),
    .A2(_1140_),
    .B1(_1141_),
    .B2(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5025_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(\reg_file.reg_storage[13][7] ),
    .I2(\reg_file.reg_storage[14][7] ),
    .I3(\reg_file.reg_storage[15][7] ),
    .S0(_0956_),
    .S1(_1137_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5026_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(\reg_file.reg_storage[9][7] ),
    .I2(\reg_file.reg_storage[10][7] ),
    .I3(\reg_file.reg_storage[11][7] ),
    .S0(_0956_),
    .S1(_1137_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5027_ (.I0(_1138_),
    .I1(_1143_),
    .I2(_1144_),
    .I3(_1145_),
    .S0(_0531_),
    .S1(_0695_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5028_ (.A1(net94),
    .A2(_0865_),
    .B1(_0614_),
    .B2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5029_ (.A1(net20),
    .A2(_0809_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5030_ (.I(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5031_ (.I(_0969_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5032_ (.I0(\reg_file.reg_storage[4][7] ),
    .I1(\reg_file.reg_storage[5][7] ),
    .I2(\reg_file.reg_storage[6][7] ),
    .I3(\reg_file.reg_storage[7][7] ),
    .S0(_0886_),
    .S1(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5033_ (.I(_0853_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5034_ (.I(_0754_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5035_ (.A1(_1153_),
    .A2(\reg_file.reg_storage[3][7] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5036_ (.A1(_0654_),
    .A2(\reg_file.reg_storage[2][7] ),
    .B(_0655_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5037_ (.A1(_1152_),
    .A2(_1140_),
    .B1(_1154_),
    .B2(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5038_ (.I(_0646_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5039_ (.I0(\reg_file.reg_storage[12][7] ),
    .I1(\reg_file.reg_storage[13][7] ),
    .I2(\reg_file.reg_storage[14][7] ),
    .I3(\reg_file.reg_storage[15][7] ),
    .S0(_0754_),
    .S1(_1157_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5040_ (.I0(\reg_file.reg_storage[8][7] ),
    .I1(\reg_file.reg_storage[9][7] ),
    .I2(\reg_file.reg_storage[10][7] ),
    .I3(\reg_file.reg_storage[11][7] ),
    .S0(_0886_),
    .S1(_1157_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5041_ (.I0(_1151_),
    .I1(_1156_),
    .I2(_1158_),
    .I3(_1159_),
    .S0(_0662_),
    .S1(_0775_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5042_ (.A1(_0641_),
    .A2(_1149_),
    .B1(_1160_),
    .B2(_0667_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5043_ (.A1(_1161_),
    .A2(_1147_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5044_ (.I(_1162_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _5045_ (.A1(_1086_),
    .A2(_1111_),
    .A3(_1136_),
    .A4(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5046_ (.A1(_1108_),
    .A2(_1109_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5047_ (.A1(net3),
    .A2(_0752_),
    .B1(_1057_),
    .B2(net17),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _5048_ (.A1(_1027_),
    .A2(_1066_),
    .A3(_1070_),
    .B1(_1166_),
    .B2(_1043_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5049_ (.I(_1167_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5050_ (.A1(_1116_),
    .A2(_1120_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5051_ (.A1(net92),
    .A2(_0672_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5052_ (.A1(_1006_),
    .A2(_1169_),
    .B(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5053_ (.I(_1134_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5054_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5055_ (.A1(_1168_),
    .A2(_1084_),
    .A3(_1135_),
    .B(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5056_ (.I(net192),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5057_ (.A1(_1175_),
    .A2(_1107_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5058_ (.A1(_1165_),
    .A2(_1174_),
    .B(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5059_ (.I(_1147_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5060_ (.I(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5061_ (.I(_1161_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5062_ (.A1(_1179_),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5063_ (.A1(_1055_),
    .A2(_1164_),
    .B1(_1177_),
    .B2(_1163_),
    .C(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5064_ (.I(_1006_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5065_ (.A1(_0873_),
    .A2(_0879_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5066_ (.I(_0672_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(net95),
    .A2(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5068_ (.A1(_1183_),
    .A2(_1184_),
    .B(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5069_ (.A1(_1187_),
    .A2(_0903_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5070_ (.A1(_0908_),
    .A2(_1182_),
    .B(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5071_ (.I(_1005_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5072_ (.A1(_0833_),
    .A2(_0840_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5073_ (.A1(net96),
    .A2(_0612_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5074_ (.A1(_1190_),
    .A2(_1191_),
    .B(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5075_ (.I(_0862_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5076_ (.A1(_1193_),
    .A2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5077_ (.A1(_0864_),
    .A2(_1189_),
    .B(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5078_ (.I(_0807_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5079_ (.A1(_1197_),
    .A2(_0820_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5080_ (.A1(_0825_),
    .A2(_1196_),
    .B(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5081_ (.I(_0744_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5082_ (.A1(_1200_),
    .A2(_0778_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5083_ (.A1(_0782_),
    .A2(_1199_),
    .B(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5084_ (.A1(_0689_),
    .A2(_0697_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5085_ (.A1(_0671_),
    .A2(_1185_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5086_ (.A1(_1183_),
    .A2(_1203_),
    .B(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5087_ (.A1(_1205_),
    .A2(_0720_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5088_ (.A1(_0724_),
    .A2(_1202_),
    .B(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5089_ (.A1(_0628_),
    .A2(_0637_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5090_ (.A1(net69),
    .A2(_0612_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5091_ (.A1(_1190_),
    .A2(_1208_),
    .B(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5092_ (.I(_0668_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5093_ (.A1(_1210_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5094_ (.A1(_0670_),
    .A2(_1207_),
    .B(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5095_ (.I(_1029_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5096_ (.A1(_1214_),
    .A2(_1034_),
    .A3(_0544_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5097_ (.I(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5098_ (.A1(_0481_),
    .A2(_0543_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5099_ (.I(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5100_ (.A1(net24),
    .A2(_1216_),
    .B1(_1218_),
    .B2(_0550_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5101_ (.I(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5102_ (.A1(net6),
    .A2(_1216_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5103_ (.I(_1221_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5104_ (.I(_1217_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5105_ (.A1(net5),
    .A2(_1216_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5106_ (.A1(_1223_),
    .A2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5107_ (.A1(net6),
    .A2(net5),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5108_ (.A1(net4),
    .A2(_1215_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5109_ (.A1(_1223_),
    .A2(_1226_),
    .B(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5110_ (.A1(_1225_),
    .A2(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5111_ (.A1(_1222_),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5112_ (.A1(_1220_),
    .A2(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5113_ (.I(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5114_ (.A1(_0610_),
    .A2(_1213_),
    .B(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5115_ (.A1(_0610_),
    .A2(net216),
    .B(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5116_ (.A1(net5),
    .A2(_1215_),
    .B(_1218_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5117_ (.A1(_1235_),
    .A2(_1228_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5118_ (.A1(_1222_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5119_ (.I(_1237_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5120_ (.I(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5121_ (.I(_1048_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5122_ (.I(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5123_ (.I(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5124_ (.I(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5125_ (.I(_1168_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_1243_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5127_ (.I(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5128_ (.I(_0951_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5129_ (.I(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5130_ (.I(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5131_ (.I(_1249_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5132_ (.I(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5133_ (.I(_1039_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5134_ (.I(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5135_ (.I(_1253_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5136_ (.I(_1003_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5137_ (.I(_1255_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5138_ (.I(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5139_ (.I(_1087_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5140_ (.I(_0726_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5141_ (.I(_1076_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5142_ (.I(_0870_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5143_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(\reg_file.reg_storage[5][30] ),
    .I2(\reg_file.reg_storage[6][30] ),
    .I3(\reg_file.reg_storage[7][30] ),
    .S0(_1260_),
    .S1(_1261_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5144_ (.I(_0733_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5145_ (.I(\reg_file.reg_storage[1][30] ),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5146_ (.I(_1090_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5147_ (.A1(_1265_),
    .A2(\reg_file.reg_storage[3][30] ),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5148_ (.I(_1078_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5149_ (.I(_0510_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5150_ (.A1(_1267_),
    .A2(\reg_file.reg_storage[2][30] ),
    .B(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5151_ (.A1(_1263_),
    .A2(_1264_),
    .B1(_1266_),
    .B2(_1269_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5152_ (.I(_0524_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5153_ (.I(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5154_ (.I(_1137_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5155_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(\reg_file.reg_storage[13][30] ),
    .I2(\reg_file.reg_storage[14][30] ),
    .I3(\reg_file.reg_storage[15][30] ),
    .S0(_1272_),
    .S1(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5156_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(\reg_file.reg_storage[9][30] ),
    .I2(\reg_file.reg_storage[10][30] ),
    .I3(\reg_file.reg_storage[11][30] ),
    .S0(_1272_),
    .S1(_1261_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5157_ (.I(_0535_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5158_ (.I0(_1262_),
    .I1(_1270_),
    .I2(_1274_),
    .I3(_1275_),
    .S0(_0690_),
    .S1(_1276_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5159_ (.A1(net88),
    .A2(_1258_),
    .B1(_1259_),
    .B2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5160_ (.I(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5161_ (.A1(_1257_),
    .A2(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5162_ (.I(_1255_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5163_ (.I(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5164_ (.I(_0491_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5165_ (.I(_1090_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5166_ (.I(_0619_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5167_ (.I(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5168_ (.I0(\reg_file.reg_storage[4][31] ),
    .I1(\reg_file.reg_storage[5][31] ),
    .I2(\reg_file.reg_storage[6][31] ),
    .I3(\reg_file.reg_storage[7][31] ),
    .S0(_1284_),
    .S1(_1286_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5169_ (.I(\reg_file.reg_storage[1][31] ),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5170_ (.A1(_1265_),
    .A2(\reg_file.reg_storage[3][31] ),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5171_ (.I(_1139_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5172_ (.A1(_1267_),
    .A2(\reg_file.reg_storage[2][31] ),
    .B(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5173_ (.A1(_1263_),
    .A2(_1288_),
    .B1(_1289_),
    .B2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5174_ (.I0(\reg_file.reg_storage[12][31] ),
    .I1(\reg_file.reg_storage[13][31] ),
    .I2(\reg_file.reg_storage[14][31] ),
    .I3(\reg_file.reg_storage[15][31] ),
    .S0(_1284_),
    .S1(_1286_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5175_ (.I0(\reg_file.reg_storage[8][31] ),
    .I1(\reg_file.reg_storage[9][31] ),
    .I2(\reg_file.reg_storage[10][31] ),
    .I3(\reg_file.reg_storage[11][31] ),
    .S0(_1284_),
    .S1(_1286_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5176_ (.I(_0804_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5177_ (.I(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5178_ (.I0(_1287_),
    .I1(_1292_),
    .I2(_1293_),
    .I3(_1294_),
    .S0(_0875_),
    .S1(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5179_ (.A1(net89),
    .A2(_1283_),
    .B1(_1259_),
    .B2(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5180_ (.I(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5181_ (.A1(_1282_),
    .A2(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5182_ (.A1(_1254_),
    .A2(_1280_),
    .A3(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5183_ (.A1(_1251_),
    .A2(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5184_ (.I(_1243_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5185_ (.I(net205),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5186_ (.I(_1304_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5187_ (.I(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5188_ (.I(_0980_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5189_ (.I(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5190_ (.I(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5191_ (.I(_1004_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5192_ (.I(_1190_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5193_ (.I(_0799_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5194_ (.I0(\reg_file.reg_storage[4][27] ),
    .I1(\reg_file.reg_storage[5][27] ),
    .I2(\reg_file.reg_storage[6][27] ),
    .I3(\reg_file.reg_storage[7][27] ),
    .S0(_0785_),
    .S1(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5195_ (.I(\reg_file.reg_storage[1][27] ),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5196_ (.A1(_0792_),
    .A2(\reg_file.reg_storage[3][27] ),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5197_ (.A1(_0794_),
    .A2(\reg_file.reg_storage[2][27] ),
    .B(_1139_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5198_ (.A1(_0789_),
    .A2(_1314_),
    .B1(_1315_),
    .B2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5199_ (.I(_0531_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5200_ (.I0(_1313_),
    .I1(_1317_),
    .S(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5201_ (.A1(_1296_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5202_ (.I(_0729_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5203_ (.I0(\reg_file.reg_storage[12][27] ),
    .I1(\reg_file.reg_storage[13][27] ),
    .I2(\reg_file.reg_storage[14][27] ),
    .I3(\reg_file.reg_storage[15][27] ),
    .S0(_0676_),
    .S1(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5204_ (.I0(\reg_file.reg_storage[8][27] ),
    .I1(\reg_file.reg_storage[9][27] ),
    .I2(\reg_file.reg_storage[10][27] ),
    .I3(\reg_file.reg_storage[11][27] ),
    .S0(_0728_),
    .S1(_1321_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5205_ (.I0(_1322_),
    .I1(_1323_),
    .S(_0629_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5206_ (.A1(_0688_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5207_ (.A1(net84),
    .A2(_1283_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5208_ (.A1(_1311_),
    .A2(_1320_),
    .A3(_1325_),
    .B(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5209_ (.I0(\reg_file.reg_storage[4][26] ),
    .I1(\reg_file.reg_storage[5][26] ),
    .I2(\reg_file.reg_storage[6][26] ),
    .I3(\reg_file.reg_storage[7][26] ),
    .S0(_0691_),
    .S1(_0679_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5210_ (.I(\reg_file.reg_storage[1][26] ),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5211_ (.A1(_1284_),
    .A2(\reg_file.reg_storage[3][26] ),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5212_ (.I(_0517_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5213_ (.A1(_1331_),
    .A2(\reg_file.reg_storage[2][26] ),
    .B(_1007_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5214_ (.A1(_1268_),
    .A2(_1329_),
    .B1(_1330_),
    .B2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5215_ (.I(_1073_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5216_ (.I(_0799_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5217_ (.I0(\reg_file.reg_storage[12][26] ),
    .I1(\reg_file.reg_storage[13][26] ),
    .I2(\reg_file.reg_storage[14][26] ),
    .I3(\reg_file.reg_storage[15][26] ),
    .S0(_1334_),
    .S1(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5218_ (.I0(\reg_file.reg_storage[8][26] ),
    .I1(\reg_file.reg_storage[9][26] ),
    .I2(\reg_file.reg_storage[10][26] ),
    .I3(\reg_file.reg_storage[11][26] ),
    .S0(_1334_),
    .S1(_1335_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5219_ (.I(_1013_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5220_ (.I0(_1328_),
    .I1(_1333_),
    .I2(_1336_),
    .I3(_1337_),
    .S0(_1338_),
    .S1(_0805_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5221_ (.A1(net83),
    .A2(_1185_),
    .B1(_0674_),
    .B2(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5222_ (.I(_1340_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5223_ (.A1(_1281_),
    .A2(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5224_ (.A1(_1310_),
    .A2(_1327_),
    .B(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5225_ (.A1(_1309_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5226_ (.I(_1256_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5227_ (.A1(net86),
    .A2(_0673_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5228_ (.I(_0799_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5229_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(\reg_file.reg_storage[5][29] ),
    .I2(\reg_file.reg_storage[6][29] ),
    .I3(\reg_file.reg_storage[7][29] ),
    .S0(_1090_),
    .S1(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5230_ (.I(\reg_file.reg_storage[1][29] ),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5231_ (.A1(_1272_),
    .A2(\reg_file.reg_storage[3][29] ),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5232_ (.A1(_1331_),
    .A2(\reg_file.reg_storage[2][29] ),
    .B(_1007_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5233_ (.A1(_1268_),
    .A2(_1349_),
    .B1(_1350_),
    .B2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5234_ (.I(_0956_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5235_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(\reg_file.reg_storage[13][29] ),
    .I2(\reg_file.reg_storage[14][29] ),
    .I3(\reg_file.reg_storage[15][29] ),
    .S0(_1353_),
    .S1(_1312_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5236_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(\reg_file.reg_storage[9][29] ),
    .I2(\reg_file.reg_storage[10][29] ),
    .I3(\reg_file.reg_storage[11][29] ),
    .S0(_1353_),
    .S1(_1347_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5237_ (.I0(_1348_),
    .I1(_1352_),
    .I2(_1354_),
    .I3(_1355_),
    .S0(_1318_),
    .S1(_0805_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5238_ (.A1(_0674_),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5239_ (.A1(_1346_),
    .A2(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5240_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5241_ (.A1(_1345_),
    .A2(_1359_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5242_ (.I(_0506_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5243_ (.I0(\reg_file.reg_storage[4][28] ),
    .I1(\reg_file.reg_storage[5][28] ),
    .I2(\reg_file.reg_storage[6][28] ),
    .I3(\reg_file.reg_storage[7][28] ),
    .S0(_0504_),
    .S1(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5244_ (.I(\reg_file.reg_storage[1][28] ),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5245_ (.A1(_0792_),
    .A2(\reg_file.reg_storage[3][28] ),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5246_ (.A1(_0518_),
    .A2(\reg_file.reg_storage[2][28] ),
    .B(_0520_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5247_ (.A1(_0511_),
    .A2(_1363_),
    .B1(_1364_),
    .B2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5248_ (.I0(\reg_file.reg_storage[12][28] ),
    .I1(\reg_file.reg_storage[13][28] ),
    .I2(\reg_file.reg_storage[14][28] ),
    .I3(\reg_file.reg_storage[15][28] ),
    .S0(_0525_),
    .S1(_0526_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5249_ (.I0(\reg_file.reg_storage[8][28] ),
    .I1(\reg_file.reg_storage[9][28] ),
    .I2(\reg_file.reg_storage[10][28] ),
    .I3(\reg_file.reg_storage[11][28] ),
    .S0(_0525_),
    .S1(_0507_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5250_ (.I0(_1362_),
    .I1(_1366_),
    .I2(_1367_),
    .I3(_1368_),
    .S0(_0532_),
    .S1(_1295_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5251_ (.A1(net85),
    .A2(_0491_),
    .B1(_0783_),
    .B2(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5252_ (.I(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5253_ (.A1(_1257_),
    .A2(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5254_ (.I(_1253_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5255_ (.A1(_1360_),
    .A2(_1372_),
    .B(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5256_ (.A1(_1344_),
    .A2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5257_ (.I(_1247_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5258_ (.I(_1376_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5259_ (.I(_1004_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5260_ (.I0(\reg_file.reg_storage[4][23] ),
    .I1(\reg_file.reg_storage[5][23] ),
    .I2(\reg_file.reg_storage[6][23] ),
    .I3(\reg_file.reg_storage[7][23] ),
    .S0(_0515_),
    .S1(_1273_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5261_ (.I(\reg_file.reg_storage[1][23] ),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5262_ (.A1(_1265_),
    .A2(\reg_file.reg_storage[3][23] ),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5263_ (.A1(_1331_),
    .A2(\reg_file.reg_storage[2][23] ),
    .B(_0511_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5264_ (.A1(_1290_),
    .A2(_1380_),
    .B1(_1381_),
    .B2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5265_ (.I0(\reg_file.reg_storage[12][23] ),
    .I1(\reg_file.reg_storage[13][23] ),
    .I2(\reg_file.reg_storage[14][23] ),
    .I3(\reg_file.reg_storage[15][23] ),
    .S0(_0736_),
    .S1(_1273_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5266_ (.I0(\reg_file.reg_storage[8][23] ),
    .I1(\reg_file.reg_storage[9][23] ),
    .I2(\reg_file.reg_storage[10][23] ),
    .I3(\reg_file.reg_storage[11][23] ),
    .S0(_0515_),
    .S1(_1273_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5267_ (.I(_0681_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5268_ (.I0(_1379_),
    .I1(_1383_),
    .I2(_1384_),
    .I3(_1385_),
    .S0(_1386_),
    .S1(_0696_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5269_ (.A1(net80),
    .A2(_1258_),
    .B1(_1259_),
    .B2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5270_ (.I(net175),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5271_ (.I(_1004_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5272_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(\reg_file.reg_storage[5][22] ),
    .I2(\reg_file.reg_storage[6][22] ),
    .I3(\reg_file.reg_storage[7][22] ),
    .S0(_1076_),
    .S1(_1312_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5273_ (.I(\reg_file.reg_storage[1][22] ),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_1272_),
    .A2(\reg_file.reg_storage[3][22] ),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5275_ (.A1(_0794_),
    .A2(\reg_file.reg_storage[2][22] ),
    .B(_0795_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5276_ (.A1(_0789_),
    .A2(_1392_),
    .B1(_1393_),
    .B2(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5277_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(\reg_file.reg_storage[13][22] ),
    .I2(\reg_file.reg_storage[14][22] ),
    .I3(\reg_file.reg_storage[15][22] ),
    .S0(_0785_),
    .S1(_0787_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5278_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(\reg_file.reg_storage[9][22] ),
    .I2(\reg_file.reg_storage[10][22] ),
    .I3(\reg_file.reg_storage[11][22] ),
    .S0(_0785_),
    .S1(_1312_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5279_ (.I0(_1391_),
    .I1(_1395_),
    .I2(_1396_),
    .I3(_1397_),
    .S0(_0803_),
    .S1(_0805_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5280_ (.A1(net79),
    .A2(_0673_),
    .B1(_0783_),
    .B2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5281_ (.I(_1399_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_1390_),
    .A2(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5283_ (.A1(_1378_),
    .A2(_1389_),
    .B(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5284_ (.I(_1006_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5285_ (.I(_0503_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5286_ (.I0(\reg_file.reg_storage[2][25] ),
    .I1(\reg_file.reg_storage[3][25] ),
    .S(_1404_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5287_ (.A1(_0800_),
    .A2(\reg_file.reg_storage[1][25] ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5288_ (.A1(_0789_),
    .A2(_1405_),
    .B(_1406_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5289_ (.I0(\reg_file.reg_storage[4][25] ),
    .I1(\reg_file.reg_storage[5][25] ),
    .I2(\reg_file.reg_storage[6][25] ),
    .I3(\reg_file.reg_storage[7][25] ),
    .S0(_0735_),
    .S1(_0870_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5290_ (.A1(_1318_),
    .A2(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5291_ (.A1(_1386_),
    .A2(_1407_),
    .B(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5292_ (.A1(_1276_),
    .A2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5293_ (.I(_0832_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5294_ (.I0(\reg_file.reg_storage[12][25] ),
    .I1(\reg_file.reg_storage[13][25] ),
    .I2(\reg_file.reg_storage[14][25] ),
    .I3(\reg_file.reg_storage[15][25] ),
    .S0(_0676_),
    .S1(_1321_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5295_ (.I0(\reg_file.reg_storage[8][25] ),
    .I1(\reg_file.reg_storage[9][25] ),
    .I2(\reg_file.reg_storage[10][25] ),
    .I3(\reg_file.reg_storage[11][25] ),
    .S0(_0728_),
    .S1(_0730_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5296_ (.I0(_1413_),
    .I1(_1414_),
    .S(_0629_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5297_ (.A1(_1412_),
    .A2(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5298_ (.A1(net82),
    .A2(_1087_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5299_ (.A1(_1403_),
    .A2(_1411_),
    .A3(_1416_),
    .B(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5300_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5301_ (.A1(_1256_),
    .A2(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5302_ (.I(_1255_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5303_ (.I0(\reg_file.reg_storage[2][24] ),
    .I1(\reg_file.reg_storage[3][24] ),
    .S(_0691_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5304_ (.A1(_0679_),
    .A2(\reg_file.reg_storage[1][24] ),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5305_ (.A1(_1290_),
    .A2(_1422_),
    .B(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5306_ (.I0(\reg_file.reg_storage[4][24] ),
    .I1(\reg_file.reg_storage[5][24] ),
    .I2(\reg_file.reg_storage[6][24] ),
    .I3(\reg_file.reg_storage[7][24] ),
    .S0(_0504_),
    .S1(_1361_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5307_ (.A1(_1338_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5308_ (.A1(_0875_),
    .A2(_1424_),
    .B(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5309_ (.A1(_1427_),
    .A2(_1296_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5310_ (.I0(\reg_file.reg_storage[12][24] ),
    .I1(\reg_file.reg_storage[13][24] ),
    .I2(\reg_file.reg_storage[14][24] ),
    .I3(\reg_file.reg_storage[15][24] ),
    .S0(_1353_),
    .S1(_1347_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5311_ (.I0(\reg_file.reg_storage[8][24] ),
    .I1(\reg_file.reg_storage[9][24] ),
    .I2(\reg_file.reg_storage[10][24] ),
    .I3(\reg_file.reg_storage[11][24] ),
    .S0(_1353_),
    .S1(_1347_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5312_ (.I0(_1429_),
    .I1(_1430_),
    .S(_1338_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5313_ (.A1(_1412_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5314_ (.A1(_1403_),
    .A2(_1428_),
    .A3(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5315_ (.A1(net81),
    .A2(_1283_),
    .B(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5316_ (.A1(_1421_),
    .A2(net212),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(_1420_),
    .A2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5318_ (.I0(_1402_),
    .I1(_1436_),
    .S(_1253_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5319_ (.A1(_1377_),
    .A2(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5320_ (.A1(_1306_),
    .A2(_1375_),
    .B(_1438_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5321_ (.I(_1240_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5322_ (.I(_1440_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5323_ (.I(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5324_ (.I(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5325_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(\reg_file.reg_storage[5][15] ),
    .I2(\reg_file.reg_storage[6][15] ),
    .I3(\reg_file.reg_storage[7][15] ),
    .S0(_1404_),
    .S1(_1361_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5326_ (.I(\reg_file.reg_storage[1][15] ),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5327_ (.A1(_0792_),
    .A2(\reg_file.reg_storage[3][15] ),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5328_ (.A1(_0794_),
    .A2(\reg_file.reg_storage[2][15] ),
    .B(_1139_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5329_ (.A1(_0511_),
    .A2(_1445_),
    .B1(_1446_),
    .B2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5330_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(\reg_file.reg_storage[13][15] ),
    .I2(\reg_file.reg_storage[14][15] ),
    .I3(\reg_file.reg_storage[15][15] ),
    .S0(_0504_),
    .S1(_0507_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5331_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(\reg_file.reg_storage[9][15] ),
    .I2(\reg_file.reg_storage[10][15] ),
    .I3(\reg_file.reg_storage[11][15] ),
    .S0(_1404_),
    .S1(_1361_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5332_ (.I0(_1444_),
    .I1(_1448_),
    .I2(_1449_),
    .I3(_1450_),
    .S0(_0532_),
    .S1(_1295_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5333_ (.A1(net71),
    .A2(_0491_),
    .B1(_0783_),
    .B2(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5334_ (.I(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5335_ (.I(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5336_ (.A1(net224),
    .A2(_1421_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5337_ (.A1(_1378_),
    .A2(_1454_),
    .B(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5338_ (.I0(\reg_file.reg_storage[4][17] ),
    .I1(\reg_file.reg_storage[5][17] ),
    .I2(\reg_file.reg_storage[6][17] ),
    .I3(\reg_file.reg_storage[7][17] ),
    .S0(_0631_),
    .S1(_0685_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5339_ (.A1(_0682_),
    .A2(_1457_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5340_ (.A1(_0676_),
    .A2(\reg_file.reg_storage[3][17] ),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5341_ (.A1(_1331_),
    .A2(\reg_file.reg_storage[2][17] ),
    .B(_1459_),
    .C(_1007_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5342_ (.A1(_0868_),
    .A2(\reg_file.reg_storage[1][17] ),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5343_ (.A1(_1460_),
    .A2(_1461_),
    .B(_1318_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5344_ (.A1(_1458_),
    .A2(_1462_),
    .B(_0696_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5345_ (.I0(\reg_file.reg_storage[12][17] ),
    .I1(\reg_file.reg_storage[13][17] ),
    .I2(\reg_file.reg_storage[14][17] ),
    .I3(\reg_file.reg_storage[15][17] ),
    .S0(_0791_),
    .S1(_0620_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5346_ (.A1(_0629_),
    .A2(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5347_ (.I0(\reg_file.reg_storage[8][17] ),
    .I1(\reg_file.reg_storage[9][17] ),
    .I2(\reg_file.reg_storage[10][17] ),
    .I3(\reg_file.reg_storage[11][17] ),
    .S0(_0683_),
    .S1(_0685_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5348_ (.A1(_0616_),
    .A2(_1466_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5349_ (.A1(_1465_),
    .A2(_1467_),
    .B(_0688_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5350_ (.A1(net73),
    .A2(_0865_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5351_ (.A1(_1190_),
    .A2(_1463_),
    .A3(_1468_),
    .B(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5352_ (.I0(\reg_file.reg_storage[2][16] ),
    .I1(\reg_file.reg_storage[3][16] ),
    .S(_0736_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5353_ (.A1(_0868_),
    .A2(\reg_file.reg_storage[1][16] ),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5354_ (.A1(_1290_),
    .A2(_1471_),
    .B(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5355_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(\reg_file.reg_storage[5][16] ),
    .I2(\reg_file.reg_storage[6][16] ),
    .I3(\reg_file.reg_storage[7][16] ),
    .S0(_0798_),
    .S1(_0787_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5356_ (.A1(_1386_),
    .A2(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5357_ (.A1(_0875_),
    .A2(_1473_),
    .B(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5358_ (.A1(_1296_),
    .A2(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5359_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(\reg_file.reg_storage[13][16] ),
    .I2(\reg_file.reg_storage[14][16] ),
    .I3(\reg_file.reg_storage[15][16] ),
    .S0(_1334_),
    .S1(_1335_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5360_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(\reg_file.reg_storage[9][16] ),
    .I2(\reg_file.reg_storage[10][16] ),
    .I3(\reg_file.reg_storage[11][16] ),
    .S0(_1334_),
    .S1(_1335_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5361_ (.I0(_1478_),
    .I1(_1479_),
    .S(_1338_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5362_ (.A1(_1412_),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5363_ (.A1(_1183_),
    .A2(_1477_),
    .A3(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5364_ (.A1(net72),
    .A2(_1283_),
    .B(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(_1421_),
    .A2(net186),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5366_ (.A1(_1378_),
    .A2(_1470_),
    .B(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5367_ (.I(_1252_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5368_ (.I(_1486_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5369_ (.I0(_1456_),
    .I1(_1485_),
    .S(_1487_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5370_ (.I0(\reg_file.reg_storage[4][19] ),
    .I1(\reg_file.reg_storage[5][19] ),
    .I2(\reg_file.reg_storage[6][19] ),
    .I3(\reg_file.reg_storage[7][19] ),
    .S0(_1260_),
    .S1(_1286_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5371_ (.I(\reg_file.reg_storage[1][19] ),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5372_ (.A1(_1265_),
    .A2(\reg_file.reg_storage[3][19] ),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5373_ (.A1(_1267_),
    .A2(\reg_file.reg_storage[2][19] ),
    .B(_1268_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5374_ (.A1(_1263_),
    .A2(_1490_),
    .B1(_1491_),
    .B2(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5375_ (.I0(\reg_file.reg_storage[12][19] ),
    .I1(\reg_file.reg_storage[13][19] ),
    .I2(\reg_file.reg_storage[14][19] ),
    .I3(\reg_file.reg_storage[15][19] ),
    .S0(_1260_),
    .S1(_1261_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5376_ (.I0(\reg_file.reg_storage[8][19] ),
    .I1(\reg_file.reg_storage[9][19] ),
    .I2(\reg_file.reg_storage[10][19] ),
    .I3(\reg_file.reg_storage[11][19] ),
    .S0(_1260_),
    .S1(_1261_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5377_ (.I0(_1489_),
    .I1(_1493_),
    .I2(_1494_),
    .I3(_1495_),
    .S0(_0690_),
    .S1(_1276_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5378_ (.A1(net75),
    .A2(_1258_),
    .B1(_1259_),
    .B2(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5379_ (.I(_1497_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5380_ (.I0(\reg_file.reg_storage[4][18] ),
    .I1(\reg_file.reg_storage[5][18] ),
    .I2(\reg_file.reg_storage[6][18] ),
    .I3(\reg_file.reg_storage[7][18] ),
    .S0(_1271_),
    .S1(_0526_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5381_ (.I(\reg_file.reg_storage[1][18] ),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5382_ (.A1(_0515_),
    .A2(\reg_file.reg_storage[3][18] ),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5383_ (.A1(_0518_),
    .A2(\reg_file.reg_storage[2][18] ),
    .B(_0520_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5384_ (.A1(_0733_),
    .A2(_1500_),
    .B1(_1501_),
    .B2(_1502_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5385_ (.I0(\reg_file.reg_storage[12][18] ),
    .I1(\reg_file.reg_storage[13][18] ),
    .I2(\reg_file.reg_storage[14][18] ),
    .I3(\reg_file.reg_storage[15][18] ),
    .S0(_1271_),
    .S1(_1321_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5386_ (.I0(\reg_file.reg_storage[8][18] ),
    .I1(\reg_file.reg_storage[9][18] ),
    .I2(\reg_file.reg_storage[10][18] ),
    .I3(\reg_file.reg_storage[11][18] ),
    .S0(_1271_),
    .S1(_0526_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5387_ (.I0(_1499_),
    .I1(_1503_),
    .I2(_1504_),
    .I3(_1505_),
    .S0(_0682_),
    .S1(_0535_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5388_ (.A1(net74),
    .A2(_0725_),
    .B1(_0501_),
    .B2(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5389_ (.I(_1507_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5390_ (.I0(_1498_),
    .I1(_1508_),
    .S(_1281_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5391_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(\reg_file.reg_storage[5][21] ),
    .I2(\reg_file.reg_storage[6][21] ),
    .I3(\reg_file.reg_storage[7][21] ),
    .S0(_0514_),
    .S1(_1285_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5392_ (.I(\reg_file.reg_storage[1][21] ),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5393_ (.A1(_0691_),
    .A2(\reg_file.reg_storage[3][21] ),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5394_ (.A1(_1078_),
    .A2(\reg_file.reg_storage[2][21] ),
    .B(_0510_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5395_ (.A1(_0733_),
    .A2(_1511_),
    .B1(_1512_),
    .B2(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5396_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(\reg_file.reg_storage[13][21] ),
    .I2(\reg_file.reg_storage[14][21] ),
    .I3(\reg_file.reg_storage[15][21] ),
    .S0(_0735_),
    .S1(_1285_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5397_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(\reg_file.reg_storage[9][21] ),
    .I2(\reg_file.reg_storage[10][21] ),
    .I3(\reg_file.reg_storage[11][21] ),
    .S0(_0514_),
    .S1(_1285_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5398_ (.I0(_1510_),
    .I1(_1514_),
    .I2(_1515_),
    .I3(_1516_),
    .S0(_0742_),
    .S1(_0636_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5399_ (.A1(net78),
    .A2(_1087_),
    .B1(_0726_),
    .B2(_1517_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5400_ (.I0(\reg_file.reg_storage[2][20] ),
    .I1(\reg_file.reg_storage[3][20] ),
    .S(_0791_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5401_ (.I0(\reg_file.reg_storage[1][20] ),
    .I1(_1519_),
    .S(_0787_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5402_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(\reg_file.reg_storage[5][20] ),
    .I2(\reg_file.reg_storage[6][20] ),
    .I3(\reg_file.reg_storage[7][20] ),
    .S0(_0503_),
    .S1(_0786_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5403_ (.A1(_0742_),
    .A2(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5404_ (.A1(_0675_),
    .A2(_1520_),
    .B(_1522_),
    .C(_0832_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5405_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(\reg_file.reg_storage[13][20] ),
    .I2(\reg_file.reg_storage[14][20] ),
    .I3(\reg_file.reg_storage[15][20] ),
    .S0(_1404_),
    .S1(_0800_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5406_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(\reg_file.reg_storage[9][20] ),
    .I2(\reg_file.reg_storage[10][20] ),
    .I3(\reg_file.reg_storage[11][20] ),
    .S0(_0524_),
    .S1(_1014_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5407_ (.A1(_0835_),
    .A2(_1525_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5408_ (.A1(_1386_),
    .A2(_1524_),
    .B(_1526_),
    .C(_1295_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5409_ (.A1(_1527_),
    .A2(_1523_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5410_ (.A1(net77),
    .A2(_0725_),
    .B1(_0501_),
    .B2(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5411_ (.I0(net220),
    .I1(net177),
    .S(_1421_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5412_ (.I0(_1509_),
    .I1(_1530_),
    .S(_1487_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5413_ (.I0(_1488_),
    .I1(_1531_),
    .S(_1306_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5414_ (.A1(_1443_),
    .A2(_1532_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5415_ (.I(_1072_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5416_ (.I(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5417_ (.I(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5418_ (.I(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5419_ (.A1(_1303_),
    .A2(_1439_),
    .B(_1533_),
    .C(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5420_ (.A1(_1246_),
    .A2(_1302_),
    .B(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5421_ (.A1(_1219_),
    .A2(_1221_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5422_ (.A1(_1236_),
    .A2(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5423_ (.A1(_1168_),
    .A2(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5424_ (.I(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5425_ (.I(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5426_ (.I(_1051_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5427_ (.I(_1545_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5428_ (.A1(_1193_),
    .A2(_1281_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5429_ (.A1(_0807_),
    .A2(_1390_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5430_ (.A1(_1547_),
    .A2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5431_ (.A1(_1345_),
    .A2(_1179_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5432_ (.A1(_0881_),
    .A2(_1310_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5433_ (.A1(_1550_),
    .A2(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5434_ (.I0(_1549_),
    .I1(_1552_),
    .S(_1486_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5435_ (.A1(net221),
    .A2(_1256_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5436_ (.A1(_1455_),
    .A2(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5437_ (.I(_1310_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5438_ (.I(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5439_ (.A1(_0699_),
    .A2(_1390_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5440_ (.A1(_1200_),
    .A2(_1557_),
    .B(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5441_ (.I0(_1555_),
    .I1(_1559_),
    .S(_1253_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5442_ (.I0(_1553_),
    .I1(_1560_),
    .S(_1249_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5443_ (.I(_1051_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5444_ (.I(_1376_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5445_ (.A1(_1345_),
    .A2(_1171_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5446_ (.A1(_1282_),
    .A2(net172),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5447_ (.A1(_1564_),
    .A2(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5448_ (.I(_1053_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5449_ (.I(_1556_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5450_ (.I(_1084_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5451_ (.A1(_1282_),
    .A2(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5452_ (.A1(_1567_),
    .A2(_1568_),
    .B(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5453_ (.I(_1252_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5454_ (.I0(_1566_),
    .I1(_1571_),
    .S(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5455_ (.I(_0980_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5456_ (.I(_1574_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5457_ (.I(_1040_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5458_ (.I(_0963_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_1390_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5460_ (.I(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5461_ (.A1(_1577_),
    .A2(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5462_ (.A1(_1576_),
    .A2(_1568_),
    .B(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5463_ (.I(_1574_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5464_ (.I(_1310_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5465_ (.A1(_1583_),
    .A2(_1025_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5466_ (.A1(_1582_),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5467_ (.A1(_1575_),
    .A2(_1581_),
    .B(_1585_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5468_ (.A1(_1563_),
    .A2(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5469_ (.A1(_1563_),
    .A2(_1573_),
    .B(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5470_ (.A1(_1562_),
    .A2(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5471_ (.A1(_1546_),
    .A2(_1561_),
    .B(_1589_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5472_ (.A1(_1223_),
    .A2(_1226_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5473_ (.A1(net4),
    .A2(_1216_),
    .B(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5474_ (.A1(net24),
    .A2(_1221_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5475_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5476_ (.A1(_1225_),
    .A2(_1592_),
    .A3(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5477_ (.I(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5478_ (.I(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5479_ (.I(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5480_ (.I(_0608_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5481_ (.A1(_1229_),
    .A2(_1594_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5482_ (.I(_1600_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5483_ (.A1(_1225_),
    .A2(_1228_),
    .A3(_1594_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5484_ (.I(_1602_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5485_ (.A1(_1599_),
    .A2(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5486_ (.A1(_1599_),
    .A2(_1601_),
    .B(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5487_ (.A1(_1598_),
    .A2(_1605_),
    .B(_0607_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5488_ (.A1(_1239_),
    .A2(_1539_),
    .B1(_1544_),
    .B2(_1590_),
    .C(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5489_ (.A1(_0608_),
    .A2(_0607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5490_ (.I(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5491_ (.A1(_1210_),
    .A2(_0668_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5492_ (.I(_0779_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5493_ (.I(_0822_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5494_ (.A1(_0842_),
    .A2(_1194_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5495_ (.I(_0904_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5496_ (.A1(_0842_),
    .A2(_1194_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5497_ (.A1(_1613_),
    .A2(_1614_),
    .B(_1615_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5498_ (.A1(_1612_),
    .A2(_1616_),
    .B(_0823_),
    .C(_0780_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5499_ (.A1(_1611_),
    .A2(_1617_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5500_ (.I(_1108_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5501_ (.A1(_1178_),
    .A2(_1180_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5502_ (.A1(_1178_),
    .A2(_1180_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5503_ (.A1(_1619_),
    .A2(_1620_),
    .B(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5504_ (.A1(_1122_),
    .A2(_1172_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5505_ (.I(_1162_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5506_ (.A1(_1240_),
    .A2(_1052_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5507_ (.I(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5508_ (.A1(_1247_),
    .A2(_1577_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5509_ (.A1(_0989_),
    .A2(_1038_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5510_ (.A1(_1403_),
    .A2(_1023_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5511_ (.A1(net65),
    .A2(_0866_),
    .B(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5512_ (.A1(_0980_),
    .A2(_0990_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5513_ (.A1(net210),
    .A2(_1255_),
    .A3(_1630_),
    .B(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5514_ (.A1(_1247_),
    .A2(net180),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5515_ (.A1(_1627_),
    .A2(_1632_),
    .B(_1633_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5516_ (.A1(_1048_),
    .A2(_1052_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5517_ (.I(_1635_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5518_ (.A1(_1626_),
    .A2(_1634_),
    .B(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5519_ (.A1(_1122_),
    .A2(_1172_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5520_ (.A1(_1534_),
    .A2(_1569_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5521_ (.A1(_1086_),
    .A2(_1637_),
    .B(_1638_),
    .C(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _5522_ (.A1(_1165_),
    .A2(_1623_),
    .A3(_1624_),
    .A4(_1640_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5523_ (.A1(_1622_),
    .A2(_1641_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5524_ (.A1(_0823_),
    .A2(_0821_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5525_ (.A1(_0782_),
    .A2(net222),
    .A3(_0864_),
    .A4(_0907_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5526_ (.A1(_1642_),
    .A2(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5527_ (.A1(_1618_),
    .A2(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5528_ (.A1(_0639_),
    .A2(_1211_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5529_ (.A1(_0639_),
    .A2(_1211_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5530_ (.A1(_1647_),
    .A2(_0721_),
    .B(_1648_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5531_ (.A1(_1610_),
    .A2(_0724_),
    .A3(_1646_),
    .B(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5532_ (.A1(_1222_),
    .A2(_1236_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5533_ (.I(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5534_ (.A1(_1220_),
    .A2(_1230_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5535_ (.A1(_1222_),
    .A2(_1592_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5536_ (.A1(_1220_),
    .A2(_1654_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5537_ (.A1(_1652_),
    .A2(_1653_),
    .A3(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5538_ (.I(_1656_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5539_ (.I(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5540_ (.A1(_1609_),
    .A2(_1650_),
    .B(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5541_ (.A1(_1609_),
    .A2(_1650_),
    .B(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5542_ (.A1(_1234_),
    .A2(_1607_),
    .A3(_1660_),
    .ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5543_ (.I(_0557_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5544_ (.I(_0559_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5545_ (.A1(_1267_),
    .A2(_1661_),
    .B(_1662_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5546_ (.I(_0703_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5547_ (.I0(\reg_file.reg_storage[4][15] ),
    .I1(\reg_file.reg_storage[5][15] ),
    .I2(\reg_file.reg_storage[6][15] ),
    .I3(\reg_file.reg_storage[7][15] ),
    .S0(_0892_),
    .S1(_1664_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5548_ (.I(_0996_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5549_ (.I(_0652_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5550_ (.A1(_1667_),
    .A2(\reg_file.reg_storage[3][15] ),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5551_ (.A1(_0591_),
    .A2(\reg_file.reg_storage[2][15] ),
    .B(_1152_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5552_ (.A1(_1666_),
    .A2(_1445_),
    .B1(_1668_),
    .B2(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5553_ (.I0(\reg_file.reg_storage[12][15] ),
    .I1(\reg_file.reg_storage[13][15] ),
    .I2(\reg_file.reg_storage[14][15] ),
    .I3(\reg_file.reg_storage[15][15] ),
    .S0(_0892_),
    .S1(_0704_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5554_ (.I0(\reg_file.reg_storage[8][15] ),
    .I1(\reg_file.reg_storage[9][15] ),
    .I2(\reg_file.reg_storage[10][15] ),
    .I3(\reg_file.reg_storage[11][15] ),
    .S0(_0892_),
    .S1(_1664_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5555_ (.I0(_1665_),
    .I1(_1670_),
    .I2(_1671_),
    .I3(_1672_),
    .S0(_0900_),
    .S1(_0718_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5556_ (.A1(_0882_),
    .A2(_1663_),
    .B1(_1673_),
    .B2(_0902_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5557_ (.A1(_1452_),
    .A2(_1674_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5558_ (.A1(_1452_),
    .A2(net229),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5559_ (.A1(_1676_),
    .A2(_1675_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5560_ (.I(_1677_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5561_ (.I(_0537_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5562_ (.A1(_1679_),
    .A2(_0606_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5563_ (.A1(_0610_),
    .A2(_1213_),
    .B(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5564_ (.A1(_1220_),
    .A2(_1230_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5565_ (.I(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5566_ (.A1(_1678_),
    .A2(_1681_),
    .B(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5567_ (.A1(_1678_),
    .A2(_1681_),
    .B(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5568_ (.I(_1652_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5569_ (.I(_1545_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5570_ (.I(_1534_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5571_ (.A1(_1687_),
    .A2(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5572_ (.I(_1689_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5573_ (.I(_1305_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5574_ (.I(_1691_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5575_ (.I(_1692_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5576_ (.I(_1308_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5577_ (.I(_1694_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5578_ (.I(_1345_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_1696_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5580_ (.A1(_1697_),
    .A2(_1299_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5581_ (.A1(_1695_),
    .A2(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5582_ (.A1(_1693_),
    .A2(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5583_ (.I(_1051_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5584_ (.I(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5585_ (.I(_1578_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5586_ (.I(_1703_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5587_ (.A1(_1697_),
    .A2(_1279_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5588_ (.A1(_1704_),
    .A2(_1359_),
    .B(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5589_ (.I(_1282_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5590_ (.A1(_1707_),
    .A2(_1371_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5591_ (.I(_1708_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5592_ (.I(_1583_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5593_ (.A1(_1710_),
    .A2(_1327_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5594_ (.A1(_1709_),
    .A2(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5595_ (.I(_1694_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5596_ (.I0(_1706_),
    .I1(_1712_),
    .S(_1713_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5597_ (.I(_1696_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5598_ (.I(_1578_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5599_ (.A1(_1716_),
    .A2(_1341_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5600_ (.A1(_1715_),
    .A2(_1419_),
    .B(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5601_ (.A1(net81),
    .A2(_1258_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5602_ (.A1(_1311_),
    .A2(net168),
    .A3(_1432_),
    .B(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(_1703_),
    .A2(net176),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5604_ (.A1(_1715_),
    .A2(net211),
    .B(_1721_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5605_ (.I0(_1718_),
    .I1(_1722_),
    .S(_1694_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5606_ (.I(_1250_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5607_ (.I0(_1714_),
    .I1(_1723_),
    .S(_1724_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5608_ (.I(_1257_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5609_ (.I(_1508_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5610_ (.A1(_1726_),
    .A2(_1727_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5611_ (.I(_1578_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5612_ (.A1(_1311_),
    .A2(_1463_),
    .A3(_1468_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5613_ (.A1(_1469_),
    .A2(_1730_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5614_ (.A1(_1729_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5615_ (.A1(_1728_),
    .A2(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5616_ (.A1(net72),
    .A2(_1185_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5617_ (.A1(_1183_),
    .A2(_1477_),
    .A3(_1481_),
    .B(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5618_ (.A1(_1579_),
    .A2(_1453_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5619_ (.A1(_1715_),
    .A2(_1735_),
    .B(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5620_ (.I0(_1733_),
    .I1(_1737_),
    .S(_1694_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5621_ (.A1(_1716_),
    .A2(_1498_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5622_ (.A1(_1523_),
    .A2(_1527_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5623_ (.I(net77),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5624_ (.A1(_1741_),
    .A2(_0866_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5625_ (.A1(_1311_),
    .A2(_1740_),
    .B(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5626_ (.A1(_1726_),
    .A2(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5627_ (.A1(_1739_),
    .A2(_1744_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5628_ (.I(_1400_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5629_ (.I(net220),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5630_ (.A1(_1716_),
    .A2(_1747_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5631_ (.A1(_1715_),
    .A2(_1746_),
    .B(_1748_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5632_ (.I0(_1745_),
    .I1(_1749_),
    .S(_1572_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5633_ (.I(_1305_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5634_ (.I0(_1738_),
    .I1(_1750_),
    .S(_1751_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5635_ (.A1(_1243_),
    .A2(_1752_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5636_ (.I(_1244_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5637_ (.A1(_1702_),
    .A2(_1725_),
    .B(_1753_),
    .C(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5638_ (.A1(_1690_),
    .A2(_1700_),
    .B(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5639_ (.I(_1308_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5640_ (.I(_1577_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5641_ (.A1(_1053_),
    .A2(_1729_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5642_ (.A1(_1758_),
    .A2(_1568_),
    .B(_1759_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5643_ (.A1(_1757_),
    .A2(_1760_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5644_ (.I(_1026_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5645_ (.A1(_1040_),
    .A2(_1729_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5646_ (.A1(_1762_),
    .A2(_1763_),
    .B(_1487_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5647_ (.A1(_1761_),
    .A2(_1764_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5648_ (.A1(_1696_),
    .A2(net199),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5649_ (.A1(_1716_),
    .A2(_1175_),
    .B(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5650_ (.I(_1569_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5651_ (.A1(_1707_),
    .A2(_1122_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5652_ (.A1(_1557_),
    .A2(_1768_),
    .B(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5653_ (.I0(_1767_),
    .I1(_1770_),
    .S(_1572_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5654_ (.I0(_1765_),
    .I1(_1771_),
    .S(_1724_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5655_ (.A1(_1187_),
    .A2(_1556_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5656_ (.A1(_0842_),
    .A2(_1707_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(_1773_),
    .A2(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5658_ (.A1(net184),
    .A2(_1579_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5659_ (.A1(_1197_),
    .A2(_1697_),
    .B(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5660_ (.I0(_1775_),
    .I1(_1777_),
    .S(_1582_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(_0639_),
    .A2(_1579_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5662_ (.A1(_1205_),
    .A2(_1726_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(_1779_),
    .A2(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5664_ (.A1(_1679_),
    .A2(_1726_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5665_ (.A1(_1736_),
    .A2(_1782_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5666_ (.I(_1307_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5667_ (.I(_1784_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5668_ (.I0(_1781_),
    .I1(_1783_),
    .S(_1785_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5669_ (.I(_1563_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5670_ (.I0(_1778_),
    .I1(_1786_),
    .S(_1787_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5671_ (.I(_1240_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5672_ (.I0(_1772_),
    .I1(_1788_),
    .S(_1789_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5673_ (.I(_1536_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5674_ (.A1(_1236_),
    .A2(_1540_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5675_ (.I(_1792_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5676_ (.I(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5677_ (.A1(_1791_),
    .A2(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5678_ (.A1(_1225_),
    .A2(_1593_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5679_ (.A1(_1592_),
    .A2(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5680_ (.I(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5681_ (.I(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5682_ (.A1(_1229_),
    .A2(_1594_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5683_ (.I(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5684_ (.I(_1801_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5685_ (.I(_1596_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5686_ (.A1(_1802_),
    .A2(_1676_),
    .B(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5687_ (.I(net213),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(_1453_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5689_ (.A1(_1799_),
    .A2(_1676_),
    .B1(_1804_),
    .B2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5690_ (.A1(_1686_),
    .A2(_1756_),
    .B1(_1790_),
    .B2(_1795_),
    .C(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _5691_ (.I(_1677_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5692_ (.A1(_1609_),
    .A2(_1650_),
    .B(_1599_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5693_ (.A1(_1651_),
    .A2(_1653_),
    .A3(_1655_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5694_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5695_ (.I(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5696_ (.A1(_1809_),
    .A2(_1810_),
    .B(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5697_ (.A1(_1809_),
    .A2(_1810_),
    .B(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5698_ (.A1(_1685_),
    .A2(_1808_),
    .A3(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5699_ (.I(_1816_),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5700_ (.I(_1812_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5701_ (.I(_1817_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5702_ (.I(_0843_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5703_ (.A1(_1263_),
    .A2(_1661_),
    .B(_1662_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5704_ (.I(_1157_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5705_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(\reg_file.reg_storage[5][16] ),
    .I2(\reg_file.reg_storage[6][16] ),
    .I3(\reg_file.reg_storage[7][16] ),
    .S0(_0813_),
    .S1(_1821_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5706_ (.I(_1152_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5707_ (.I(\reg_file.reg_storage[1][16] ),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5708_ (.I(_0645_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5709_ (.A1(_1825_),
    .A2(\reg_file.reg_storage[3][16] ),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5710_ (.I(_0852_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5711_ (.A1(_1827_),
    .A2(\reg_file.reg_storage[2][16] ),
    .B(_1666_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5712_ (.A1(_1823_),
    .A2(_1824_),
    .B1(_1826_),
    .B2(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5713_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(\reg_file.reg_storage[13][16] ),
    .I2(\reg_file.reg_storage[14][16] ),
    .I3(\reg_file.reg_storage[15][16] ),
    .S0(_0587_),
    .S1(_1821_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5714_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(\reg_file.reg_storage[9][16] ),
    .I2(\reg_file.reg_storage[10][16] ),
    .I3(\reg_file.reg_storage[11][16] ),
    .S0(_0587_),
    .S1(_1821_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5715_ (.I(_0662_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5716_ (.I(_0775_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _5717_ (.I0(_1822_),
    .I1(_1829_),
    .I2(_1830_),
    .I3(_1831_),
    .S0(_1832_),
    .S1(_1833_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5718_ (.I(_0861_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5719_ (.A1(_1819_),
    .A2(_1820_),
    .B1(_1834_),
    .B2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5720_ (.A1(_1483_),
    .A2(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5721_ (.A1(_1483_),
    .A2(_1836_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5722_ (.A1(_1837_),
    .A2(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5723_ (.I(_1839_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5724_ (.A1(_1609_),
    .A2(_0670_),
    .A3(_0723_),
    .A4(_1678_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5725_ (.A1(_1622_),
    .A2(_1641_),
    .B(_1644_),
    .C(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5726_ (.I(_1618_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5727_ (.I(_1649_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5728_ (.A1(_0607_),
    .A2(_1675_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5729_ (.A1(_1599_),
    .A2(_1844_),
    .B(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5730_ (.A1(_1453_),
    .A2(_1805_),
    .B1(_1841_),
    .B2(_1843_),
    .C(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5731_ (.A1(_1842_),
    .A2(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5732_ (.A1(_1840_),
    .A2(_1848_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5733_ (.I(_1839_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5734_ (.A1(_1608_),
    .A2(_0669_),
    .A3(_0723_),
    .A4(_1677_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5735_ (.A1(_0781_),
    .A2(_1643_),
    .A3(_0863_),
    .A4(_0906_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5736_ (.A1(_1851_),
    .A2(_1852_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5737_ (.A1(_1187_),
    .A2(_0903_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5738_ (.A1(_0863_),
    .A2(_1854_),
    .B(_1195_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5739_ (.A1(_0824_),
    .A2(_1855_),
    .B(_1198_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5740_ (.A1(_0781_),
    .A2(_1856_),
    .B(_1201_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5741_ (.A1(_1205_),
    .A2(_0720_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5742_ (.A1(_0670_),
    .A2(_1858_),
    .B(_1212_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5743_ (.A1(_0610_),
    .A2(_1859_),
    .B(_1680_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(_1454_),
    .A2(_1805_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5745_ (.A1(_1678_),
    .A2(_1860_),
    .B(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5746_ (.A1(_1182_),
    .A2(_1853_),
    .B1(_1857_),
    .B2(net171),
    .C(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5747_ (.A1(_1850_),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5748_ (.A1(_0964_),
    .A2(_0935_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5749_ (.A1(_1003_),
    .A2(_1025_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5750_ (.A1(_1039_),
    .A2(_0990_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5751_ (.A1(_1628_),
    .A2(_1866_),
    .B(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5752_ (.A1(_1049_),
    .A2(_1047_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5753_ (.A1(_1050_),
    .A2(_1052_),
    .B1(_1865_),
    .B2(_1868_),
    .C(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5754_ (.A1(_1085_),
    .A2(_1110_),
    .A3(_1135_),
    .A4(_1162_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5755_ (.A1(_1171_),
    .A2(_1134_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5756_ (.A1(_1167_),
    .A2(_1084_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5757_ (.A1(_1171_),
    .A2(_1172_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5758_ (.A1(_1872_),
    .A2(_1873_),
    .B(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5759_ (.A1(_1175_),
    .A2(_1107_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5760_ (.A1(_1110_),
    .A2(_1875_),
    .B(_1876_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5761_ (.A1(_1179_),
    .A2(_1180_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5762_ (.A1(_1870_),
    .A2(_1871_),
    .B1(_1877_),
    .B2(_1624_),
    .C(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5763_ (.A1(_1852_),
    .A2(_1851_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5764_ (.A1(_1611_),
    .A2(_0780_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5765_ (.A1(_1193_),
    .A2(_0862_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5766_ (.A1(_1193_),
    .A2(_1194_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5767_ (.A1(_1882_),
    .A2(_1188_),
    .B(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5768_ (.A1(_1197_),
    .A2(_0820_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5769_ (.A1(_1643_),
    .A2(_1884_),
    .B(_1885_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5770_ (.A1(_1200_),
    .A2(_0778_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5771_ (.A1(_1881_),
    .A2(_1886_),
    .B(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5772_ (.A1(_0609_),
    .A2(_1610_),
    .A3(_0724_),
    .A4(_1809_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5773_ (.A1(_1210_),
    .A2(_1211_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5774_ (.A1(_1610_),
    .A2(_1206_),
    .B(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5775_ (.A1(_1679_),
    .A2(_0606_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5776_ (.A1(_1608_),
    .A2(_1891_),
    .B(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5777_ (.A1(_1454_),
    .A2(_1805_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5778_ (.A1(_1809_),
    .A2(_1893_),
    .B(_1894_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5779_ (.A1(_1879_),
    .A2(_1880_),
    .B1(_1888_),
    .B2(_1889_),
    .C(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5780_ (.I(_1231_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5781_ (.I(_1897_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5782_ (.A1(_1840_),
    .A2(_1896_),
    .B(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _5783_ (.A1(_1535_),
    .A2(_1237_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5784_ (.A1(_1280_),
    .A2(_1300_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5785_ (.A1(_1360_),
    .A2(_1372_),
    .B(_1307_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5786_ (.A1(_1784_),
    .A2(_1901_),
    .B(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5787_ (.I(_1039_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5788_ (.I0(_1436_),
    .I1(_1343_),
    .S(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5789_ (.A1(_1248_),
    .A2(_1905_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5790_ (.A1(_1304_),
    .A2(_1903_),
    .B(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5791_ (.I0(_1485_),
    .I1(_1509_),
    .S(_1904_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5792_ (.I0(_1530_),
    .I1(_1402_),
    .S(_1904_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5793_ (.I0(_1908_),
    .I1(_1909_),
    .S(net206),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5794_ (.A1(_1440_),
    .A2(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5795_ (.A1(_1241_),
    .A2(_1907_),
    .B(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _5796_ (.I(_1797_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5797_ (.I(_1838_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5798_ (.A1(_1801_),
    .A2(_1914_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5799_ (.A1(_1228_),
    .A2(_1796_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5800_ (.I(_1916_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5801_ (.A1(_1913_),
    .A2(_1914_),
    .B(_1915_),
    .C(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5802_ (.I(_1792_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5803_ (.A1(_1248_),
    .A2(_1784_),
    .A3(_1584_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5804_ (.A1(_1557_),
    .A2(_1454_),
    .B(_1484_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5805_ (.I0(_1555_),
    .I1(_1921_),
    .S(_1785_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5806_ (.I(_1784_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5807_ (.I0(_1549_),
    .I1(_1559_),
    .S(_1923_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5808_ (.I0(_1922_),
    .I1(_1924_),
    .S(_1691_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5809_ (.I0(_1581_),
    .I1(_1571_),
    .S(_1923_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5810_ (.I0(_1552_),
    .I1(_1566_),
    .S(_1486_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5811_ (.I(_1376_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5812_ (.I0(_1926_),
    .I1(_1927_),
    .S(_1928_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5813_ (.I0(_1925_),
    .I1(_1929_),
    .S(_1545_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(_1244_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5815_ (.A1(_1245_),
    .A2(_1920_),
    .B1(_1930_),
    .B2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5816_ (.A1(_1919_),
    .A2(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5817_ (.A1(_1900_),
    .A2(_1912_),
    .B1(_1918_),
    .B2(_1837_),
    .C(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5818_ (.A1(_1818_),
    .A2(_1849_),
    .B1(_1864_),
    .B2(_1899_),
    .C(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5819_ (.I(net165),
    .ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5820_ (.A1(_0690_),
    .A2(_0558_),
    .B(_0560_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5821_ (.I0(\reg_file.reg_storage[4][17] ),
    .I1(\reg_file.reg_storage[5][17] ),
    .I2(\reg_file.reg_storage[6][17] ),
    .I3(\reg_file.reg_storage[7][17] ),
    .S0(_0596_),
    .S1(_0597_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5822_ (.I(\reg_file.reg_storage[1][17] ),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5823_ (.A1(_0587_),
    .A2(\reg_file.reg_storage[3][17] ),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5824_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][17] ),
    .B(_0770_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5825_ (.A1(_0584_),
    .A2(_1938_),
    .B1(_1939_),
    .B2(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _5826_ (.I(_0574_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5827_ (.I(_0763_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5828_ (.I0(\reg_file.reg_storage[12][17] ),
    .I1(\reg_file.reg_storage[13][17] ),
    .I2(\reg_file.reg_storage[14][17] ),
    .I3(\reg_file.reg_storage[15][17] ),
    .S0(_1942_),
    .S1(_1943_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5829_ (.I0(\reg_file.reg_storage[8][17] ),
    .I1(\reg_file.reg_storage[9][17] ),
    .I2(\reg_file.reg_storage[10][17] ),
    .I3(\reg_file.reg_storage[11][17] ),
    .S0(_1942_),
    .S1(_0597_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5830_ (.I0(_1937_),
    .I1(_1941_),
    .I2(_1944_),
    .I3(_1945_),
    .S0(_0602_),
    .S1(_0604_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5831_ (.A1(_0549_),
    .A2(_1936_),
    .B1(_1946_),
    .B2(_0571_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5832_ (.A1(_1470_),
    .A2(_1947_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5833_ (.I(_1948_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5834_ (.I(_1949_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5835_ (.A1(_1840_),
    .A2(_1848_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5836_ (.A1(_1914_),
    .A2(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5837_ (.I(_1657_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5838_ (.A1(_1950_),
    .A2(_1952_),
    .B(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5839_ (.A1(_1950_),
    .A2(_1952_),
    .B(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5840_ (.A1(_1735_),
    .A2(_1836_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5841_ (.A1(_1850_),
    .A2(_1863_),
    .B(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5842_ (.A1(_1950_),
    .A2(_1957_),
    .B(_1232_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5843_ (.A1(_1950_),
    .A2(_1957_),
    .B(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5844_ (.I(_1913_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5845_ (.A1(_1731_),
    .A2(_1947_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(_1731_),
    .A2(_1947_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5847_ (.I(_1800_),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5848_ (.I(_1963_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5849_ (.A1(_1964_),
    .A2(_1961_),
    .B(_1598_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5850_ (.A1(_1960_),
    .A2(_1961_),
    .B1(_1962_),
    .B2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5851_ (.I(_1793_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5852_ (.A1(_1486_),
    .A2(_1762_),
    .A3(_1763_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5853_ (.A1(_1251_),
    .A2(_1968_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5854_ (.I(_1242_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5855_ (.I(_1970_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5856_ (.I0(_1760_),
    .I1(_1770_),
    .S(_1785_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5857_ (.I(_1574_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5858_ (.I0(_1767_),
    .I1(_1775_),
    .S(_1973_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5859_ (.A1(_1377_),
    .A2(_1974_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5860_ (.A1(_1306_),
    .A2(_1972_),
    .B(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5861_ (.I(_1241_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5862_ (.I(_1977_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5863_ (.A1(_1568_),
    .A2(_1735_),
    .B(_1732_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5864_ (.I0(_1783_),
    .I1(_1979_),
    .S(_1923_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5865_ (.I0(_1777_),
    .I1(_1781_),
    .S(_1582_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5866_ (.I0(_1980_),
    .I1(_1981_),
    .S(_1751_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5867_ (.A1(_1978_),
    .A2(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5868_ (.A1(_1971_),
    .A2(_1976_),
    .B(_1983_),
    .C(_1537_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5869_ (.A1(_1246_),
    .A2(_1969_),
    .B(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5870_ (.I(_1441_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5871_ (.I(_1986_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5872_ (.I(_1376_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5873_ (.I(_1988_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5874_ (.I(_1989_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5875_ (.A1(_1309_),
    .A2(_1698_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5876_ (.A1(_1757_),
    .A2(_1706_),
    .B(_1991_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5877_ (.I(_1249_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5878_ (.I(_1582_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5879_ (.I0(_1712_),
    .I1(_1718_),
    .S(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5880_ (.A1(_1993_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5881_ (.A1(_1990_),
    .A2(_1992_),
    .B(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5882_ (.I(_1242_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5883_ (.I(_1998_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5884_ (.I0(_1733_),
    .I1(_1745_),
    .S(_1572_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5885_ (.I0(_1749_),
    .I1(_1722_),
    .S(_1373_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5886_ (.A1(_1692_),
    .A2(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5887_ (.A1(_1993_),
    .A2(_2000_),
    .B(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5888_ (.A1(_1999_),
    .A2(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5889_ (.A1(_1987_),
    .A2(_1997_),
    .B(_2004_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _5890_ (.A1(_1244_),
    .A2(_1652_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5891_ (.I(_2006_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5892_ (.A1(_1967_),
    .A2(_1985_),
    .B1(_2005_),
    .B2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5893_ (.A1(_1955_),
    .A2(_1959_),
    .A3(_1966_),
    .A4(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5894_ (.I(_2009_),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5895_ (.A1(_1412_),
    .A2(_1661_),
    .B(_1662_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5896_ (.I(_1125_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5897_ (.I0(\reg_file.reg_storage[4][18] ),
    .I1(\reg_file.reg_storage[5][18] ),
    .I2(\reg_file.reg_storage[6][18] ),
    .I3(\reg_file.reg_storage[7][18] ),
    .S0(_0767_),
    .S1(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5898_ (.I(_0755_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5899_ (.A1(_2013_),
    .A2(\reg_file.reg_storage[3][18] ),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5900_ (.A1(_0895_),
    .A2(\reg_file.reg_storage[2][18] ),
    .B(_0766_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5901_ (.A1(_0890_),
    .A2(_1500_),
    .B1(_2014_),
    .B2(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5902_ (.I(_1125_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5903_ (.I0(\reg_file.reg_storage[12][18] ),
    .I1(\reg_file.reg_storage[13][18] ),
    .I2(\reg_file.reg_storage[14][18] ),
    .I3(\reg_file.reg_storage[15][18] ),
    .S0(_0887_),
    .S1(_2017_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5904_ (.I0(\reg_file.reg_storage[8][18] ),
    .I1(\reg_file.reg_storage[9][18] ),
    .I2(\reg_file.reg_storage[10][18] ),
    .I3(\reg_file.reg_storage[11][18] ),
    .S0(_0887_),
    .S1(_2017_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5905_ (.I(_0859_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5906_ (.I0(_2012_),
    .I1(_2016_),
    .I2(_2018_),
    .I3(_2019_),
    .S0(_0900_),
    .S1(_2020_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5907_ (.A1(_0882_),
    .A2(_2010_),
    .B1(_2021_),
    .B2(_0902_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5908_ (.A1(_1507_),
    .A2(_2022_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5909_ (.A1(_1508_),
    .A2(_2022_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5910_ (.A1(_2024_),
    .A2(_2023_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5911_ (.I(net195),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5912_ (.I(_2026_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5913_ (.A1(_1914_),
    .A2(_1961_),
    .B(_1962_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5914_ (.A1(_1840_),
    .A2(_1848_),
    .A3(_1949_),
    .B(_2028_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5915_ (.A1(_2027_),
    .A2(_2029_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5916_ (.A1(_2027_),
    .A2(_2029_),
    .B(_1813_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5917_ (.A1(_1470_),
    .A2(_1947_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5918_ (.A1(_1949_),
    .A2(_1957_),
    .B(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5919_ (.A1(_2027_),
    .A2(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5920_ (.I(_1683_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5921_ (.A1(_2027_),
    .A2(_2033_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5922_ (.A1(_2035_),
    .A2(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5923_ (.I(_1535_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5924_ (.I(_2038_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5925_ (.A1(_1729_),
    .A2(_1508_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5926_ (.A1(_1557_),
    .A2(_1470_),
    .B(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5927_ (.I0(_1921_),
    .I1(_2041_),
    .S(_1973_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5928_ (.I0(_1560_),
    .I1(_2042_),
    .S(_1989_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5929_ (.I0(_1553_),
    .I1(_1573_),
    .S(_1751_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5930_ (.I0(_2043_),
    .I1(_2044_),
    .S(_1562_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5931_ (.I(_1688_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5932_ (.A1(_1970_),
    .A2(_1251_),
    .A3(_1586_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5933_ (.A1(_2046_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5934_ (.A1(_2039_),
    .A2(_2045_),
    .B(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5935_ (.I(_1562_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5936_ (.I(_1304_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5937_ (.I(_2051_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5938_ (.I0(_1531_),
    .I1(_1437_),
    .S(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5939_ (.I(_1687_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5940_ (.I(_1928_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5941_ (.A1(_2055_),
    .A2(_1301_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5942_ (.A1(_1251_),
    .A2(_1375_),
    .B(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5943_ (.A1(_2054_),
    .A2(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5944_ (.A1(_2050_),
    .A2(_2053_),
    .B(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5945_ (.I(_1595_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5946_ (.I(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5947_ (.I(_1600_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5948_ (.I(_2024_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5949_ (.I(_1602_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5950_ (.A1(_2064_),
    .A2(_2063_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5951_ (.A1(_2062_),
    .A2(_2063_),
    .B(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5952_ (.A1(_2061_),
    .A2(_2066_),
    .B(_2023_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5953_ (.A1(_1967_),
    .A2(_2049_),
    .B1(_2059_),
    .B2(_2007_),
    .C(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5954_ (.A1(_2030_),
    .A2(_2031_),
    .B1(_2034_),
    .B2(_2037_),
    .C(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5955_ (.I(_2069_),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5956_ (.I(_0745_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5957_ (.A1(_0496_),
    .A2(_1661_),
    .B(_1662_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5958_ (.I(_0702_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5959_ (.I(_1150_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5960_ (.I0(\reg_file.reg_storage[4][19] ),
    .I1(\reg_file.reg_storage[5][19] ),
    .I2(\reg_file.reg_storage[6][19] ),
    .I3(\reg_file.reg_storage[7][19] ),
    .S0(_2072_),
    .S1(_2073_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5961_ (.A1(_0756_),
    .A2(\reg_file.reg_storage[3][19] ),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5962_ (.I(_0654_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5963_ (.A1(_2076_),
    .A2(\reg_file.reg_storage[2][19] ),
    .B(_1666_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5964_ (.A1(_1823_),
    .A2(_1490_),
    .B1(_2075_),
    .B2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5965_ (.I(_1157_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5966_ (.I0(\reg_file.reg_storage[12][19] ),
    .I1(\reg_file.reg_storage[13][19] ),
    .I2(\reg_file.reg_storage[14][19] ),
    .I3(\reg_file.reg_storage[15][19] ),
    .S0(_0711_),
    .S1(_2079_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5967_ (.I0(\reg_file.reg_storage[8][19] ),
    .I1(\reg_file.reg_storage[9][19] ),
    .I2(\reg_file.reg_storage[10][19] ),
    .I3(\reg_file.reg_storage[11][19] ),
    .S0(_0711_),
    .S1(_2079_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5968_ (.I(_0717_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _5969_ (.I0(_2074_),
    .I1(_2078_),
    .I2(_2080_),
    .I3(_2081_),
    .S0(_2082_),
    .S1(_1833_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5970_ (.I(_0777_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5971_ (.A1(_2070_),
    .A2(_2071_),
    .B1(_2083_),
    .B2(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5972_ (.A1(_1497_),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5973_ (.A1(_1497_),
    .A2(_2085_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5974_ (.A1(_2086_),
    .A2(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5975_ (.I(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5976_ (.A1(_1727_),
    .A2(_2022_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5977_ (.A1(_2026_),
    .A2(_2033_),
    .B(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5978_ (.A1(_2089_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5979_ (.A1(_2089_),
    .A2(_2091_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5980_ (.A1(_2035_),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5981_ (.A1(_2063_),
    .A2(_2030_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5982_ (.I(_1657_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5983_ (.A1(_2089_),
    .A2(_2095_),
    .B(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5984_ (.A1(_2089_),
    .A2(_2095_),
    .B(_2097_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5985_ (.I(_2038_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5986_ (.I(_2052_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5987_ (.A1(_1702_),
    .A2(_2100_),
    .A3(_1765_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5988_ (.I0(_1771_),
    .I1(_1778_),
    .S(_1377_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5989_ (.I(_1441_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5990_ (.A1(_1728_),
    .A2(_1739_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5991_ (.I0(_1979_),
    .I1(_2104_),
    .S(_1994_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5992_ (.A1(_1250_),
    .A2(_1786_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5993_ (.A1(_1692_),
    .A2(_2105_),
    .B(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5994_ (.A1(_2103_),
    .A2(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5995_ (.I(_1688_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5996_ (.A1(_1999_),
    .A2(_2102_),
    .B(_2108_),
    .C(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5997_ (.A1(_2099_),
    .A2(_2101_),
    .B(_2110_),
    .C(_1967_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5998_ (.I(_2086_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5999_ (.I(_2087_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6000_ (.A1(_1802_),
    .A2(_2112_),
    .B(_1803_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6001_ (.I(_1977_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6002_ (.I0(_1699_),
    .I1(_1714_),
    .S(_1724_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6003_ (.I0(_1750_),
    .I1(_1723_),
    .S(_2051_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6004_ (.A1(_1687_),
    .A2(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6005_ (.A1(_2115_),
    .A2(_2116_),
    .B(_2118_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6006_ (.A1(_1799_),
    .A2(_2112_),
    .B1(_2113_),
    .B2(_2114_),
    .C1(_2119_),
    .C2(_2007_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6007_ (.A1(_2111_),
    .A2(_2120_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6008_ (.A1(_2092_),
    .A2(_2094_),
    .B(_2098_),
    .C(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6009_ (.I(_2122_),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6010_ (.I(_0769_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6011_ (.I(_0910_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6012_ (.A1(_0746_),
    .A2(_0910_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6013_ (.I(_2125_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6014_ (.A1(_2123_),
    .A2(_2124_),
    .B(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6015_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(\reg_file.reg_storage[5][20] ),
    .I2(\reg_file.reg_storage[6][20] ),
    .I3(\reg_file.reg_storage[7][20] ),
    .S0(_1942_),
    .S1(_1943_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6016_ (.I(\reg_file.reg_storage[1][20] ),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6017_ (.I(_0886_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6018_ (.A1(_2130_),
    .A2(\reg_file.reg_storage[3][20] ),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6019_ (.A1(_0769_),
    .A2(\reg_file.reg_storage[2][20] ),
    .B(_0770_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6020_ (.A1(_0584_),
    .A2(_2129_),
    .B1(_2131_),
    .B2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6021_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(\reg_file.reg_storage[13][20] ),
    .I2(\reg_file.reg_storage[14][20] ),
    .I3(\reg_file.reg_storage[15][20] ),
    .S0(net185),
    .S1(_1943_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6022_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(\reg_file.reg_storage[9][20] ),
    .I2(\reg_file.reg_storage[10][20] ),
    .I3(\reg_file.reg_storage[11][20] ),
    .S0(_1942_),
    .S1(_1943_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6023_ (.I0(_2128_),
    .I1(_2133_),
    .I2(_2134_),
    .I3(_2135_),
    .S0(_0602_),
    .S1(_0604_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6024_ (.A1(_0745_),
    .A2(_2127_),
    .B1(_2136_),
    .B2(_0777_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6025_ (.A1(_2137_),
    .A2(_1529_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6026_ (.A1(_1529_),
    .A2(_2137_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6027_ (.I(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6028_ (.A1(net193),
    .A2(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6029_ (.I(_2085_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6030_ (.A1(_1498_),
    .A2(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6031_ (.A1(_2088_),
    .A2(_2091_),
    .B(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6032_ (.A1(_2141_),
    .A2(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6033_ (.A1(_2141_),
    .A2(_2144_),
    .B(_1898_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6034_ (.A1(_1839_),
    .A2(_1949_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6035_ (.A1(_2087_),
    .A2(_2112_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6036_ (.A1(_2026_),
    .A2(_2147_),
    .A3(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6037_ (.I(_2063_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6038_ (.A1(_2150_),
    .A2(_2028_),
    .B(_2087_),
    .C(_2023_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6039_ (.A1(_2112_),
    .A2(_2151_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6040_ (.I(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6041_ (.A1(_1848_),
    .A2(_2149_),
    .B(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6042_ (.A1(_2141_),
    .A2(_2154_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6043_ (.A1(_2141_),
    .A2(_2154_),
    .B(_1817_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6044_ (.A1(_2155_),
    .A2(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6045_ (.I(_1306_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6046_ (.A1(_2158_),
    .A2(_1903_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6047_ (.I(_2051_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6048_ (.I0(_1909_),
    .I1(_1905_),
    .S(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6049_ (.A1(_2115_),
    .A2(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6050_ (.A1(_1971_),
    .A2(_2159_),
    .B(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6051_ (.A1(_1963_),
    .A2(_2140_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6052_ (.A1(_1913_),
    .A2(_2140_),
    .B(_2164_),
    .C(_1917_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(_1695_),
    .A2(_1584_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6054_ (.I(_1988_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _6055_ (.I0(_2166_),
    .I1(_1926_),
    .S(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6056_ (.I(_1441_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6057_ (.I0(_1924_),
    .I1(_1927_),
    .S(_1691_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6058_ (.I(_2170_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6059_ (.I0(_1498_),
    .I1(net178),
    .S(_1703_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6060_ (.I0(_2041_),
    .I1(_2172_),
    .S(_1785_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6061_ (.I0(_1922_),
    .I1(_2173_),
    .S(_1928_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6062_ (.A1(_1442_),
    .A2(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6063_ (.I(_1535_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6064_ (.A1(_2169_),
    .A2(_2171_),
    .B(_2175_),
    .C(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6065_ (.A1(_1245_),
    .A2(_2168_),
    .B(_2177_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6066_ (.A1(_1794_),
    .A2(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6067_ (.A1(_1900_),
    .A2(_2163_),
    .B1(_2165_),
    .B2(net194),
    .C(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6068_ (.A1(_2145_),
    .A2(_2146_),
    .B(_2157_),
    .C(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6069_ (.I(net164),
    .ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6070_ (.I(_0649_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6071_ (.A1(_2182_),
    .A2(_2124_),
    .B(_2125_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6072_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(\reg_file.reg_storage[5][21] ),
    .I2(\reg_file.reg_storage[6][21] ),
    .I3(\reg_file.reg_storage[7][21] ),
    .S0(_0658_),
    .S1(_1103_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6073_ (.A1(_0702_),
    .A2(\reg_file.reg_storage[3][21] ),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6074_ (.A1(_0852_),
    .A2(\reg_file.reg_storage[2][21] ),
    .B(_0583_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6075_ (.A1(_0593_),
    .A2(_1511_),
    .B1(_2185_),
    .B2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6076_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(\reg_file.reg_storage[13][21] ),
    .I2(\reg_file.reg_storage[14][21] ),
    .I3(\reg_file.reg_storage[15][21] ),
    .S0(_0846_),
    .S1(_0848_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6077_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(\reg_file.reg_storage[9][21] ),
    .I2(\reg_file.reg_storage[10][21] ),
    .I3(\reg_file.reg_storage[11][21] ),
    .S0(_0846_),
    .S1(_1103_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6078_ (.I0(_2184_),
    .I1(_2187_),
    .I2(_2188_),
    .I3(_2189_),
    .S0(_0858_),
    .S1(_0664_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6079_ (.A1(_0641_),
    .A2(_2183_),
    .B1(_2190_),
    .B2(_0667_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6080_ (.A1(_1518_),
    .A2(_2191_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6081_ (.I(_2192_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6082_ (.A1(_1743_),
    .A2(_2137_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6083_ (.A1(_2145_),
    .A2(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6084_ (.A1(_2193_),
    .A2(_2195_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6085_ (.A1(_2193_),
    .A2(_2195_),
    .B(_1898_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6086_ (.A1(_2140_),
    .A2(_2155_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6087_ (.A1(_2193_),
    .A2(_2198_),
    .B(_1817_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6088_ (.A1(_2193_),
    .A2(_2198_),
    .B(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6089_ (.I(_1998_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6090_ (.A1(_1744_),
    .A2(_1748_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6091_ (.I0(_2104_),
    .I1(_2202_),
    .S(_1923_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6092_ (.I0(_1980_),
    .I1(_2203_),
    .S(_1988_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6093_ (.A1(_2201_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6094_ (.I0(_1981_),
    .I1(_1974_),
    .S(_1691_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6095_ (.A1(_1546_),
    .A2(_2206_),
    .B(_1931_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6096_ (.A1(_1305_),
    .A2(_1968_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6097_ (.A1(_1751_),
    .A2(_1972_),
    .B(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6098_ (.A1(_2103_),
    .A2(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6099_ (.A1(_2205_),
    .A2(_2207_),
    .B1(_2210_),
    .B2(_1754_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6100_ (.A1(_1989_),
    .A2(_1992_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6101_ (.I0(_1995_),
    .I1(_2001_),
    .S(_1989_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6102_ (.A1(_1978_),
    .A2(_2213_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6103_ (.A1(_1303_),
    .A2(_2212_),
    .B(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6104_ (.I(_1797_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6105_ (.A1(_1747_),
    .A2(_2191_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6106_ (.A1(_1963_),
    .A2(_2217_),
    .B(_1597_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6107_ (.A1(_1747_),
    .A2(_2191_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6108_ (.A1(_2216_),
    .A2(_2217_),
    .B1(_2218_),
    .B2(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6109_ (.A1(_1541_),
    .A2(_2211_),
    .B1(_2215_),
    .B2(_1900_),
    .C(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6110_ (.A1(_2196_),
    .A2(_2197_),
    .B(_2200_),
    .C(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6111_ (.I(net162),
    .ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6112_ (.I(_0717_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6113_ (.A1(_2223_),
    .A2(_2124_),
    .B(_2126_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6114_ (.I(_0762_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6115_ (.I(_0993_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6116_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(\reg_file.reg_storage[5][22] ),
    .I2(\reg_file.reg_storage[6][22] ),
    .I3(\reg_file.reg_storage[7][22] ),
    .S0(_2225_),
    .S1(_2226_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6117_ (.A1(_1825_),
    .A2(\reg_file.reg_storage[3][22] ),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6118_ (.A1(_1827_),
    .A2(\reg_file.reg_storage[2][22] ),
    .B(_0706_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6119_ (.A1(_2182_),
    .A2(_1392_),
    .B1(_2228_),
    .B2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6120_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(\reg_file.reg_storage[13][22] ),
    .I2(\reg_file.reg_storage[14][22] ),
    .I3(\reg_file.reg_storage[15][22] ),
    .S0(_2225_),
    .S1(_2226_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6121_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(\reg_file.reg_storage[9][22] ),
    .I2(\reg_file.reg_storage[10][22] ),
    .I3(\reg_file.reg_storage[11][22] ),
    .S0(_2225_),
    .S1(_2226_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6122_ (.I0(_2227_),
    .I1(_2230_),
    .I2(_2231_),
    .I3(_2232_),
    .S0(_1832_),
    .S1(_2020_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6123_ (.A1(_1819_),
    .A2(_2224_),
    .B1(_2233_),
    .B2(_1835_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _6124_ (.A1(_1399_),
    .A2(_2234_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6125_ (.A1(_1400_),
    .A2(_2234_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6126_ (.I(_2236_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6127_ (.A1(_2235_),
    .A2(_2237_),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6128_ (.A1(_2138_),
    .A2(_2139_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6129_ (.A1(_2239_),
    .A2(_2192_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6130_ (.A1(_2139_),
    .A2(_2217_),
    .B(_2219_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6131_ (.I(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6132_ (.A1(_2154_),
    .A2(_2240_),
    .B(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6133_ (.A1(_2238_),
    .A2(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6134_ (.I(_2238_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6135_ (.A1(_2245_),
    .A2(_2243_),
    .B(_1812_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6136_ (.A1(_2239_),
    .A2(_2192_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6137_ (.A1(_1743_),
    .A2(_2137_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6138_ (.I(_0745_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6139_ (.I(_0777_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6140_ (.A1(_2249_),
    .A2(_2183_),
    .B1(net203),
    .B2(_2250_),
    .C(net219),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6141_ (.A1(_2192_),
    .A2(_2248_),
    .B(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6142_ (.A1(_2144_),
    .A2(_2247_),
    .B(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6143_ (.A1(_2238_),
    .A2(_2253_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6144_ (.A1(_2245_),
    .A2(_2253_),
    .B(_1682_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6145_ (.A1(_1701_),
    .A2(_1561_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6146_ (.I0(_1747_),
    .I1(_1400_),
    .S(_1703_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6147_ (.I0(_2172_),
    .I1(_2257_),
    .S(_1973_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6148_ (.I0(_2042_),
    .I1(_2258_),
    .S(_1928_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6149_ (.A1(_1442_),
    .A2(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6150_ (.A1(_1536_),
    .A2(_2256_),
    .A3(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6151_ (.A1(_1970_),
    .A2(_1931_),
    .A3(_1588_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6152_ (.A1(_2261_),
    .A2(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6153_ (.I(_1242_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6154_ (.A1(_2264_),
    .A2(_1439_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6155_ (.A1(_1986_),
    .A2(_1302_),
    .B(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6156_ (.A1(_1602_),
    .A2(_2237_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6157_ (.A1(_1600_),
    .A2(_2237_),
    .B(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6158_ (.A1(_2060_),
    .A2(_2268_),
    .B(_2235_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6159_ (.A1(_1919_),
    .A2(_2263_),
    .B1(_2266_),
    .B2(_2006_),
    .C(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6160_ (.A1(_2244_),
    .A2(_2246_),
    .B1(_2254_),
    .B2(_2255_),
    .C(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6161_ (.I(_2271_),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6162_ (.I(_2125_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6163_ (.A1(_0944_),
    .A2(_2124_),
    .B(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6164_ (.I0(\reg_file.reg_storage[4][23] ),
    .I1(\reg_file.reg_storage[5][23] ),
    .I2(\reg_file.reg_storage[6][23] ),
    .I3(\reg_file.reg_storage[7][23] ),
    .S0(_2225_),
    .S1(_2226_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6165_ (.A1(_1825_),
    .A2(\reg_file.reg_storage[3][23] ),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6166_ (.A1(_1827_),
    .A2(\reg_file.reg_storage[2][23] ),
    .B(_0706_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6167_ (.A1(_2182_),
    .A2(_1380_),
    .B1(_2275_),
    .B2(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6168_ (.I0(\reg_file.reg_storage[12][23] ),
    .I1(\reg_file.reg_storage[13][23] ),
    .I2(\reg_file.reg_storage[14][23] ),
    .I3(\reg_file.reg_storage[15][23] ),
    .S0(_2130_),
    .S1(_2011_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6169_ (.I0(\reg_file.reg_storage[8][23] ),
    .I1(\reg_file.reg_storage[9][23] ),
    .I2(\reg_file.reg_storage[10][23] ),
    .I3(\reg_file.reg_storage[11][23] ),
    .S0(_2130_),
    .S1(_2011_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6170_ (.I0(_2274_),
    .I1(_2277_),
    .I2(_2278_),
    .I3(_2279_),
    .S0(_1832_),
    .S1(_2020_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6171_ (.A1(_1819_),
    .A2(_2273_),
    .B1(_2280_),
    .B2(_1835_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _6172_ (.A1(_1388_),
    .A2(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6173_ (.A1(net179),
    .A2(net174),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6174_ (.A1(_2283_),
    .A2(_2282_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6175_ (.I(_2284_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6176_ (.I(_2237_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6177_ (.A1(_2245_),
    .A2(_2243_),
    .B(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6178_ (.A1(_2285_),
    .A2(_2287_),
    .B(_1658_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6179_ (.A1(_2285_),
    .A2(_2287_),
    .B(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6180_ (.I(_1931_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6181_ (.A1(_1710_),
    .A2(_1746_),
    .B(_1721_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6182_ (.I0(_2202_),
    .I1(_2291_),
    .S(_1994_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6183_ (.I0(_2105_),
    .I1(_2292_),
    .S(_2055_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6184_ (.I0(_1788_),
    .I1(_2293_),
    .S(_1443_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6185_ (.A1(_1546_),
    .A2(_1772_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6186_ (.A1(_2290_),
    .A2(_2295_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6187_ (.A1(_2290_),
    .A2(_2294_),
    .B(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6188_ (.A1(_2050_),
    .A2(_1700_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6189_ (.A1(_2050_),
    .A2(_1725_),
    .B(_2298_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6190_ (.A1(_1802_),
    .A2(net190),
    .B(_1803_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6191_ (.I(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6192_ (.I(_1798_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6193_ (.A1(_2302_),
    .A2(net190),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6194_ (.A1(_2282_),
    .A2(_2301_),
    .B(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6195_ (.A1(_1967_),
    .A2(_2297_),
    .B1(_2299_),
    .B2(_2007_),
    .C(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6196_ (.A1(_1746_),
    .A2(_2234_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6197_ (.A1(_2245_),
    .A2(_2253_),
    .B(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6198_ (.I(_1897_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6199_ (.A1(_2285_),
    .A2(_2307_),
    .B(_2308_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6200_ (.A1(_2285_),
    .A2(_2307_),
    .B(_2309_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6201_ (.A1(_2289_),
    .A2(_2305_),
    .A3(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6202_ (.I(_2311_),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6203_ (.I(_2126_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6204_ (.A1(net17),
    .A2(_0810_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6205_ (.A1(_2312_),
    .A2(_2313_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6206_ (.I(_0652_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6207_ (.I(_1150_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6208_ (.I0(\reg_file.reg_storage[4][24] ),
    .I1(\reg_file.reg_storage[5][24] ),
    .I2(\reg_file.reg_storage[6][24] ),
    .I3(\reg_file.reg_storage[7][24] ),
    .S0(_2315_),
    .S1(_2316_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6209_ (.I(_0766_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6210_ (.I(\reg_file.reg_storage[1][24] ),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6211_ (.I(_2130_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6212_ (.A1(_2320_),
    .A2(\reg_file.reg_storage[3][24] ),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6213_ (.I(_0996_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6214_ (.A1(_2123_),
    .A2(\reg_file.reg_storage[2][24] ),
    .B(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6215_ (.A1(_2318_),
    .A2(_2319_),
    .B1(_2321_),
    .B2(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6216_ (.I(_1150_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6217_ (.I0(\reg_file.reg_storage[12][24] ),
    .I1(\reg_file.reg_storage[13][24] ),
    .I2(\reg_file.reg_storage[14][24] ),
    .I3(\reg_file.reg_storage[15][24] ),
    .S0(_2315_),
    .S1(_2325_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6218_ (.I0(\reg_file.reg_storage[8][24] ),
    .I1(\reg_file.reg_storage[9][24] ),
    .I2(\reg_file.reg_storage[10][24] ),
    .I3(\reg_file.reg_storage[11][24] ),
    .S0(_2315_),
    .S1(_2316_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6219_ (.I(_0775_),
    .Z(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6220_ (.I0(_2317_),
    .I1(_2324_),
    .I2(_2326_),
    .I3(_2327_),
    .S0(_2223_),
    .S1(_2328_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6221_ (.A1(_2249_),
    .A2(_2314_),
    .B1(_2329_),
    .B2(_2250_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6222_ (.A1(_1434_),
    .A2(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6223_ (.A1(_2330_),
    .A2(_1434_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6224_ (.A1(_2331_),
    .A2(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6225_ (.A1(_1839_),
    .A2(_1948_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6226_ (.A1(_2236_),
    .A2(_2235_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6227_ (.A1(_2335_),
    .A2(_2247_),
    .A3(_2284_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6228_ (.A1(net196),
    .A2(_2148_),
    .A3(_2334_),
    .A4(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6229_ (.A1(_1735_),
    .A2(_1836_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6230_ (.A1(_1948_),
    .A2(_2338_),
    .B(_2032_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6231_ (.A1(_2025_),
    .A2(_2339_),
    .B(_2090_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6232_ (.A1(_2088_),
    .A2(_2340_),
    .B(_2143_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6233_ (.A1(_2335_),
    .A2(_2252_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6234_ (.A1(_2306_),
    .A2(_2342_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6235_ (.A1(_1389_),
    .A2(net179),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6236_ (.A1(_2341_),
    .A2(net167),
    .B1(_2343_),
    .B2(_2284_),
    .C(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6237_ (.A1(_1896_),
    .A2(_2337_),
    .B(_2345_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6238_ (.A1(_2333_),
    .A2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6239_ (.I(_2333_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6240_ (.A1(_2348_),
    .A2(_2346_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6241_ (.A1(_2035_),
    .A2(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6242_ (.A1(_2335_),
    .A2(_2240_),
    .A3(_2284_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6243_ (.A1(_2026_),
    .A2(_2147_),
    .A3(_2148_),
    .A4(_2351_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6244_ (.A1(_1842_),
    .A2(_1847_),
    .B(_2352_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6245_ (.A1(_2286_),
    .A2(_2241_),
    .B(_2282_),
    .C(_2235_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6246_ (.A1(_2152_),
    .A2(_2351_),
    .B(_2354_),
    .C(net189),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6247_ (.A1(_2353_),
    .A2(_2355_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6248_ (.A1(_2348_),
    .A2(_2356_),
    .B(_2096_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6249_ (.A1(_2348_),
    .A2(_2356_),
    .B(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6250_ (.A1(_1704_),
    .A2(_1389_),
    .B(_1435_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6251_ (.I0(_2257_),
    .I1(_2359_),
    .S(_1713_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6252_ (.I0(_2173_),
    .I1(_2360_),
    .S(_1993_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6253_ (.A1(_1978_),
    .A2(_1925_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6254_ (.I(_2038_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6255_ (.A1(_2050_),
    .A2(_2361_),
    .B(_2362_),
    .C(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6256_ (.I0(_1920_),
    .I1(_1929_),
    .S(_1986_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6257_ (.A1(_2290_),
    .A2(_2365_),
    .B(_1541_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6258_ (.A1(_1701_),
    .A2(_1900_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6259_ (.I(_2367_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6260_ (.I(_1597_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(_2332_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_2064_),
    .A2(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6263_ (.A1(_2062_),
    .A2(_2370_),
    .B(_2371_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6264_ (.A1(_2369_),
    .A2(_2372_),
    .B(_2331_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6265_ (.A1(_2364_),
    .A2(_2366_),
    .B1(_2368_),
    .B2(_1907_),
    .C(_2373_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6266_ (.A1(_2347_),
    .A2(_2350_),
    .B(_2358_),
    .C(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6267_ (.I(_2375_),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6268_ (.A1(net18),
    .A2(_0810_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6269_ (.A1(_2126_),
    .A2(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6270_ (.I0(\reg_file.reg_storage[4][25] ),
    .I1(\reg_file.reg_storage[5][25] ),
    .I2(\reg_file.reg_storage[6][25] ),
    .I3(\reg_file.reg_storage[7][25] ),
    .S0(_1153_),
    .S1(_0888_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6271_ (.I(\reg_file.reg_storage[1][25] ),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6272_ (.A1(_2315_),
    .A2(\reg_file.reg_storage[3][25] ),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6273_ (.A1(_0895_),
    .A2(\reg_file.reg_storage[2][25] ),
    .B(_1152_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6274_ (.A1(_2322_),
    .A2(_2379_),
    .B1(_2380_),
    .B2(_2381_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6275_ (.I0(\reg_file.reg_storage[12][25] ),
    .I1(\reg_file.reg_storage[13][25] ),
    .I2(\reg_file.reg_storage[14][25] ),
    .I3(\reg_file.reg_storage[15][25] ),
    .S0(_1153_),
    .S1(_1664_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6276_ (.I0(\reg_file.reg_storage[8][25] ),
    .I1(\reg_file.reg_storage[9][25] ),
    .I2(\reg_file.reg_storage[10][25] ),
    .I3(\reg_file.reg_storage[11][25] ),
    .S0(_1153_),
    .S1(_1664_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6277_ (.I0(_2378_),
    .I1(_2382_),
    .I2(_2383_),
    .I3(_2384_),
    .S0(_0900_),
    .S1(_0718_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6278_ (.A1(_0882_),
    .A2(_2377_),
    .B1(_2385_),
    .B2(_0902_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6279_ (.A1(_1418_),
    .A2(_2386_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6280_ (.I(_2387_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6281_ (.A1(_1720_),
    .A2(_2330_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6282_ (.A1(_2347_),
    .A2(_2389_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6283_ (.A1(_2388_),
    .A2(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6284_ (.I(_1682_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6285_ (.A1(_2388_),
    .A2(_2390_),
    .B(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6286_ (.A1(_2348_),
    .A2(_2356_),
    .B(_2370_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6287_ (.A1(_2388_),
    .A2(_2394_),
    .B(_2096_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6288_ (.A1(_2388_),
    .A2(_2394_),
    .B(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6289_ (.I(_2386_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6290_ (.A1(_1418_),
    .A2(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6291_ (.I(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6292_ (.A1(_1601_),
    .A2(_2398_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6293_ (.A1(_1419_),
    .A2(_2397_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6294_ (.A1(_2369_),
    .A2(_2400_),
    .B(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6295_ (.A1(_2201_),
    .A2(_2006_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6296_ (.A1(_1243_),
    .A2(_1976_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6297_ (.A1(_1789_),
    .A2(_1969_),
    .B(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6298_ (.I(_1419_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6299_ (.A1(_1707_),
    .A2(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6300_ (.A1(_1710_),
    .A2(net211),
    .B(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6301_ (.I0(_2291_),
    .I1(_2408_),
    .S(_1973_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6302_ (.A1(_2167_),
    .A2(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6303_ (.A1(_2160_),
    .A2(_2203_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6304_ (.A1(_1998_),
    .A2(_2410_),
    .A3(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6305_ (.A1(_1789_),
    .A2(_1982_),
    .B(_2412_),
    .C(_2176_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6306_ (.A1(_2046_),
    .A2(_2405_),
    .B(_2413_),
    .C(_1919_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6307_ (.A1(_1997_),
    .A2(_2403_),
    .B(_2414_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6308_ (.A1(_1960_),
    .A2(_2399_),
    .B(_2402_),
    .C(_2415_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6309_ (.A1(_2391_),
    .A2(_2393_),
    .B(_2396_),
    .C(_2416_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6310_ (.I(_2417_),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6311_ (.I(_0844_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6312_ (.A1(net19),
    .A2(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6313_ (.A1(_2272_),
    .A2(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6314_ (.I0(\reg_file.reg_storage[4][26] ),
    .I1(\reg_file.reg_storage[5][26] ),
    .I2(\reg_file.reg_storage[6][26] ),
    .I3(\reg_file.reg_storage[7][26] ),
    .S0(_1667_),
    .S1(_2325_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6315_ (.A1(_0756_),
    .A2(\reg_file.reg_storage[3][26] ),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6316_ (.A1(_2076_),
    .A2(\reg_file.reg_storage[2][26] ),
    .B(_2322_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6317_ (.A1(_1823_),
    .A2(_1329_),
    .B1(_2422_),
    .B2(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6318_ (.I0(\reg_file.reg_storage[12][26] ),
    .I1(\reg_file.reg_storage[13][26] ),
    .I2(\reg_file.reg_storage[14][26] ),
    .I3(\reg_file.reg_storage[15][26] ),
    .S0(_2072_),
    .S1(_2073_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6319_ (.I0(\reg_file.reg_storage[8][26] ),
    .I1(\reg_file.reg_storage[9][26] ),
    .I2(\reg_file.reg_storage[10][26] ),
    .I3(\reg_file.reg_storage[11][26] ),
    .S0(_2072_),
    .S1(_2073_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6320_ (.I0(_2421_),
    .I1(_2424_),
    .I2(_2425_),
    .I3(_2426_),
    .S0(_2082_),
    .S1(_1833_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6321_ (.A1(_2070_),
    .A2(_2420_),
    .B1(_2427_),
    .B2(_2084_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6322_ (.A1(_1340_),
    .A2(_2428_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6323_ (.A1(_1341_),
    .A2(net169),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6324_ (.A1(_2429_),
    .A2(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6325_ (.I(_2431_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6326_ (.I(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6327_ (.A1(_2331_),
    .A2(_2370_),
    .A3(_2387_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6328_ (.I(_2332_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6329_ (.A1(_2435_),
    .A2(_2398_),
    .B(_2401_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6330_ (.A1(_2356_),
    .A2(_2434_),
    .B(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6331_ (.A1(_2433_),
    .A2(_2437_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6332_ (.I(_1813_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6333_ (.A1(_2433_),
    .A2(_2437_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(_2439_),
    .A2(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6335_ (.A1(_1418_),
    .A2(_2386_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6336_ (.A1(_2391_),
    .A2(_2433_),
    .A3(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6337_ (.A1(_2391_),
    .A2(_2442_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6338_ (.A1(_2432_),
    .A2(_2444_),
    .B(_2392_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6339_ (.A1(_1420_),
    .A2(_1342_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6340_ (.I0(_2359_),
    .I1(_2446_),
    .S(_1309_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6341_ (.I0(_2258_),
    .I1(_2447_),
    .S(_2167_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6342_ (.I0(_2043_),
    .I1(_2448_),
    .S(_2169_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6343_ (.A1(_1687_),
    .A2(_1586_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _6344_ (.A1(_1562_),
    .A2(_2044_),
    .B1(_2450_),
    .B2(_2158_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6345_ (.A1(_2046_),
    .A2(_2451_),
    .B(_1793_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6346_ (.A1(_2039_),
    .A2(_2449_),
    .B(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6347_ (.I(_2430_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6348_ (.A1(_2064_),
    .A2(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6349_ (.A1(_2062_),
    .A2(_2454_),
    .B(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6350_ (.A1(_2369_),
    .A2(_2456_),
    .B(_2429_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6351_ (.A1(_2057_),
    .A2(_2368_),
    .B(_2453_),
    .C(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6352_ (.A1(_2438_),
    .A2(_2441_),
    .B1(_2443_),
    .B2(_2445_),
    .C(_2458_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6353_ (.I(_2459_),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6354_ (.A1(_1276_),
    .A2(_1319_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6355_ (.A1(_1403_),
    .A2(_1325_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6356_ (.A1(net84),
    .A2(_0866_),
    .B1(_2460_),
    .B2(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6357_ (.A1(net20),
    .A2(_0810_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6358_ (.A1(_2272_),
    .A2(_2463_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6359_ (.I0(\reg_file.reg_storage[4][27] ),
    .I1(\reg_file.reg_storage[5][27] ),
    .I2(\reg_file.reg_storage[6][27] ),
    .I3(\reg_file.reg_storage[7][27] ),
    .S0(_0767_),
    .S1(_2011_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6360_ (.A1(_2013_),
    .A2(\reg_file.reg_storage[3][27] ),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6361_ (.A1(_1827_),
    .A2(\reg_file.reg_storage[2][27] ),
    .B(_0584_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6362_ (.A1(_0890_),
    .A2(_1314_),
    .B1(_2466_),
    .B2(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6363_ (.I0(\reg_file.reg_storage[12][27] ),
    .I1(\reg_file.reg_storage[13][27] ),
    .I2(\reg_file.reg_storage[14][27] ),
    .I3(\reg_file.reg_storage[15][27] ),
    .S0(_0887_),
    .S1(_2017_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _6364_ (.I0(\reg_file.reg_storage[8][27] ),
    .I1(\reg_file.reg_storage[9][27] ),
    .I2(\reg_file.reg_storage[10][27] ),
    .I3(\reg_file.reg_storage[11][27] ),
    .S0(_0767_),
    .S1(_2017_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6365_ (.I0(_2465_),
    .I1(_2468_),
    .I2(_2469_),
    .I3(_2470_),
    .S0(_1832_),
    .S1(_2020_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6366_ (.A1(_1819_),
    .A2(_2464_),
    .B1(_2471_),
    .B2(_1835_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6367_ (.A1(_2462_),
    .A2(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6368_ (.A1(_2462_),
    .A2(_2472_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6369_ (.A1(_2473_),
    .A2(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6370_ (.A1(_2454_),
    .A2(_2438_),
    .A3(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6371_ (.A1(_2454_),
    .A2(_2438_),
    .B(_2475_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6372_ (.A1(_2439_),
    .A2(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6373_ (.A1(_2052_),
    .A2(_1765_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6374_ (.A1(_1998_),
    .A2(_2102_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6375_ (.A1(_2169_),
    .A2(_2479_),
    .B(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6376_ (.A1(_1711_),
    .A2(_1717_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6377_ (.I0(_2408_),
    .I1(_2482_),
    .S(_1309_),
    .Z(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6378_ (.A1(_1692_),
    .A2(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6379_ (.A1(_1787_),
    .A2(_2292_),
    .B(_1977_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6380_ (.A1(_1970_),
    .A2(_2107_),
    .B1(_2484_),
    .B2(_2485_),
    .C(_1536_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6381_ (.A1(_2109_),
    .A2(_2481_),
    .B(_2486_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6382_ (.A1(_1794_),
    .A2(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6383_ (.I(_2474_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6384_ (.I(_1801_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6385_ (.I(_1596_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6386_ (.A1(_2490_),
    .A2(_2489_),
    .B(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6387_ (.A1(_2462_),
    .A2(_2472_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6388_ (.A1(_2302_),
    .A2(_2489_),
    .B1(_2492_),
    .B2(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6389_ (.A1(_2116_),
    .A2(_2403_),
    .B(_2488_),
    .C(_2494_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6390_ (.I(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6391_ (.A1(_2473_),
    .A2(_2489_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6392_ (.I(_1341_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6393_ (.A1(_2498_),
    .A2(_2428_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6394_ (.A1(_2432_),
    .A2(_2444_),
    .B(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6395_ (.I(_1231_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6396_ (.A1(_2497_),
    .A2(_2500_),
    .B(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6397_ (.A1(_2497_),
    .A2(_2500_),
    .B(_2502_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6398_ (.A1(_2476_),
    .A2(_2478_),
    .B(_2496_),
    .C(_2503_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6399_ (.I(_2504_),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6400_ (.I(_1657_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6401_ (.I(_2505_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6402_ (.A1(net21),
    .A2(_2418_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6403_ (.A1(_2272_),
    .A2(_2507_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6404_ (.I0(\reg_file.reg_storage[4][28] ),
    .I1(\reg_file.reg_storage[5][28] ),
    .I2(\reg_file.reg_storage[6][28] ),
    .I3(\reg_file.reg_storage[7][28] ),
    .S0(_0711_),
    .S1(_2079_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6405_ (.A1(_0756_),
    .A2(\reg_file.reg_storage[3][28] ),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6406_ (.A1(_2076_),
    .A2(\reg_file.reg_storage[2][28] ),
    .B(_1666_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6407_ (.A1(_1823_),
    .A2(_1363_),
    .B1(_2510_),
    .B2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6408_ (.I0(\reg_file.reg_storage[12][28] ),
    .I1(\reg_file.reg_storage[13][28] ),
    .I2(\reg_file.reg_storage[14][28] ),
    .I3(\reg_file.reg_storage[15][28] ),
    .S0(_0813_),
    .S1(_1821_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6409_ (.I0(\reg_file.reg_storage[8][28] ),
    .I1(\reg_file.reg_storage[9][28] ),
    .I2(\reg_file.reg_storage[10][28] ),
    .I3(\reg_file.reg_storage[11][28] ),
    .S0(_0813_),
    .S1(_2079_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6410_ (.I0(_2509_),
    .I1(_2512_),
    .I2(_2513_),
    .I3(_2514_),
    .S0(_2082_),
    .S1(_1833_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6411_ (.A1(_2070_),
    .A2(_2508_),
    .B1(_2515_),
    .B2(_2084_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6412_ (.A1(_1371_),
    .A2(_2516_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6413_ (.I(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6414_ (.A1(_1370_),
    .A2(_2516_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6415_ (.I(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6416_ (.A1(_2518_),
    .A2(_2520_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6417_ (.I(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6418_ (.A1(_2432_),
    .A2(_2434_),
    .A3(_2475_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6419_ (.A1(_2353_),
    .A2(_2355_),
    .B(_2523_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6420_ (.A1(_2430_),
    .A2(_2436_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6421_ (.A1(_2429_),
    .A2(_2525_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6422_ (.A1(_2489_),
    .A2(_2526_),
    .B(_2493_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6423_ (.I(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6424_ (.A1(_2524_),
    .A2(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6425_ (.A1(_2522_),
    .A2(_2529_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6426_ (.A1(_2401_),
    .A2(_2399_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _6427_ (.A1(_2333_),
    .A2(_2531_),
    .A3(_2431_),
    .A4(_2475_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6428_ (.A1(_2387_),
    .A2(_2389_),
    .B(_2442_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6429_ (.A1(_2431_),
    .A2(_2533_),
    .B(_2499_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6430_ (.A1(_1327_),
    .A2(_2472_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6431_ (.A1(_2497_),
    .A2(_2534_),
    .B(_2535_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6432_ (.A1(net202),
    .A2(_2532_),
    .B(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6433_ (.A1(_2521_),
    .A2(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6434_ (.A1(_2537_),
    .A2(_2521_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6435_ (.A1(_2392_),
    .A2(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6436_ (.A1(_1986_),
    .A2(_2171_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6437_ (.A1(_1978_),
    .A2(_2168_),
    .B(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6438_ (.A1(_2115_),
    .A2(_2174_),
    .B(_2109_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6439_ (.I(_2055_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6440_ (.I(_1695_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6441_ (.A1(_1704_),
    .A2(_1327_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6442_ (.A1(_2546_),
    .A2(_1372_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6443_ (.I(_1713_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6444_ (.A1(_2548_),
    .A2(_2446_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6445_ (.A1(_2545_),
    .A2(_2547_),
    .B(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6446_ (.A1(_2052_),
    .A2(_2360_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6447_ (.A1(_2544_),
    .A2(_2550_),
    .B(_2551_),
    .C(_1546_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6448_ (.A1(_2363_),
    .A2(_2542_),
    .B1(_2543_),
    .B2(_2552_),
    .C(_1794_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6449_ (.I(_1801_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6450_ (.A1(_2554_),
    .A2(_2519_),
    .B(_2491_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6451_ (.A1(_2159_),
    .A2(_2368_),
    .B1(_2518_),
    .B2(_2555_),
    .C1(_2519_),
    .C2(_2302_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6452_ (.A1(_2553_),
    .A2(_2556_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6453_ (.A1(_2506_),
    .A2(_2530_),
    .B1(_2538_),
    .B2(_2540_),
    .C(_2557_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6454_ (.I(_2558_),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6455_ (.A1(net22),
    .A2(_2418_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6456_ (.A1(_2312_),
    .A2(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6457_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(\reg_file.reg_storage[5][29] ),
    .I2(\reg_file.reg_storage[6][29] ),
    .I3(\reg_file.reg_storage[7][29] ),
    .S0(_1667_),
    .S1(_2325_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6458_ (.A1(_2320_),
    .A2(\reg_file.reg_storage[3][29] ),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6459_ (.A1(_2076_),
    .A2(\reg_file.reg_storage[2][29] ),
    .B(_2322_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6460_ (.A1(_2318_),
    .A2(_1349_),
    .B1(_2562_),
    .B2(_2563_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6461_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(\reg_file.reg_storage[13][29] ),
    .I2(\reg_file.reg_storage[14][29] ),
    .I3(\reg_file.reg_storage[15][29] ),
    .S0(_2072_),
    .S1(_2073_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6462_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(\reg_file.reg_storage[9][29] ),
    .I2(\reg_file.reg_storage[10][29] ),
    .I3(\reg_file.reg_storage[11][29] ),
    .S0(_1667_),
    .S1(_2325_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6463_ (.I0(_2561_),
    .I1(_2564_),
    .I2(_2565_),
    .I3(_2566_),
    .S0(_2082_),
    .S1(_2328_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6464_ (.A1(_2070_),
    .A2(_2560_),
    .B1(_2567_),
    .B2(_2084_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6465_ (.I(_2568_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6466_ (.A1(_1359_),
    .A2(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6467_ (.I(_1358_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6468_ (.A1(_2571_),
    .A2(_2568_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6469_ (.A1(_2570_),
    .A2(_2572_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6470_ (.A1(_2524_),
    .A2(_2528_),
    .B(_2518_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6471_ (.A1(_2520_),
    .A2(_2573_),
    .A3(_2574_),
    .Z(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6472_ (.A1(_2520_),
    .A2(_2574_),
    .B(_2573_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6473_ (.I(_2573_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6474_ (.I(_1371_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6475_ (.A1(_2578_),
    .A2(_2516_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6476_ (.A1(_2539_),
    .A2(_2577_),
    .A3(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6477_ (.A1(_2539_),
    .A2(_2579_),
    .B(_2577_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6478_ (.A1(_1897_),
    .A2(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6479_ (.A1(_1545_),
    .A2(_2209_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6480_ (.A1(_1701_),
    .A2(_2206_),
    .B(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6481_ (.A1(_2051_),
    .A2(_2409_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6482_ (.A1(_1710_),
    .A2(_1359_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6483_ (.A1(_2586_),
    .A2(_1708_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6484_ (.A1(_1575_),
    .A2(_2587_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6485_ (.A1(_1994_),
    .A2(_2482_),
    .B(_2588_),
    .C(_1988_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6486_ (.A1(_1977_),
    .A2(_2585_),
    .A3(_2589_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6487_ (.A1(_1442_),
    .A2(_2204_),
    .B(_2590_),
    .C(_1688_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6488_ (.A1(_2176_),
    .A2(_2584_),
    .B(_2591_),
    .C(_1793_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6489_ (.I(_2570_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6490_ (.I(_2572_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6491_ (.A1(_1800_),
    .A2(_2594_),
    .B(_1596_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6492_ (.A1(_2212_),
    .A2(_2367_),
    .B1(_2593_),
    .B2(_2595_),
    .C1(_2594_),
    .C2(_1798_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6493_ (.A1(_2592_),
    .A2(_2596_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6494_ (.A1(_2580_),
    .A2(_2582_),
    .B(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _6495_ (.A1(_2096_),
    .A2(_2575_),
    .A3(_2576_),
    .B(_2598_),
    .ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6496_ (.A1(net24),
    .A2(_2418_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6497_ (.A1(_2312_),
    .A2(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6498_ (.I(_0764_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6499_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(\reg_file.reg_storage[5][30] ),
    .I2(\reg_file.reg_storage[6][30] ),
    .I3(\reg_file.reg_storage[7][30] ),
    .S0(_0893_),
    .S1(_2601_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6500_ (.A1(_2320_),
    .A2(\reg_file.reg_storage[3][30] ),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6501_ (.A1(_2123_),
    .A2(\reg_file.reg_storage[2][30] ),
    .B(_0890_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6502_ (.A1(_2318_),
    .A2(_1264_),
    .B1(_2603_),
    .B2(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6503_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(\reg_file.reg_storage[13][30] ),
    .I2(\reg_file.reg_storage[14][30] ),
    .I3(\reg_file.reg_storage[15][30] ),
    .S0(_0893_),
    .S1(_2316_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6504_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(\reg_file.reg_storage[9][30] ),
    .I2(\reg_file.reg_storage[10][30] ),
    .I3(\reg_file.reg_storage[11][30] ),
    .S0(_0893_),
    .S1(_2316_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6505_ (.I0(_2602_),
    .I1(_2605_),
    .I2(_2606_),
    .I3(_2607_),
    .S0(_2223_),
    .S1(_2328_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6506_ (.A1(_2249_),
    .A2(_2600_),
    .B1(_2608_),
    .B2(_2250_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6507_ (.A1(_1279_),
    .A2(_2609_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6508_ (.A1(net200),
    .A2(_2609_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6509_ (.I(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6510_ (.A1(_2612_),
    .A2(_2610_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6511_ (.I(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6512_ (.A1(_2520_),
    .A2(_2574_),
    .B(_2570_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6513_ (.A1(_2594_),
    .A2(_2615_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6514_ (.A1(_2614_),
    .A2(_2616_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6515_ (.A1(_2571_),
    .A2(_2569_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6516_ (.A1(_2581_),
    .A2(_2613_),
    .A3(_2618_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6517_ (.A1(_2581_),
    .A2(_2618_),
    .B(_2613_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6518_ (.A1(_2392_),
    .A2(_2619_),
    .A3(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6519_ (.A1(_1280_),
    .A2(_1360_),
    .B(_1575_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6520_ (.A1(_1713_),
    .A2(_2547_),
    .B(_2622_),
    .C(_1377_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6521_ (.A1(_2167_),
    .A2(_2447_),
    .B(_2623_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6522_ (.A1(_2264_),
    .A2(_2624_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6523_ (.A1(_1789_),
    .A2(_2259_),
    .B(_2625_),
    .C(_2176_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6524_ (.A1(_1537_),
    .A2(_1590_),
    .B(_2626_),
    .C(_1919_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6525_ (.A1(_1798_),
    .A2(_2611_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6526_ (.A1(_2490_),
    .A2(_2611_),
    .B(_2628_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6527_ (.A1(_1917_),
    .A2(_2629_),
    .B(_2610_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6528_ (.A1(_2544_),
    .A2(_1301_),
    .A3(_2368_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6529_ (.A1(_2505_),
    .A2(_2627_),
    .A3(_2630_),
    .A4(_2631_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6530_ (.A1(_2621_),
    .A2(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6531_ (.A1(_2506_),
    .A2(_2617_),
    .B(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _6532_ (.I(_2634_),
    .ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6533_ (.A1(_2594_),
    .A2(_2615_),
    .B(_2614_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6534_ (.I0(\reg_file.reg_storage[4][31] ),
    .I1(\reg_file.reg_storage[5][31] ),
    .I2(\reg_file.reg_storage[6][31] ),
    .I3(\reg_file.reg_storage[7][31] ),
    .S0(_1825_),
    .S1(_2601_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6535_ (.A1(_2320_),
    .A2(\reg_file.reg_storage[3][31] ),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6536_ (.A1(_2123_),
    .A2(\reg_file.reg_storage[2][31] ),
    .B(_2182_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6537_ (.A1(_2318_),
    .A2(_1288_),
    .B1(_2637_),
    .B2(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6538_ (.I0(\reg_file.reg_storage[12][31] ),
    .I1(\reg_file.reg_storage[13][31] ),
    .I2(\reg_file.reg_storage[14][31] ),
    .I3(\reg_file.reg_storage[15][31] ),
    .S0(_2013_),
    .S1(_2601_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6539_ (.I0(\reg_file.reg_storage[8][31] ),
    .I1(\reg_file.reg_storage[9][31] ),
    .I2(\reg_file.reg_storage[10][31] ),
    .I3(\reg_file.reg_storage[11][31] ),
    .S0(_2013_),
    .S1(_2601_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _6540_ (.I0(_2636_),
    .I1(_2639_),
    .I2(_2640_),
    .I3(_2641_),
    .S0(_2223_),
    .S1(_2328_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6541_ (.A1(_0746_),
    .A2(_2249_),
    .B1(_2250_),
    .B2(_2642_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6542_ (.A1(_1298_),
    .A2(_2643_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6543_ (.A1(_1298_),
    .A2(_2643_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6544_ (.A1(_2644_),
    .A2(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6545_ (.I(_2646_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6546_ (.A1(_2612_),
    .A2(_2635_),
    .B(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6547_ (.A1(_2612_),
    .A2(_2635_),
    .A3(_2647_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6548_ (.I(_1443_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6549_ (.A1(_1254_),
    .A2(_2586_),
    .A3(_1708_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6550_ (.A1(_1254_),
    .A2(_1705_),
    .B(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6551_ (.A1(_1990_),
    .A2(_1699_),
    .A3(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6552_ (.A1(_1693_),
    .A2(_2483_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6553_ (.A1(_1303_),
    .A2(_2653_),
    .A3(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6554_ (.A1(_2650_),
    .A2(_2293_),
    .B(_2655_),
    .C(_2099_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6555_ (.A1(_2290_),
    .A2(_1790_),
    .B(_1541_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _6556_ (.I(_2647_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6557_ (.I(_2609_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6558_ (.A1(_1279_),
    .A2(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6559_ (.I(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6560_ (.A1(_2620_),
    .A2(_2658_),
    .A3(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6561_ (.A1(_2620_),
    .A2(_2661_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6562_ (.A1(_2647_),
    .A2(_2663_),
    .B(_2501_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6563_ (.I(_2643_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6564_ (.A1(_1299_),
    .A2(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6565_ (.A1(_2064_),
    .A2(_2645_),
    .B(_2060_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6566_ (.A1(_1601_),
    .A2(_2645_),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6567_ (.A1(_2100_),
    .A2(_1699_),
    .A3(_2403_),
    .B1(_2666_),
    .B2(_2668_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6568_ (.A1(_2656_),
    .A2(_2657_),
    .B1(_2662_),
    .B2(_2664_),
    .C(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _6569_ (.A1(_2506_),
    .A2(_2648_),
    .A3(_2649_),
    .B(_2670_),
    .ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6570_ (.A1(_2613_),
    .A2(_2646_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6571_ (.A1(_2522_),
    .A2(_2536_),
    .B(_2579_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6572_ (.A1(_2573_),
    .A2(_2672_),
    .B(_2618_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _6573_ (.A1(_2522_),
    .A2(_2532_),
    .A3(_2577_),
    .A4(_2671_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _6574_ (.A1(_1298_),
    .A2(_2665_),
    .B1(_2671_),
    .B2(_2673_),
    .C1(_2674_),
    .C2(_2346_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6575_ (.A1(_1592_),
    .A2(_2658_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6576_ (.A1(_2658_),
    .A2(_2661_),
    .B(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6577_ (.I(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6578_ (.A1(_1235_),
    .A2(_1540_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6579_ (.A1(_2675_),
    .A2(_2678_),
    .B(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6580_ (.A1(net215),
    .A2(_2676_),
    .B(_2680_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6581_ (.A1(_1564_),
    .A2(_1570_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6582_ (.A1(_1550_),
    .A2(_1565_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6583_ (.I0(_2682_),
    .I1(_2683_),
    .S(_1252_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6584_ (.A1(_1567_),
    .A2(_1583_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6585_ (.A1(_1577_),
    .A2(_1696_),
    .B(_2685_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6586_ (.A1(_1576_),
    .A2(_1583_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6587_ (.A1(_1257_),
    .A2(_1630_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6588_ (.A1(_2687_),
    .A2(_2688_),
    .B(_1574_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6589_ (.A1(_1308_),
    .A2(_2686_),
    .B(_2689_),
    .C(_1248_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6590_ (.A1(_1249_),
    .A2(_2684_),
    .B(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6591_ (.A1(_1547_),
    .A2(_1551_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6592_ (.A1(_1200_),
    .A2(_1378_),
    .B(_1548_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6593_ (.I0(_2692_),
    .I1(_2693_),
    .S(_1904_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6594_ (.A1(_1554_),
    .A2(_1558_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6595_ (.I0(_1456_),
    .I1(_2695_),
    .S(_1307_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6596_ (.I0(_2694_),
    .I1(_2696_),
    .S(_1304_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6597_ (.A1(_1440_),
    .A2(_2697_),
    .B(_1534_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6598_ (.A1(_1241_),
    .A2(_2691_),
    .B(_2698_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6599_ (.A1(_1168_),
    .A2(_1912_),
    .B(_2699_),
    .C(_1652_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6600_ (.A1(_1556_),
    .A2(_1630_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6601_ (.I(_2701_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6602_ (.A1(_1231_),
    .A2(_1800_),
    .B(_2702_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6603_ (.A1(_1916_),
    .A2(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6604_ (.A1(_1440_),
    .A2(_1542_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6605_ (.A1(_1920_),
    .A2(_2705_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6606_ (.A1(_1797_),
    .A2(_2702_),
    .B(_1811_),
    .C(_2706_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6607_ (.A1(_2701_),
    .A2(_2688_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6608_ (.A1(_0991_),
    .A2(_1235_),
    .A3(_1655_),
    .A4(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _6609_ (.A1(net195),
    .A2(_2148_),
    .A3(_2334_),
    .A4(_2336_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6610_ (.A1(net204),
    .A2(_2710_),
    .A3(_2674_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6611_ (.A1(_0965_),
    .A2(net217),
    .A3(_2709_),
    .A4(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6612_ (.A1(_2688_),
    .A2(_2704_),
    .B(_2707_),
    .C(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _6613_ (.A1(_2681_),
    .A2(_2700_),
    .A3(_2713_),
    .B1(_2708_),
    .B2(_1656_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _6614_ (.I(_2714_),
    .ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6615_ (.I(_2046_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6616_ (.A1(_1197_),
    .A2(_1704_),
    .B(_1774_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6617_ (.A1(_1776_),
    .A2(_1780_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6618_ (.I0(_2716_),
    .I1(_2717_),
    .S(_1487_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6619_ (.A1(_1779_),
    .A2(_1782_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6620_ (.I0(_1737_),
    .I1(_2719_),
    .S(_1575_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6621_ (.I0(_2718_),
    .I1(_2720_),
    .S(_2160_),
    .Z(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6622_ (.A1(_1766_),
    .A2(_1773_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6623_ (.I(_1697_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6624_ (.A1(_2723_),
    .A2(_1175_),
    .B(_1769_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6625_ (.I0(_2722_),
    .I1(_2724_),
    .S(_1757_),
    .Z(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6626_ (.A1(_2723_),
    .A2(_1768_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6627_ (.A1(_1053_),
    .A2(_2723_),
    .B(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6628_ (.A1(_1758_),
    .A2(_2723_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6629_ (.A1(_2728_),
    .A2(_1763_),
    .B(_1757_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6630_ (.A1(_2548_),
    .A2(_2727_),
    .B(_2729_),
    .C(_2055_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6631_ (.A1(_1993_),
    .A2(_2725_),
    .B(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6632_ (.A1(_2201_),
    .A2(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6633_ (.A1(_1987_),
    .A2(_2721_),
    .B(_2732_),
    .C(_1791_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6634_ (.A1(_2715_),
    .A2(_2005_),
    .B(_2733_),
    .C(_1238_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6635_ (.A1(_1969_),
    .A2(_2705_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6636_ (.I0(_1603_),
    .I1(_2490_),
    .S(_1631_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6637_ (.A1(_2545_),
    .A2(_1040_),
    .B1(_2061_),
    .B2(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6638_ (.A1(_2735_),
    .A2(_2737_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6639_ (.I(_0991_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6640_ (.A1(_2739_),
    .A2(_2702_),
    .B(_2505_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6641_ (.A1(_2739_),
    .A2(_2702_),
    .B(_2740_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6642_ (.A1(_2739_),
    .A2(_1762_),
    .B(_1897_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6643_ (.A1(_2739_),
    .A2(_1762_),
    .B(_2742_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _6644_ (.A1(_2734_),
    .A2(_2738_),
    .A3(_2741_),
    .A4(_2743_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6645_ (.I(_2744_),
    .ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6646_ (.I(net227),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6647_ (.A1(_2745_),
    .A2(_1632_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6648_ (.I0(_2693_),
    .I1(_2695_),
    .S(_1373_),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6649_ (.I0(_1488_),
    .I1(_2747_),
    .S(_1787_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6650_ (.A1(_2548_),
    .A2(_2686_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6651_ (.A1(_2545_),
    .A2(_2682_),
    .B(_2749_),
    .C(_1990_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6652_ (.I0(_2683_),
    .I1(_2692_),
    .S(_1373_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6653_ (.A1(_1693_),
    .A2(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6654_ (.A1(_1303_),
    .A2(_2750_),
    .A3(_2752_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6655_ (.A1(_2650_),
    .A2(_2748_),
    .B(_2753_),
    .C(_2039_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6656_ (.A1(_2715_),
    .A2(_2059_),
    .B(_2754_),
    .C(_1239_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6657_ (.A1(_1633_),
    .A2(_2554_),
    .B(_2491_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6658_ (.A1(_1633_),
    .A2(_2216_),
    .B1(_2756_),
    .B2(_1627_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6659_ (.A1(_1953_),
    .A2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6660_ (.A1(_2745_),
    .A2(_1868_),
    .B(_1682_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6661_ (.A1(_2745_),
    .A2(_1868_),
    .B(_2759_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6662_ (.A1(_1544_),
    .A2(_2047_),
    .B(_2758_),
    .C(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6663_ (.A1(_2439_),
    .A2(_2746_),
    .B1(_2755_),
    .B2(_2761_),
    .ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6664_ (.I0(_2717_),
    .I1(_2719_),
    .S(_1254_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6665_ (.I0(_1738_),
    .I1(_2762_),
    .S(_1787_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6666_ (.A1(_2548_),
    .A2(_2727_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6667_ (.A1(_2545_),
    .A2(_2724_),
    .B(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6668_ (.I0(_2716_),
    .I1(_2722_),
    .S(_1695_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6669_ (.A1(_2158_),
    .A2(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6670_ (.A1(_2100_),
    .A2(_2765_),
    .B(_2767_),
    .C(_2201_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6671_ (.A1(_1987_),
    .A2(_2763_),
    .B(_2768_),
    .C(_2363_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6672_ (.A1(_2715_),
    .A2(_2119_),
    .B(_2769_),
    .C(_1238_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6673_ (.A1(net197),
    .A2(_1634_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6674_ (.A1(_1818_),
    .A2(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6675_ (.I(_1047_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6676_ (.A1(_2745_),
    .A2(_1868_),
    .B(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6677_ (.A1(net197),
    .A2(_2774_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6678_ (.A1(_2035_),
    .A2(_2775_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6679_ (.I(_1542_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6680_ (.A1(_1635_),
    .A2(_1802_),
    .B(_2061_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _6681_ (.A1(_1635_),
    .A2(_1799_),
    .B1(_2101_),
    .B2(_2777_),
    .C1(_2778_),
    .C2(_1625_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6682_ (.A1(_2770_),
    .A2(_2772_),
    .A3(_2776_),
    .A4(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6683_ (.I(_2780_),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6684_ (.I(_1754_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6685_ (.A1(_2781_),
    .A2(_2163_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6686_ (.A1(_2544_),
    .A2(_2694_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6687_ (.A1(_1693_),
    .A2(_2684_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6688_ (.I0(_1908_),
    .I1(_2696_),
    .S(_1250_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6689_ (.A1(_1702_),
    .A2(_2785_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6690_ (.A1(_2054_),
    .A2(_2783_),
    .A3(_2784_),
    .B(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6691_ (.A1(_2099_),
    .A2(_2787_),
    .B(_1686_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6692_ (.I(_1086_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6693_ (.A1(_1870_),
    .A2(_2789_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6694_ (.A1(_1639_),
    .A2(_1913_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6695_ (.I(_1639_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6696_ (.A1(_2792_),
    .A2(_1600_),
    .B(_1916_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6697_ (.A1(_2109_),
    .A2(_1569_),
    .B1(_2791_),
    .B2(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6698_ (.I(_2794_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6699_ (.A1(_2168_),
    .A2(_2705_),
    .B1(_2790_),
    .B2(_2501_),
    .C(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6700_ (.A1(_2789_),
    .A2(_1637_),
    .B(_1817_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6701_ (.A1(_2789_),
    .A2(_1637_),
    .B(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6702_ (.A1(_2782_),
    .A2(_2788_),
    .B(_2796_),
    .C(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6703_ (.I(net166),
    .ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6704_ (.I(_1238_),
    .Z(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6705_ (.I0(_2000_),
    .I1(_2720_),
    .S(_1563_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6706_ (.A1(_2544_),
    .A2(_2725_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6707_ (.A1(_2100_),
    .A2(_2718_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6708_ (.A1(_1987_),
    .A2(_2802_),
    .A3(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6709_ (.A1(_2650_),
    .A2(_2801_),
    .B(_2804_),
    .C(_2099_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6710_ (.A1(_2781_),
    .A2(_2215_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6711_ (.A1(_2800_),
    .A2(_2805_),
    .A3(_2806_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6712_ (.A1(_1638_),
    .A2(_1964_),
    .B(_2369_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6713_ (.I(_1623_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _6714_ (.A1(_1638_),
    .A2(_1960_),
    .B1(_2210_),
    .B2(_2777_),
    .C1(_2808_),
    .C2(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6715_ (.A1(_2789_),
    .A2(_1637_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6716_ (.A1(_2792_),
    .A2(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6717_ (.A1(_1136_),
    .A2(_2812_),
    .Z(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6718_ (.I(_1086_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6719_ (.A1(_1870_),
    .A2(_2814_),
    .B(_1873_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6720_ (.A1(_1136_),
    .A2(_2815_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6721_ (.A1(_1136_),
    .A2(_2815_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6722_ (.A1(_1898_),
    .A2(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6723_ (.A1(_1818_),
    .A2(_2813_),
    .B1(_2816_),
    .B2(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6724_ (.A1(_2807_),
    .A2(_2810_),
    .A3(_2819_),
    .ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6725_ (.A1(_1165_),
    .A2(_1623_),
    .A3(_1640_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6726_ (.A1(_1623_),
    .A2(_1640_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6727_ (.A1(_1111_),
    .A2(_2821_),
    .B(_1818_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6728_ (.A1(_1874_),
    .A2(_2817_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6729_ (.A1(_1111_),
    .A2(_2823_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6730_ (.A1(_1111_),
    .A2(_2823_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6731_ (.A1(_2308_),
    .A2(_2825_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6732_ (.A1(_1619_),
    .A2(_2490_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6733_ (.A1(_1619_),
    .A2(_2216_),
    .B(_2827_),
    .C(_1917_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6734_ (.A1(_1971_),
    .A2(_1543_),
    .A3(_1588_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6735_ (.A1(_2160_),
    .A2(_2747_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6736_ (.A1(_1724_),
    .A2(_2751_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6737_ (.A1(_2264_),
    .A2(_2830_),
    .A3(_2831_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6738_ (.A1(_2103_),
    .A2(_1532_),
    .B(_2832_),
    .C(_2038_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6739_ (.A1(_1791_),
    .A2(_2266_),
    .B(_2833_),
    .C(_1237_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6740_ (.A1(_1109_),
    .A2(_2828_),
    .B(_2829_),
    .C(_2834_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6741_ (.A1(_2824_),
    .A2(_2826_),
    .B(_2835_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6742_ (.A1(_2820_),
    .A2(_2822_),
    .B(_2836_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6743_ (.I(_2837_),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6744_ (.A1(_1619_),
    .A2(_2820_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6745_ (.A1(_1624_),
    .A2(_2838_),
    .B(_1953_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6746_ (.A1(_1624_),
    .A2(_2838_),
    .B(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6747_ (.A1(_2158_),
    .A2(_2766_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6748_ (.A1(_1990_),
    .A2(_2762_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6749_ (.A1(_2841_),
    .A2(_2842_),
    .B(_1999_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6750_ (.A1(_2650_),
    .A2(_1752_),
    .B(_2843_),
    .C(_2039_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6751_ (.A1(_2715_),
    .A2(_2299_),
    .B(_2844_),
    .C(_1239_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6752_ (.A1(_1620_),
    .A2(_1964_),
    .B(_2061_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _6753_ (.A1(_1620_),
    .A2(_1799_),
    .B1(_2295_),
    .B2(_2777_),
    .C1(_2846_),
    .C2(_1621_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6754_ (.A1(_1176_),
    .A2(_2825_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6755_ (.A1(_1163_),
    .A2(_2848_),
    .B(_1232_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6756_ (.A1(_1163_),
    .A2(_2848_),
    .B(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6757_ (.A1(_2840_),
    .A2(_2845_),
    .A3(_2847_),
    .A4(_2850_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6758_ (.I(_2851_),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6759_ (.I(_0908_),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6760_ (.I(_1642_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6761_ (.A1(_2852_),
    .A2(_2853_),
    .B(_1658_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6762_ (.A1(_2852_),
    .A2(_2853_),
    .B(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6763_ (.A1(_0907_),
    .A2(net170),
    .B(_2308_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6764_ (.A1(_0907_),
    .A2(net170),
    .B(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6765_ (.I(_2365_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6766_ (.I0(_1910_),
    .I1(_2697_),
    .S(_1443_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6767_ (.A1(_1689_),
    .A2(_1907_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6768_ (.A1(_2781_),
    .A2(_2859_),
    .B(_2860_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6769_ (.A1(_1614_),
    .A2(_1603_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6770_ (.A1(_1614_),
    .A2(_1601_),
    .B(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6771_ (.A1(_1598_),
    .A2(_2863_),
    .B(_0905_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6772_ (.A1(_1544_),
    .A2(_2858_),
    .B1(_2861_),
    .B2(_2800_),
    .C(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6773_ (.A1(_2855_),
    .A2(_2857_),
    .A3(_2865_),
    .ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6774_ (.A1(_2852_),
    .A2(_2853_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6775_ (.A1(_1614_),
    .A2(_2866_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6776_ (.A1(_1882_),
    .A2(_2867_),
    .B(_1953_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6777_ (.A1(_1882_),
    .A2(_2867_),
    .B(_2868_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6778_ (.A1(_0864_),
    .A2(_1189_),
    .B(_1232_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6779_ (.A1(_0864_),
    .A2(_1189_),
    .B(_2870_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6780_ (.A1(_1613_),
    .A2(_1964_),
    .B(_1598_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6781_ (.A1(_1613_),
    .A2(_1960_),
    .B1(_2872_),
    .B2(_1615_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6782_ (.A1(_2115_),
    .A2(_2721_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6783_ (.A1(_1971_),
    .A2(_2003_),
    .B(_2874_),
    .C(_1537_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6784_ (.A1(_1246_),
    .A2(_1997_),
    .B(_2875_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6785_ (.A1(_1544_),
    .A2(_2405_),
    .B1(_2876_),
    .B2(_2800_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6786_ (.A1(_2869_),
    .A2(_2871_),
    .A3(_2873_),
    .A4(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6787_ (.I(_2878_),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6788_ (.A1(_1882_),
    .A2(_2852_),
    .A3(_2853_),
    .B(_1616_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6789_ (.A1(_0825_),
    .A2(_2879_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6790_ (.A1(_0825_),
    .A2(net183),
    .B(_2501_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6791_ (.A1(_0825_),
    .A2(net183),
    .B(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6792_ (.A1(_1690_),
    .A2(_2057_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6793_ (.A1(_1999_),
    .A2(_2748_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6794_ (.A1(_2054_),
    .A2(_2053_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6795_ (.A1(_1791_),
    .A2(_2884_),
    .A3(_2885_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6796_ (.A1(_2883_),
    .A2(_2886_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6797_ (.A1(_0822_),
    .A2(_1963_),
    .B(_2060_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6798_ (.I(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6799_ (.A1(_1612_),
    .A2(_1603_),
    .B1(_2889_),
    .B2(_0823_),
    .C(_2505_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6800_ (.A1(_2777_),
    .A2(_2451_),
    .B1(_2887_),
    .B2(_1239_),
    .C(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6801_ (.A1(_2439_),
    .A2(_2880_),
    .B1(_2882_),
    .B2(_2891_),
    .ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6802_ (.A1(net223),
    .A2(_2879_),
    .B(_0822_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6803_ (.A1(_1881_),
    .A2(_2892_),
    .B(_1658_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6804_ (.A1(_1881_),
    .A2(_2892_),
    .B(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6805_ (.A1(_0782_),
    .A2(_1199_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6806_ (.A1(_0782_),
    .A2(_1199_),
    .B(_2308_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6807_ (.I0(_2117_),
    .I1(_2763_),
    .S(_2103_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6808_ (.A1(_1246_),
    .A2(_2116_),
    .B1(_2897_),
    .B2(_2781_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6809_ (.A1(_1611_),
    .A2(_2554_),
    .B(_1597_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6810_ (.I(_0780_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6811_ (.A1(_1611_),
    .A2(_2216_),
    .B1(_2899_),
    .B2(_2900_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6812_ (.A1(_1795_),
    .A2(_2481_),
    .B(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6813_ (.A1(_2895_),
    .A2(_2896_),
    .B1(_2898_),
    .B2(_2800_),
    .C(_2902_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _6814_ (.A1(_2894_),
    .A2(_2903_),
    .ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6815_ (.I(_0724_),
    .Z(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6816_ (.A1(_2904_),
    .A2(_1646_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6817_ (.A1(_2904_),
    .A2(net182),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6818_ (.A1(_2904_),
    .A2(net182),
    .B(_1683_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6819_ (.A1(_2264_),
    .A2(_2785_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6820_ (.A1(_1702_),
    .A2(_2161_),
    .B(_2908_),
    .C(_1754_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6821_ (.A1(_1690_),
    .A2(_2159_),
    .B(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6822_ (.I(_0721_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6823_ (.A1(_2911_),
    .A2(_1602_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6824_ (.A1(_2911_),
    .A2(_2062_),
    .B(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6825_ (.A1(_1803_),
    .A2(_2913_),
    .B(_0722_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6826_ (.A1(_1543_),
    .A2(_2542_),
    .B(_2914_),
    .C(_1812_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6827_ (.A1(_2906_),
    .A2(_2907_),
    .B1(_2910_),
    .B2(_1686_),
    .C(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6828_ (.A1(_2506_),
    .A2(_2905_),
    .B(_2916_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6829_ (.I(_2917_),
    .ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6830_ (.I(_0670_),
    .Z(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6831_ (.A1(_2918_),
    .A2(_1207_),
    .B(_1683_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6832_ (.A1(_2918_),
    .A2(_1207_),
    .B(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6833_ (.A1(_2904_),
    .A2(_1646_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6834_ (.A1(_2918_),
    .A2(_2911_),
    .A3(_2921_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6835_ (.A1(_2911_),
    .A2(_2921_),
    .B(_2918_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6836_ (.A1(_1813_),
    .A2(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6837_ (.A1(_2169_),
    .A2(_2801_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6838_ (.A1(_2054_),
    .A2(_2213_),
    .B(_2925_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6839_ (.A1(_1690_),
    .A2(_2212_),
    .B1(_2926_),
    .B2(_2363_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6840_ (.A1(_1647_),
    .A2(_2554_),
    .B(_2491_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _6841_ (.A1(_1647_),
    .A2(_2302_),
    .B1(_2584_),
    .B2(_1543_),
    .C1(_2928_),
    .C2(_1648_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6842_ (.A1(_2922_),
    .A2(_2924_),
    .B1(_2927_),
    .B2(_1686_),
    .C(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6843_ (.A1(_2920_),
    .A2(_2930_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6844_ (.I(_2931_),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6845_ (.A1(_0808_),
    .A2(_1030_),
    .A3(_0759_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6846_ (.A1(net4),
    .A2(_2714_),
    .Z(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6847_ (.A1(_0487_),
    .A2(_2932_),
    .B1(_2933_),
    .B2(_1223_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6848_ (.A1(net12),
    .A2(net1),
    .A3(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6849_ (.I(_2935_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6850_ (.I(_2936_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6851_ (.I(net65),
    .Z(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6852_ (.A1(_2938_),
    .A2(_0992_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6853_ (.A1(_0808_),
    .A2(_1030_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6854_ (.A1(_0757_),
    .A2(_0758_),
    .A3(_2940_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6855_ (.I(_2941_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6856_ (.A1(_0487_),
    .A2(net12),
    .A3(net1),
    .A4(_2942_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _6857_ (.A1(_2935_),
    .A2(_2943_),
    .Z(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6858_ (.I(_2944_),
    .Z(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6859_ (.I(_2945_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6860_ (.A1(_2938_),
    .A2(_2946_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6861_ (.A1(_2937_),
    .A2(_2939_),
    .B(_2947_),
    .ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6862_ (.I(_2943_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6863_ (.I(_2948_),
    .Z(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6864_ (.I(net76),
    .Z(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6865_ (.I(net208),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6866_ (.A1(_2938_),
    .A2(_0992_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6867_ (.A1(_2950_),
    .A2(_2951_),
    .A3(_2952_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6868_ (.I(_2936_),
    .Z(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6869_ (.I(_2945_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6870_ (.A1(_2950_),
    .A2(_2955_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6871_ (.A1(_2744_),
    .A2(_2949_),
    .B1(_2953_),
    .B2(_2954_),
    .C(_2956_),
    .ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6872_ (.I(net87),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6873_ (.I(_2957_),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6874_ (.A1(_2935_),
    .A2(_2948_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6875_ (.I(_2959_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6876_ (.I(_2960_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6877_ (.A1(net76),
    .A2(_2951_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6878_ (.A1(_2950_),
    .A2(_2951_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6879_ (.A1(_2952_),
    .A2(_2962_),
    .B(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6880_ (.A1(_2958_),
    .A2(_1044_),
    .A3(_2964_),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6881_ (.I(_2932_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _6882_ (.I(_2966_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6883_ (.A1(net12),
    .A2(net1),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6884_ (.A1(_0554_),
    .A2(_2967_),
    .A3(_2968_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6885_ (.I(_2969_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6886_ (.I(_2970_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6887_ (.A1(net119),
    .A2(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6888_ (.A1(_2958_),
    .A2(_2961_),
    .B1(_2965_),
    .B2(_2954_),
    .C(_2972_),
    .ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6889_ (.I(net90),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6890_ (.A1(_2958_),
    .A2(_2973_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6891_ (.I(_0913_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6892_ (.A1(_2957_),
    .A2(_0938_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6893_ (.A1(_2957_),
    .A2(_0938_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6894_ (.A1(_2976_),
    .A2(_2964_),
    .B(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6895_ (.A1(_2973_),
    .A2(_2975_),
    .A3(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6896_ (.I(_2936_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6897_ (.I(_2970_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6898_ (.A1(net122),
    .A2(_2981_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6899_ (.A1(_2961_),
    .A2(_2974_),
    .B1(_2979_),
    .B2(_2980_),
    .C(_2982_),
    .ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6900_ (.I(net91),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6901_ (.A1(net90),
    .A2(_2975_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6902_ (.A1(_2973_),
    .A2(_2975_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6903_ (.A1(_2984_),
    .A2(_2978_),
    .B(_2985_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6904_ (.A1(_2983_),
    .A2(_1166_),
    .A3(_2986_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6905_ (.I(_2945_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6906_ (.A1(_2957_),
    .A2(_2973_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6907_ (.A1(_2983_),
    .A2(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6908_ (.A1(_2988_),
    .A2(_2990_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6909_ (.A1(_2799_),
    .A2(_2949_),
    .B1(_2987_),
    .B2(_2980_),
    .C(_2991_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6910_ (.I(net92),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6911_ (.A1(net87),
    .A2(net90),
    .A3(net91),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6912_ (.A1(_2992_),
    .A2(_2993_),
    .Z(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6913_ (.A1(_2983_),
    .A2(_1059_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6914_ (.A1(_2983_),
    .A2(_1059_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6915_ (.A1(_2995_),
    .A2(_2986_),
    .B(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6916_ (.A1(_2992_),
    .A2(_1124_),
    .A3(_2997_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6917_ (.A1(net124),
    .A2(_2981_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6918_ (.A1(_2961_),
    .A2(_2994_),
    .B1(_2998_),
    .B2(_2980_),
    .C(_2999_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6919_ (.I(_2935_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6920_ (.I(_3000_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6921_ (.I(net93),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6922_ (.A1(_3002_),
    .A2(_1098_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6923_ (.A1(_2992_),
    .A2(_1124_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6924_ (.A1(_2992_),
    .A2(_1124_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6925_ (.A1(_3004_),
    .A2(_2997_),
    .B(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6926_ (.A1(_3003_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6927_ (.A1(net125),
    .A2(_2971_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6928_ (.I(net92),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6929_ (.A1(_3009_),
    .A2(_2993_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6930_ (.A1(_3002_),
    .A2(_3010_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6931_ (.A1(_2946_),
    .A2(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6932_ (.A1(_3001_),
    .A2(_3007_),
    .B(_3008_),
    .C(_3012_),
    .ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6933_ (.I(_2959_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6934_ (.A1(net94),
    .A2(net93),
    .A3(_3010_),
    .Z(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6935_ (.I(net94),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6936_ (.A1(_3002_),
    .A2(_3010_),
    .B(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6937_ (.A1(_3014_),
    .A2(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6938_ (.A1(_3002_),
    .A2(_1098_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6939_ (.A1(_3003_),
    .A2(_3006_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6940_ (.A1(_3018_),
    .A2(_3019_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6941_ (.A1(_3015_),
    .A2(_1148_),
    .A3(_3020_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6942_ (.A1(net126),
    .A2(_2981_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6943_ (.A1(_3013_),
    .A2(_3017_),
    .B1(_3021_),
    .B2(_2980_),
    .C(_3022_),
    .ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6944_ (.I(net95),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6945_ (.A1(_3023_),
    .A2(_3014_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6946_ (.A1(_3023_),
    .A2(_0883_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6947_ (.A1(_3015_),
    .A2(_1149_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6948_ (.I(_3015_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6949_ (.A1(_3027_),
    .A2(_1148_),
    .B(_3018_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6950_ (.A1(_3003_),
    .A2(_3006_),
    .B(_3028_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6951_ (.A1(_3026_),
    .A2(_3029_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6952_ (.A1(_3025_),
    .A2(_3030_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6953_ (.I(_3000_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6954_ (.A1(net127),
    .A2(_2981_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6955_ (.A1(_3013_),
    .A2(_3024_),
    .B1(_3031_),
    .B2(_3032_),
    .C(_3033_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6956_ (.A1(_3023_),
    .A2(_3014_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6957_ (.A1(_0826_),
    .A2(_3034_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6958_ (.A1(_0826_),
    .A2(_0845_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6959_ (.A1(_0826_),
    .A2(_0845_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6960_ (.A1(_3036_),
    .A2(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6961_ (.A1(_3023_),
    .A2(_0884_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6962_ (.A1(_3026_),
    .A2(_3025_),
    .A3(_3029_),
    .B(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6963_ (.A1(_3038_),
    .A2(_3040_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6964_ (.I(_2970_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6965_ (.A1(net128),
    .A2(_3042_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6966_ (.A1(_3013_),
    .A2(_3035_),
    .B1(_3041_),
    .B2(_3032_),
    .C(_3043_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6967_ (.I(_0811_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6968_ (.A1(net66),
    .A2(_3044_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6969_ (.A1(_3039_),
    .A2(_3036_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6970_ (.A1(_3026_),
    .A2(_3025_),
    .A3(_3029_),
    .B(_3046_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6971_ (.A1(_3037_),
    .A2(_3045_),
    .A3(_3047_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6972_ (.A1(_3037_),
    .A2(_3047_),
    .B(_3045_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6973_ (.A1(_3048_),
    .A2(_3049_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6974_ (.A1(net98),
    .A2(_2971_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6975_ (.I(net66),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6976_ (.A1(net96),
    .A2(net95),
    .A3(_3014_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6977_ (.A1(_3052_),
    .A2(_3053_),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6978_ (.A1(_2946_),
    .A2(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6979_ (.A1(_3001_),
    .A2(_3050_),
    .B(_3051_),
    .C(_3055_),
    .ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6980_ (.A1(net67),
    .A2(net66),
    .A3(_3053_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6981_ (.I(net67),
    .Z(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6982_ (.I(_3057_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6983_ (.A1(_3052_),
    .A2(_3053_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6984_ (.A1(_3058_),
    .A2(_3059_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6985_ (.A1(_3056_),
    .A2(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6986_ (.I(_0761_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6987_ (.A1(_3052_),
    .A2(_3044_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6988_ (.A1(_3037_),
    .A2(_3045_),
    .A3(_3047_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6989_ (.A1(_3063_),
    .A2(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6990_ (.A1(_3058_),
    .A2(_3062_),
    .A3(_3065_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6991_ (.A1(net99),
    .A2(_3042_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6992_ (.A1(_3013_),
    .A2(_3061_),
    .B1(_3066_),
    .B2(_3032_),
    .C(_3067_),
    .ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6993_ (.A1(_0671_),
    .A2(_0701_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6994_ (.A1(_3057_),
    .A2(_0761_),
    .B1(_3044_),
    .B2(_3052_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6995_ (.A1(_3057_),
    .A2(_3062_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6996_ (.A1(_3064_),
    .A2(_3069_),
    .B(_3070_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6997_ (.A1(_3068_),
    .A2(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6998_ (.I(net68),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6999_ (.A1(_3073_),
    .A2(_3056_),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7000_ (.A1(_2988_),
    .A2(_3074_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7001_ (.A1(_2917_),
    .A2(_2949_),
    .B1(_3072_),
    .B2(_3032_),
    .C(_3075_),
    .ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7002_ (.I(_3000_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7003_ (.I(net69),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7004_ (.I(_0643_),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7005_ (.A1(_3077_),
    .A2(_3078_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7006_ (.A1(_0671_),
    .A2(_0701_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7007_ (.A1(_3068_),
    .A2(_3071_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7008_ (.A1(_3080_),
    .A2(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7009_ (.A1(_3079_),
    .A2(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7010_ (.A1(net101),
    .A2(_2971_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7011_ (.A1(_3073_),
    .A2(_3056_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7012_ (.A1(_3077_),
    .A2(_3085_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7013_ (.A1(_2946_),
    .A2(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7014_ (.A1(_3076_),
    .A2(_3083_),
    .B(_3084_),
    .C(_3087_),
    .ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7015_ (.I(net70),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7016_ (.A1(net69),
    .A2(_3085_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7017_ (.A1(_3088_),
    .A2(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7018_ (.I(_0561_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7019_ (.A1(net70),
    .A2(_3091_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7020_ (.I(_3069_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7021_ (.A1(_3068_),
    .A2(_3079_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7022_ (.A1(_3057_),
    .A2(_3062_),
    .B1(_3048_),
    .B2(_3093_),
    .C(_3094_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7023_ (.A1(_3077_),
    .A2(_3078_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7024_ (.A1(_3077_),
    .A2(_3078_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7025_ (.A1(_3080_),
    .A2(_3096_),
    .B(_3097_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7026_ (.I(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7027_ (.A1(_3095_),
    .A2(_3099_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7028_ (.A1(_3092_),
    .A2(_3100_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7029_ (.I(_3000_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7030_ (.A1(net102),
    .A2(_3042_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7031_ (.A1(_2960_),
    .A2(_3090_),
    .B1(_3101_),
    .B2(_3102_),
    .C(_3103_),
    .ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7032_ (.I(net71),
    .Z(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7033_ (.I(_1663_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7034_ (.A1(_3104_),
    .A2(_3105_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7035_ (.I(_3092_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7036_ (.A1(_3107_),
    .A2(_3100_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7037_ (.A1(_3088_),
    .A2(_3091_),
    .B(_3108_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7038_ (.A1(_3106_),
    .A2(_3109_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7039_ (.A1(net71),
    .A2(net70),
    .A3(_3089_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7040_ (.A1(_3088_),
    .A2(_3089_),
    .B(_3104_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7041_ (.A1(_3111_),
    .A2(_3112_),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7042_ (.A1(net103),
    .A2(_3042_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7043_ (.A1(_3076_),
    .A2(_3110_),
    .B1(_3113_),
    .B2(_2961_),
    .C(_3114_),
    .ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7044_ (.I(net72),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7045_ (.A1(_3115_),
    .A2(_1820_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7046_ (.A1(_3092_),
    .A2(_3106_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7047_ (.A1(_3095_),
    .A2(_3099_),
    .B(_3117_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7048_ (.A1(_3104_),
    .A2(_3105_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7049_ (.A1(_3104_),
    .A2(_3105_),
    .B(_3091_),
    .C(_3088_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7050_ (.A1(_3119_),
    .A2(_3120_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7051_ (.A1(_3118_),
    .A2(_3121_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7052_ (.A1(_3116_),
    .A2(_3122_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7053_ (.A1(_3115_),
    .A2(_3111_),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7054_ (.A1(_2988_),
    .A2(_3124_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7055_ (.A1(_1935_),
    .A2(_2949_),
    .B1(_3123_),
    .B2(_3102_),
    .C(_3125_),
    .ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7056_ (.I(net73),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7057_ (.A1(_3115_),
    .A2(_3111_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7058_ (.A1(_3126_),
    .A2(_3127_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7059_ (.A1(_3126_),
    .A2(_1936_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7060_ (.A1(_3126_),
    .A2(_1936_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7061_ (.A1(_3129_),
    .A2(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7062_ (.A1(_3115_),
    .A2(_1820_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7063_ (.A1(_3118_),
    .A2(_3121_),
    .B(_3116_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7064_ (.A1(_3132_),
    .A2(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7065_ (.A1(_3131_),
    .A2(_3134_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7066_ (.I(_2969_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7067_ (.A1(net105),
    .A2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7068_ (.A1(_2960_),
    .A2(_3128_),
    .B1(_3135_),
    .B2(_3102_),
    .C(_3137_),
    .ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7069_ (.I(net74),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7070_ (.I(_2010_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7071_ (.A1(_3138_),
    .A2(_3139_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7072_ (.A1(_3132_),
    .A2(_3133_),
    .A3(_3129_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7073_ (.A1(_3130_),
    .A2(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7074_ (.A1(_3140_),
    .A2(_3142_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7075_ (.I(_3138_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7076_ (.A1(_3126_),
    .A2(net72),
    .A3(_3111_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7077_ (.A1(_3144_),
    .A2(_3145_),
    .Z(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7078_ (.A1(net106),
    .A2(_3136_),
    .B1(_2955_),
    .B2(_3146_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7079_ (.A1(_2937_),
    .A2(_3143_),
    .B(_3147_),
    .ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7080_ (.I(net75),
    .Z(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7081_ (.I(_2071_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7082_ (.A1(_3148_),
    .A2(_3149_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7083_ (.I(_3140_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7084_ (.A1(_3151_),
    .A2(_3142_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7085_ (.A1(_3138_),
    .A2(_3139_),
    .B(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7086_ (.A1(_3150_),
    .A2(_3153_),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7087_ (.A1(_3144_),
    .A2(_3145_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7088_ (.A1(_3148_),
    .A2(_3155_),
    .Z(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7089_ (.A1(net107),
    .A2(_3136_),
    .B1(_2955_),
    .B2(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7090_ (.A1(_2937_),
    .A2(_3154_),
    .B(_3157_),
    .ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7091_ (.I(_2127_),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7092_ (.A1(_1741_),
    .A2(_3158_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7093_ (.A1(_3140_),
    .A2(_3150_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7094_ (.I(_3160_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7095_ (.A1(_3116_),
    .A2(_3129_),
    .A3(_3130_),
    .A4(_3161_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7096_ (.A1(_3132_),
    .A2(_3129_),
    .B(_3160_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7097_ (.A1(_3148_),
    .A2(_3149_),
    .B(_3139_),
    .C(_3138_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7098_ (.I(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7099_ (.A1(_3148_),
    .A2(_3149_),
    .B1(_3130_),
    .B2(_3163_),
    .C(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7100_ (.A1(_3122_),
    .A2(_3162_),
    .B(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7101_ (.A1(_3159_),
    .A2(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7102_ (.I(_1741_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7103_ (.A1(net75),
    .A2(_3155_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7104_ (.A1(_3169_),
    .A2(_3170_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7105_ (.A1(_2988_),
    .A2(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7106_ (.A1(_2181_),
    .A2(_2948_),
    .B1(_3168_),
    .B2(_3102_),
    .C(_3172_),
    .ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7107_ (.I(net78),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7108_ (.I(_2183_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7109_ (.A1(_3173_),
    .A2(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7110_ (.A1(_3173_),
    .A2(_3174_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7111_ (.A1(_3175_),
    .A2(_3176_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7112_ (.A1(_3169_),
    .A2(_3158_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7113_ (.A1(_3159_),
    .A2(_3167_),
    .B(_3178_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7114_ (.A1(_3177_),
    .A2(_3179_),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7115_ (.A1(net78),
    .A2(_1741_),
    .A3(_3170_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7116_ (.A1(_3169_),
    .A2(_3170_),
    .B(_3173_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7117_ (.A1(_3181_),
    .A2(_3182_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7118_ (.A1(_2955_),
    .A2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7119_ (.A1(_2222_),
    .A2(_2948_),
    .B1(_3180_),
    .B2(_3001_),
    .C(_3184_),
    .ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7120_ (.I(net79),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7121_ (.A1(_3185_),
    .A2(_2224_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7122_ (.I(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7123_ (.A1(_3173_),
    .A2(_3174_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7124_ (.A1(_3175_),
    .A2(_3179_),
    .B(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7125_ (.A1(_3187_),
    .A2(_3189_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7126_ (.I(_2969_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7127_ (.I(_2944_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7128_ (.A1(_3185_),
    .A2(_3181_),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7129_ (.A1(net111),
    .A2(_3191_),
    .B1(_3192_),
    .B2(_3193_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7130_ (.A1(_2937_),
    .A2(_3190_),
    .B(_3194_),
    .ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7131_ (.I(net80),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7132_ (.I(_2273_),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7133_ (.A1(_3195_),
    .A2(_3196_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7134_ (.I(_3197_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7135_ (.A1(_3185_),
    .A2(_2224_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7136_ (.A1(_3186_),
    .A2(_3189_),
    .B(_3199_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7137_ (.A1(_3198_),
    .A2(_3200_),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7138_ (.A1(_3198_),
    .A2(_3200_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7139_ (.I(_2969_),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7140_ (.I(_2944_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7141_ (.A1(_3185_),
    .A2(_3181_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7142_ (.A1(_3195_),
    .A2(_3205_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7143_ (.A1(net112),
    .A2(_3203_),
    .B1(_3204_),
    .B2(_3206_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7144_ (.A1(_3076_),
    .A2(_3201_),
    .A3(_3202_),
    .B(_3207_),
    .ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7145_ (.I(net81),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7146_ (.A1(net80),
    .A2(net79),
    .A3(_3181_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7147_ (.A1(_3208_),
    .A2(_3209_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7148_ (.A1(_3208_),
    .A2(_2314_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7149_ (.A1(_3159_),
    .A2(_3177_),
    .A3(_3186_),
    .A4(_3197_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7150_ (.A1(_3162_),
    .A2(_3212_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7151_ (.I(_3213_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7152_ (.A1(_3118_),
    .A2(_3121_),
    .B(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7153_ (.A1(_3169_),
    .A2(_3158_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7154_ (.A1(_3216_),
    .A2(_3175_),
    .B(_3187_),
    .C(_3198_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7155_ (.A1(_3195_),
    .A2(_3196_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7156_ (.A1(_3195_),
    .A2(_3196_),
    .B(_3199_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7157_ (.A1(_3218_),
    .A2(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7158_ (.A1(_3166_),
    .A2(_3212_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7159_ (.A1(_3176_),
    .A2(_3217_),
    .B(_3220_),
    .C(_3221_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7160_ (.A1(_3215_),
    .A2(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7161_ (.A1(_3211_),
    .A2(_3223_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7162_ (.A1(net113),
    .A2(_3136_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7163_ (.A1(_2960_),
    .A2(_3210_),
    .B1(_3224_),
    .B2(_3001_),
    .C(_3225_),
    .ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7164_ (.I(_2936_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7165_ (.I(net82),
    .Z(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7166_ (.I(_2377_),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7167_ (.A1(_3227_),
    .A2(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7168_ (.A1(_3227_),
    .A2(_3228_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7169_ (.A1(_3229_),
    .A2(_3230_),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7170_ (.I(_3208_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7171_ (.A1(_3232_),
    .A2(_2312_),
    .A3(_2313_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7172_ (.A1(_3211_),
    .A2(_3223_),
    .B(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7173_ (.A1(_3231_),
    .A2(_3234_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7174_ (.A1(_3232_),
    .A2(_3209_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7175_ (.A1(_3227_),
    .A2(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7176_ (.A1(net114),
    .A2(_3191_),
    .B1(_3192_),
    .B2(_3237_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7177_ (.A1(_3226_),
    .A2(_3235_),
    .B(_3238_),
    .ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7178_ (.I(net83),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7179_ (.A1(_3239_),
    .A2(_2420_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7180_ (.A1(_3227_),
    .A2(_3228_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7181_ (.A1(_3229_),
    .A2(_3234_),
    .B(_3241_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7182_ (.A1(_3240_),
    .A2(_3242_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7183_ (.A1(net82),
    .A2(_3236_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7184_ (.A1(_3239_),
    .A2(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7185_ (.A1(net115),
    .A2(_3191_),
    .B1(_3192_),
    .B2(_3245_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7186_ (.A1(_3226_),
    .A2(_3243_),
    .B(_3246_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7187_ (.I(net84),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7188_ (.I(_2464_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7189_ (.A1(_3247_),
    .A2(_3248_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7190_ (.A1(_3239_),
    .A2(_2420_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7191_ (.I(_3250_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7192_ (.A1(_3240_),
    .A2(_3242_),
    .B(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7193_ (.A1(_3249_),
    .A2(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7194_ (.A1(net84),
    .A2(net83),
    .A3(_3244_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7195_ (.I(_3254_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7196_ (.A1(_3239_),
    .A2(_3244_),
    .B(_3247_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7197_ (.A1(_3255_),
    .A2(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7198_ (.A1(net116),
    .A2(_3191_),
    .B1(_3192_),
    .B2(_3257_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7199_ (.A1(_3226_),
    .A2(_3253_),
    .B(_3258_),
    .ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7200_ (.I(net85),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7201_ (.A1(_3259_),
    .A2(_2508_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7202_ (.A1(_3259_),
    .A2(_2508_),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7203_ (.A1(_3260_),
    .A2(_3261_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7204_ (.A1(_3240_),
    .A2(_3249_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7205_ (.A1(_3211_),
    .A2(_3231_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7206_ (.A1(_3215_),
    .A2(_3222_),
    .B(_3263_),
    .C(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7207_ (.A1(_3208_),
    .A2(_2314_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7208_ (.A1(_3266_),
    .A2(_3229_),
    .B(_3263_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7209_ (.A1(_3247_),
    .A2(_3248_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7210_ (.A1(_3250_),
    .A2(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7211_ (.A1(_3247_),
    .A2(_3248_),
    .B1(_3230_),
    .B2(_3267_),
    .C(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7212_ (.I(_3270_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7213_ (.A1(_3265_),
    .A2(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7214_ (.A1(_3262_),
    .A2(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7215_ (.A1(_3259_),
    .A2(_3255_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7216_ (.A1(net117),
    .A2(_3203_),
    .B1(_3204_),
    .B2(_3274_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7217_ (.A1(_3226_),
    .A2(_3273_),
    .B(_3275_),
    .ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7218_ (.I(net86),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7219_ (.A1(_3276_),
    .A2(_2560_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7220_ (.I(_3277_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7221_ (.A1(_3276_),
    .A2(_2560_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7222_ (.A1(_3278_),
    .A2(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7223_ (.A1(_3265_),
    .A2(_3271_),
    .B(_3261_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7224_ (.A1(_3260_),
    .A2(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7225_ (.A1(_3280_),
    .A2(_3282_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7226_ (.A1(net85),
    .A2(_3255_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7227_ (.A1(_3276_),
    .A2(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7228_ (.A1(net118),
    .A2(_3203_),
    .B1(_3204_),
    .B2(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7229_ (.A1(_2954_),
    .A2(_3283_),
    .B(_3286_),
    .ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7230_ (.I(net88),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7231_ (.A1(_3287_),
    .A2(_2600_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7232_ (.A1(_3260_),
    .A2(_3281_),
    .B(_3278_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7233_ (.A1(_3279_),
    .A2(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7234_ (.A1(_3288_),
    .A2(_3290_),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7235_ (.A1(net86),
    .A2(net85),
    .A3(_3254_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7236_ (.A1(_3287_),
    .A2(_3292_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7237_ (.A1(net120),
    .A2(_3203_),
    .B1(_3204_),
    .B2(_3293_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7238_ (.A1(_2954_),
    .A2(_3291_),
    .B(_3294_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7239_ (.A1(_3287_),
    .A2(_2600_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7240_ (.A1(_3279_),
    .A2(_3289_),
    .B(_3288_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7241_ (.A1(_0747_),
    .A2(net89),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7242_ (.A1(_3295_),
    .A2(_3296_),
    .A3(_3297_),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7243_ (.A1(_3295_),
    .A2(_3296_),
    .B(_3297_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7244_ (.A1(_3276_),
    .A2(_3259_),
    .A3(_3287_),
    .A4(_3255_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7245_ (.A1(net89),
    .A2(_3300_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7246_ (.I(_3301_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7247_ (.A1(net121),
    .A2(_2970_),
    .B1(_2945_),
    .B2(_3302_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7248_ (.A1(_3076_),
    .A2(_3298_),
    .A3(_3299_),
    .B(_3303_),
    .ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7249_ (.A1(_0554_),
    .A2(_0551_),
    .A3(_0480_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7250_ (.A1(_2940_),
    .A2(_3304_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7251_ (.I(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7252_ (.I(_3306_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7253_ (.I(_1214_),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7254_ (.I(_3308_),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7255_ (.I(_2941_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7256_ (.I(_3305_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7257_ (.A1(net33),
    .A2(_3309_),
    .B1(_3310_),
    .B2(_2938_),
    .C(_3311_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7258_ (.A1(_1214_),
    .A2(_2941_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7259_ (.I(_3313_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7260_ (.I(_3314_),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7261_ (.A1(_0992_),
    .A2(_3315_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7262_ (.A1(_2714_),
    .A2(_3307_),
    .B1(_3312_),
    .B2(_3316_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7263_ (.I(_3317_),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7264_ (.I(_3318_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _7265_ (.I(net31),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7266_ (.I(net30),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7267_ (.I(net32),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7268_ (.I(_3304_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7269_ (.A1(_3313_),
    .A2(_3323_),
    .B(net3),
    .C(_2968_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7270_ (.A1(net2),
    .A2(_3322_),
    .A3(_3324_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _7271_ (.A1(_3320_),
    .A2(_3321_),
    .A3(_3325_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7272_ (.I(_3326_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7273_ (.I(_3327_),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7274_ (.I0(\reg_file.reg_storage[14][0] ),
    .I1(_3319_),
    .S(_3328_),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7275_ (.I(_3329_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7276_ (.A1(_2951_),
    .A2(_3315_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7277_ (.I(_3308_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7278_ (.I(_3305_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7279_ (.I(_3332_),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7280_ (.A1(net44),
    .A2(_3331_),
    .B1(_3310_),
    .B2(_2950_),
    .C(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7281_ (.A1(_2744_),
    .A2(_3307_),
    .B1(_3330_),
    .B2(_3334_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7282_ (.I(_3335_),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7283_ (.I(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7284_ (.I0(\reg_file.reg_storage[14][1] ),
    .I1(_3337_),
    .S(_3328_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7285_ (.I(_3338_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7286_ (.I(_3326_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7287_ (.I(_3339_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7288_ (.I(_3340_),
    .Z(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7289_ (.A1(_2940_),
    .A2(_3304_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7290_ (.I(_3342_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7291_ (.I(_3343_),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7292_ (.I(_1214_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7293_ (.I(_3345_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7294_ (.I(_3314_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7295_ (.I(_3342_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7296_ (.A1(_2958_),
    .A2(_2966_),
    .B(_3348_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7297_ (.A1(net55),
    .A2(_3346_),
    .B1(_0938_),
    .B2(_3347_),
    .C(_3349_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7298_ (.I(_3350_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7299_ (.A1(net119),
    .A2(_3344_),
    .B(_3351_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7300_ (.I(_3352_),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7301_ (.I(_3326_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7302_ (.I(_3354_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7303_ (.A1(\reg_file.reg_storage[14][2] ),
    .A2(_3355_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7304_ (.A1(_3341_),
    .A2(_3353_),
    .B(_3356_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7305_ (.I(_3342_),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7306_ (.A1(_2975_),
    .A2(_3347_),
    .A3(_3357_),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7307_ (.I(_3345_),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7308_ (.A1(net58),
    .A2(_3359_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7309_ (.A1(_2967_),
    .A2(_2974_),
    .B(_3357_),
    .C(_3360_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _7310_ (.A1(net122),
    .A2(_3357_),
    .B1(_3358_),
    .B2(_3361_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7311_ (.I(_3362_),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7312_ (.A1(\reg_file.reg_storage[14][3] ),
    .A2(_3355_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7313_ (.A1(_3341_),
    .A2(_3363_),
    .B(_3364_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7314_ (.A1(_1059_),
    .A2(_3315_),
    .A3(_3348_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7315_ (.A1(net59),
    .A2(_3331_),
    .B1(_3310_),
    .B2(_2990_),
    .C(_3333_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7316_ (.A1(net166),
    .A2(_3307_),
    .B1(_3365_),
    .B2(_3366_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7317_ (.I(_3367_),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7318_ (.I(_3368_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7319_ (.I0(\reg_file.reg_storage[14][4] ),
    .I1(_3369_),
    .S(_3328_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7320_ (.I(_3370_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7321_ (.A1(_3315_),
    .A2(_3348_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7322_ (.I(_3332_),
    .Z(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7323_ (.A1(net60),
    .A2(_3331_),
    .B(_3372_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7324_ (.A1(_2967_),
    .A2(_2994_),
    .B1(_3371_),
    .B2(_1123_),
    .C(_3373_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7325_ (.A1(net124),
    .A2(_3344_),
    .B(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7326_ (.I(_3375_),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7327_ (.I(_3327_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7328_ (.A1(\reg_file.reg_storage[14][5] ),
    .A2(_3377_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7329_ (.A1(_3341_),
    .A2(_3376_),
    .B(_3378_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7330_ (.I(_2942_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7331_ (.A1(_3379_),
    .A2(_3011_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7332_ (.I(_3332_),
    .Z(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7333_ (.A1(net61),
    .A2(_3346_),
    .B1(_1098_),
    .B2(_3347_),
    .C(_3381_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7334_ (.A1(_3380_),
    .A2(_3382_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7335_ (.A1(net125),
    .A2(_3344_),
    .B(_3383_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7336_ (.I(_3384_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7337_ (.A1(\reg_file.reg_storage[14][6] ),
    .A2(_3377_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7338_ (.A1(_3341_),
    .A2(_3385_),
    .B(_3386_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7339_ (.I(_3340_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7340_ (.I(_2966_),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7341_ (.I(_3345_),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7342_ (.I(_3313_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7343_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7344_ (.A1(net62),
    .A2(_3389_),
    .B1(_1149_),
    .B2(_3391_),
    .C(_3372_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7345_ (.A1(_3388_),
    .A2(_3017_),
    .B(_3392_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7346_ (.A1(net126),
    .A2(_3344_),
    .B(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7347_ (.I(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7348_ (.A1(\reg_file.reg_storage[14][7] ),
    .A2(_3377_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7349_ (.A1(_3387_),
    .A2(_3395_),
    .B(_3396_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7350_ (.I(_3343_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7351_ (.A1(net63),
    .A2(_3389_),
    .B1(_0884_),
    .B2(_3391_),
    .C(_3372_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7352_ (.A1(_3388_),
    .A2(_3024_),
    .B(_3398_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7353_ (.A1(net127),
    .A2(_3397_),
    .B(_3399_),
    .ZN(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7354_ (.I(_3400_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7355_ (.A1(\reg_file.reg_storage[14][8] ),
    .A2(_3377_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7356_ (.A1(_3387_),
    .A2(_3401_),
    .B(_3402_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7357_ (.A1(net64),
    .A2(_3389_),
    .B1(_0845_),
    .B2(_3391_),
    .C(_3372_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7358_ (.A1(_3388_),
    .A2(_3035_),
    .B(_3403_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7359_ (.A1(net128),
    .A2(_3397_),
    .B(_3404_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7360_ (.I(_3405_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7361_ (.I(_3327_),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7362_ (.A1(\reg_file.reg_storage[14][9] ),
    .A2(_3407_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7363_ (.A1(_3387_),
    .A2(_3406_),
    .B(_3408_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7364_ (.A1(_3379_),
    .A2(_3054_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7365_ (.A1(net34),
    .A2(_3346_),
    .B1(_3044_),
    .B2(_3347_),
    .C(_3381_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7366_ (.A1(_3409_),
    .A2(_3410_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7367_ (.A1(net98),
    .A2(_3397_),
    .B(_3411_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7368_ (.I(_3412_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7369_ (.A1(\reg_file.reg_storage[14][10] ),
    .A2(_3407_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7370_ (.A1(_3387_),
    .A2(_3413_),
    .B(_3414_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7371_ (.I(_3354_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7372_ (.I(_3332_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7373_ (.A1(net35),
    .A2(_3389_),
    .B1(_3062_),
    .B2(_3391_),
    .C(_3416_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7374_ (.A1(_3388_),
    .A2(_3061_),
    .B(_3417_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7375_ (.A1(net99),
    .A2(_3397_),
    .B(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7376_ (.I(_3419_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7377_ (.A1(\reg_file.reg_storage[14][11] ),
    .A2(_3407_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7378_ (.A1(_3415_),
    .A2(_3420_),
    .B(_3421_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7379_ (.I(_2942_),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7380_ (.A1(_3422_),
    .A2(_3074_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7381_ (.I(_3308_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7382_ (.I(_3390_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7383_ (.I(_3305_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7384_ (.A1(net36),
    .A2(_3424_),
    .B1(_0701_),
    .B2(_3425_),
    .C(_3426_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7385_ (.A1(_2917_),
    .A2(_3307_),
    .B1(_3423_),
    .B2(_3427_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7386_ (.I(_3428_),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7387_ (.I(_3429_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7388_ (.I0(\reg_file.reg_storage[14][12] ),
    .I1(_3430_),
    .S(_3328_),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7389_ (.I(_3431_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7390_ (.I(_3343_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7391_ (.A1(_3379_),
    .A2(_3086_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7392_ (.I(_3314_),
    .Z(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7393_ (.I(_3306_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7394_ (.A1(net37),
    .A2(_3346_),
    .B1(_3078_),
    .B2(_3434_),
    .C(_3435_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7395_ (.A1(_3433_),
    .A2(_3436_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7396_ (.A1(net101),
    .A2(_3432_),
    .B(_3437_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7397_ (.I(_3438_),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7398_ (.A1(\reg_file.reg_storage[14][13] ),
    .A2(_3407_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7399_ (.A1(_3415_),
    .A2(_3439_),
    .B(_3440_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7400_ (.I(_2966_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7401_ (.I(_3308_),
    .Z(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7402_ (.I(_3390_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7403_ (.A1(net38),
    .A2(_3442_),
    .B1(_3091_),
    .B2(_3443_),
    .C(_3416_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7404_ (.A1(_3441_),
    .A2(_3090_),
    .B(_3444_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7405_ (.A1(net102),
    .A2(_3432_),
    .B(_3445_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7406_ (.I(_3446_),
    .Z(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7407_ (.I(_3339_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7408_ (.A1(\reg_file.reg_storage[14][14] ),
    .A2(_3448_),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7409_ (.A1(_3415_),
    .A2(_3447_),
    .B(_3449_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7410_ (.A1(net39),
    .A2(_3442_),
    .B1(_3105_),
    .B2(_3443_),
    .C(_3416_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7411_ (.A1(_3441_),
    .A2(_3113_),
    .B(_3450_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7412_ (.A1(net103),
    .A2(_3432_),
    .B(_3451_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7413_ (.I(_3452_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7414_ (.A1(\reg_file.reg_storage[14][15] ),
    .A2(_3448_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7415_ (.A1(_3415_),
    .A2(_3453_),
    .B(_3454_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7416_ (.I(_3306_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7417_ (.A1(_3422_),
    .A2(_3124_),
    .ZN(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7418_ (.A1(net40),
    .A2(_3424_),
    .B1(_1820_),
    .B2(_3425_),
    .C(_3426_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7419_ (.A1(_1935_),
    .A2(_3455_),
    .B1(_3456_),
    .B2(_3457_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7420_ (.I(_3458_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7421_ (.I(_3459_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _7422_ (.I(_3327_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7423_ (.I0(\reg_file.reg_storage[14][16] ),
    .I1(_3460_),
    .S(_3461_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7424_ (.I(_3462_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7425_ (.I(_3354_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7426_ (.A1(net41),
    .A2(_3442_),
    .B1(_1936_),
    .B2(_3443_),
    .C(_3416_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7427_ (.A1(_3441_),
    .A2(_3128_),
    .B(_3464_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7428_ (.A1(net105),
    .A2(_3432_),
    .B(_3465_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7429_ (.I(_3466_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7430_ (.A1(\reg_file.reg_storage[14][17] ),
    .A2(_3448_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7431_ (.A1(_3463_),
    .A2(_3467_),
    .B(_3468_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7432_ (.I(_3343_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7433_ (.A1(_3379_),
    .A2(_3146_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7434_ (.I(_3345_),
    .Z(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7435_ (.A1(net42),
    .A2(_3471_),
    .B1(_3139_),
    .B2(_3434_),
    .C(_3435_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7436_ (.A1(_3470_),
    .A2(_3472_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7437_ (.A1(net106),
    .A2(_3469_),
    .B(_3473_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7438_ (.I(_3474_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7439_ (.A1(\reg_file.reg_storage[14][18] ),
    .A2(_3448_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7440_ (.A1(_3463_),
    .A2(_3475_),
    .B(_3476_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7441_ (.I(_2942_),
    .Z(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7442_ (.A1(_3477_),
    .A2(_3156_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7443_ (.A1(net43),
    .A2(_3471_),
    .B1(_3149_),
    .B2(_3434_),
    .C(_3435_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7444_ (.A1(_3478_),
    .A2(_3479_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7445_ (.A1(net107),
    .A2(_3469_),
    .B(_3480_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7446_ (.I(_3481_),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7447_ (.I(_3339_),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7448_ (.A1(\reg_file.reg_storage[14][19] ),
    .A2(_3483_),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7449_ (.A1(_3463_),
    .A2(_3482_),
    .B(_3484_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7450_ (.I(_2941_),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7451_ (.A1(_3485_),
    .A2(_3171_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7452_ (.A1(net45),
    .A2(_3424_),
    .B1(_3158_),
    .B2(_3425_),
    .C(_3426_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7453_ (.A1(_2181_),
    .A2(_3455_),
    .B1(_3486_),
    .B2(_3487_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7454_ (.I(_3488_),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7455_ (.I(_3489_),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7456_ (.I0(\reg_file.reg_storage[14][20] ),
    .I1(_3490_),
    .S(_3461_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7457_ (.I(_3491_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7458_ (.A1(_3485_),
    .A2(_3183_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7459_ (.I(_3390_),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7460_ (.A1(net46),
    .A2(_3424_),
    .B1(_3174_),
    .B2(_3493_),
    .C(_3426_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7461_ (.A1(net225),
    .A2(_3455_),
    .B1(_3492_),
    .B2(_3494_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7462_ (.I(_3495_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7463_ (.I(_3496_),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7464_ (.I0(\reg_file.reg_storage[14][21] ),
    .I1(_3497_),
    .S(_3461_),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7465_ (.I(_3498_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7466_ (.I(net111),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7467_ (.A1(_3485_),
    .A2(_3193_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7468_ (.A1(net47),
    .A2(_3309_),
    .B1(_2224_),
    .B2(_3493_),
    .C(_3311_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7469_ (.A1(_3499_),
    .A2(_3455_),
    .B1(_3500_),
    .B2(_3501_),
    .ZN(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7470_ (.I(_3502_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7471_ (.I(_3503_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7472_ (.I0(\reg_file.reg_storage[14][22] ),
    .I1(_3504_),
    .S(_3461_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7473_ (.I(_3505_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7474_ (.A1(_3477_),
    .A2(_3206_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7475_ (.A1(net48),
    .A2(_3471_),
    .B1(_3196_),
    .B2(_3434_),
    .C(_3435_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7476_ (.A1(_3506_),
    .A2(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7477_ (.A1(net112),
    .A2(_3469_),
    .B(_3508_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7478_ (.I(_3509_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7479_ (.A1(\reg_file.reg_storage[14][23] ),
    .A2(_3483_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7480_ (.A1(_3463_),
    .A2(_3510_),
    .B(_3511_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7481_ (.I(_3354_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7482_ (.A1(net49),
    .A2(_3442_),
    .B1(_2314_),
    .B2(_3443_),
    .C(_3333_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7483_ (.A1(_3441_),
    .A2(_3210_),
    .B(_3513_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7484_ (.A1(net113),
    .A2(_3469_),
    .B(_3514_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7485_ (.I(_3515_),
    .Z(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7486_ (.A1(\reg_file.reg_storage[14][24] ),
    .A2(_3483_),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7487_ (.A1(_3512_),
    .A2(_3516_),
    .B(_3517_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7488_ (.I(_3348_),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7489_ (.A1(_3477_),
    .A2(_3237_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7490_ (.I(_3314_),
    .Z(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7491_ (.I(_3306_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7492_ (.A1(net50),
    .A2(_3471_),
    .B1(_3228_),
    .B2(_3520_),
    .C(_3521_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7493_ (.A1(_3519_),
    .A2(_3522_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7494_ (.A1(net114),
    .A2(_3518_),
    .B(_3523_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7495_ (.I(_3524_),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7496_ (.A1(\reg_file.reg_storage[14][25] ),
    .A2(_3483_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7497_ (.A1(_3512_),
    .A2(_3525_),
    .B(_3526_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7498_ (.A1(_3477_),
    .A2(_3245_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7499_ (.A1(net51),
    .A2(_3359_),
    .B1(_2420_),
    .B2(_3520_),
    .C(_3521_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7500_ (.A1(_3527_),
    .A2(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7501_ (.A1(net115),
    .A2(_3518_),
    .B(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7502_ (.I(_3530_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7503_ (.I(_3339_),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7504_ (.A1(\reg_file.reg_storage[14][26] ),
    .A2(_3532_),
    .ZN(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7505_ (.A1(_3512_),
    .A2(_3531_),
    .B(_3533_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7506_ (.A1(_3422_),
    .A2(_3257_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7507_ (.A1(net52),
    .A2(_3359_),
    .B1(_3248_),
    .B2(_3520_),
    .C(_3521_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7508_ (.A1(_3534_),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7509_ (.A1(net116),
    .A2(_3518_),
    .B(_3536_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7510_ (.I(_3537_),
    .Z(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7511_ (.A1(\reg_file.reg_storage[14][27] ),
    .A2(_3532_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7512_ (.A1(_3512_),
    .A2(_3538_),
    .B(_3539_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7513_ (.A1(_3422_),
    .A2(_3274_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7514_ (.A1(net53),
    .A2(_3359_),
    .B1(_2508_),
    .B2(_3520_),
    .C(_3521_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7515_ (.A1(_3540_),
    .A2(_3541_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7516_ (.A1(net117),
    .A2(_3518_),
    .B(_3542_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7517_ (.I(_3543_),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7518_ (.A1(\reg_file.reg_storage[14][28] ),
    .A2(_3532_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7519_ (.A1(_3355_),
    .A2(_3544_),
    .B(_3545_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7520_ (.I(net118),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7521_ (.A1(_3485_),
    .A2(_3285_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7522_ (.A1(net54),
    .A2(_3309_),
    .B1(_2560_),
    .B2(_3493_),
    .C(_3311_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7523_ (.A1(_3546_),
    .A2(_3381_),
    .B1(_3547_),
    .B2(_3548_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7524_ (.I(_3549_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7525_ (.I(_3550_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7526_ (.I0(\reg_file.reg_storage[14][29] ),
    .I1(_3551_),
    .S(_3340_),
    .Z(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7527_ (.I(_3552_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7528_ (.A1(_3310_),
    .A2(_3293_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7529_ (.A1(net56),
    .A2(_3309_),
    .B1(_2600_),
    .B2(_3493_),
    .C(_3311_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _7530_ (.A1(_2634_),
    .A2(_3381_),
    .B1(_3553_),
    .B2(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7531_ (.I(_3555_),
    .Z(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7532_ (.I(_3556_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7533_ (.I0(\reg_file.reg_storage[14][30] ),
    .I1(_3557_),
    .S(_3340_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7534_ (.I(_3558_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7535_ (.A1(net57),
    .A2(_3331_),
    .B1(_3425_),
    .B2(_0746_),
    .C(_3333_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7536_ (.A1(_2967_),
    .A2(_3301_),
    .B(_3559_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7537_ (.A1(net218),
    .A2(_3357_),
    .B(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7538_ (.I(_3561_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7539_ (.A1(\reg_file.reg_storage[14][31] ),
    .A2(_3532_),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7540_ (.A1(_3355_),
    .A2(_3562_),
    .B(_3563_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7541_ (.I(net31),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _7542_ (.I(net30),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _7543_ (.A1(_3564_),
    .A2(_3565_),
    .A3(_3325_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7544_ (.I(_3566_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7545_ (.I(_3567_),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7546_ (.I0(\reg_file.reg_storage[13][0] ),
    .I1(_3319_),
    .S(_3568_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7547_ (.I(_3569_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7548_ (.I0(\reg_file.reg_storage[13][1] ),
    .I1(_3337_),
    .S(_3568_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7549_ (.I(_3570_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7550_ (.I(_3566_),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7551_ (.I(_3571_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7552_ (.I(_3572_),
    .Z(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7553_ (.I(_3566_),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7554_ (.I(_3574_),
    .Z(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7555_ (.A1(\reg_file.reg_storage[13][2] ),
    .A2(_3575_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7556_ (.A1(_3353_),
    .A2(_3573_),
    .B(_3576_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7557_ (.A1(\reg_file.reg_storage[13][3] ),
    .A2(_3575_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7558_ (.A1(_3363_),
    .A2(_3573_),
    .B(_3577_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7559_ (.I0(\reg_file.reg_storage[13][4] ),
    .I1(_3369_),
    .S(_3568_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7560_ (.I(_3578_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7561_ (.I(_3567_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7562_ (.A1(\reg_file.reg_storage[13][5] ),
    .A2(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7563_ (.A1(_3376_),
    .A2(_3573_),
    .B(_3580_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7564_ (.A1(\reg_file.reg_storage[13][6] ),
    .A2(_3579_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7565_ (.A1(_3385_),
    .A2(_3573_),
    .B(_3581_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7566_ (.I(_3572_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7567_ (.A1(\reg_file.reg_storage[13][7] ),
    .A2(_3579_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7568_ (.A1(_3395_),
    .A2(_3582_),
    .B(_3583_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7569_ (.A1(\reg_file.reg_storage[13][8] ),
    .A2(_3579_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7570_ (.A1(_3401_),
    .A2(_3582_),
    .B(_3584_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7571_ (.I(_3567_),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7572_ (.A1(\reg_file.reg_storage[13][9] ),
    .A2(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7573_ (.A1(_3406_),
    .A2(_3582_),
    .B(_3586_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7574_ (.A1(\reg_file.reg_storage[13][10] ),
    .A2(_3585_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7575_ (.A1(_3413_),
    .A2(_3582_),
    .B(_3587_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7576_ (.I(_3572_),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7577_ (.A1(\reg_file.reg_storage[13][11] ),
    .A2(_3585_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7578_ (.A1(_3420_),
    .A2(_3588_),
    .B(_3589_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7579_ (.I(_3567_),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7580_ (.I0(\reg_file.reg_storage[13][12] ),
    .I1(_3430_),
    .S(_3590_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7581_ (.I(_3591_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7582_ (.A1(\reg_file.reg_storage[13][13] ),
    .A2(_3585_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7583_ (.A1(_3439_),
    .A2(_3588_),
    .B(_3592_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7584_ (.I(_3571_),
    .Z(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7585_ (.A1(\reg_file.reg_storage[13][14] ),
    .A2(_3593_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7586_ (.A1(_3447_),
    .A2(_3588_),
    .B(_3594_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7587_ (.A1(\reg_file.reg_storage[13][15] ),
    .A2(_3593_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7588_ (.A1(_3453_),
    .A2(_3588_),
    .B(_3595_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7589_ (.I0(\reg_file.reg_storage[13][16] ),
    .I1(_3460_),
    .S(_3590_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7590_ (.I(_3596_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7591_ (.I(_3572_),
    .Z(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7592_ (.A1(\reg_file.reg_storage[13][17] ),
    .A2(_3593_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7593_ (.A1(_3467_),
    .A2(_3597_),
    .B(_3598_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7594_ (.A1(\reg_file.reg_storage[13][18] ),
    .A2(_3593_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7595_ (.A1(_3475_),
    .A2(_3597_),
    .B(_3599_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7596_ (.I(_3571_),
    .Z(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7597_ (.A1(\reg_file.reg_storage[13][19] ),
    .A2(_3600_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7598_ (.A1(_3482_),
    .A2(_3597_),
    .B(_3601_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7599_ (.I0(\reg_file.reg_storage[13][20] ),
    .I1(_3490_),
    .S(_3590_),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7600_ (.I(_3602_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7601_ (.I0(\reg_file.reg_storage[13][21] ),
    .I1(_3497_),
    .S(_3590_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7602_ (.I(_3603_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7603_ (.I0(\reg_file.reg_storage[13][22] ),
    .I1(_3504_),
    .S(_3574_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7604_ (.I(_3604_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7605_ (.A1(\reg_file.reg_storage[13][23] ),
    .A2(_3600_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7606_ (.A1(_3510_),
    .A2(_3597_),
    .B(_3605_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7607_ (.I(_3568_),
    .Z(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7608_ (.A1(\reg_file.reg_storage[13][24] ),
    .A2(_3600_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7609_ (.A1(_3516_),
    .A2(_3606_),
    .B(_3607_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7610_ (.A1(\reg_file.reg_storage[13][25] ),
    .A2(_3600_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7611_ (.A1(_3525_),
    .A2(_3606_),
    .B(_3608_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7612_ (.I(_3571_),
    .Z(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7613_ (.A1(\reg_file.reg_storage[13][26] ),
    .A2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7614_ (.A1(_3531_),
    .A2(_3606_),
    .B(_3610_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7615_ (.A1(\reg_file.reg_storage[13][27] ),
    .A2(_3609_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7616_ (.A1(_3538_),
    .A2(_3606_),
    .B(_3611_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7617_ (.A1(\reg_file.reg_storage[13][28] ),
    .A2(_3609_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7618_ (.A1(_3544_),
    .A2(_3575_),
    .B(_3612_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7619_ (.I0(\reg_file.reg_storage[13][29] ),
    .I1(_3551_),
    .S(_3574_),
    .Z(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7620_ (.I(_3613_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7621_ (.I0(\reg_file.reg_storage[13][30] ),
    .I1(_3557_),
    .S(_3574_),
    .Z(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7622_ (.I(_3614_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7623_ (.A1(\reg_file.reg_storage[13][31] ),
    .A2(_3609_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7624_ (.A1(_3562_),
    .A2(_3575_),
    .B(_3615_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7625_ (.I(net2),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7626_ (.I(net32),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7627_ (.A1(_3616_),
    .A2(_3617_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7628_ (.I(_3324_),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7629_ (.A1(_3320_),
    .A2(_3565_),
    .A3(_3619_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7630_ (.A1(_3618_),
    .A2(_3620_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7631_ (.I(_3621_),
    .Z(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7632_ (.I(_3622_),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7633_ (.I0(\reg_file.reg_storage[8][0] ),
    .I1(_3319_),
    .S(_3623_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7634_ (.I(_3624_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7635_ (.I0(\reg_file.reg_storage[8][1] ),
    .I1(_3337_),
    .S(_3623_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7636_ (.I(_3625_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7637_ (.I(_3621_),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _7638_ (.I(_3626_),
    .Z(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7639_ (.I(_3627_),
    .Z(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7640_ (.I(_3621_),
    .Z(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7641_ (.I(_3629_),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7642_ (.A1(\reg_file.reg_storage[8][2] ),
    .A2(_3630_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7643_ (.A1(_3353_),
    .A2(_3628_),
    .B(_3631_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7644_ (.A1(\reg_file.reg_storage[8][3] ),
    .A2(_3630_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7645_ (.A1(_3363_),
    .A2(_3628_),
    .B(_3632_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7646_ (.I0(\reg_file.reg_storage[8][4] ),
    .I1(_3369_),
    .S(_3623_),
    .Z(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7647_ (.I(_3633_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7648_ (.I(_3622_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7649_ (.A1(\reg_file.reg_storage[8][5] ),
    .A2(_3634_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7650_ (.A1(_3376_),
    .A2(_3628_),
    .B(_3635_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7651_ (.A1(\reg_file.reg_storage[8][6] ),
    .A2(_3634_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7652_ (.A1(_3385_),
    .A2(_3628_),
    .B(_3636_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7653_ (.I(_3627_),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7654_ (.A1(\reg_file.reg_storage[8][7] ),
    .A2(_3634_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7655_ (.A1(_3395_),
    .A2(_3637_),
    .B(_3638_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7656_ (.A1(\reg_file.reg_storage[8][8] ),
    .A2(_3634_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7657_ (.A1(_3401_),
    .A2(_3637_),
    .B(_3639_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7658_ (.I(_3622_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7659_ (.A1(\reg_file.reg_storage[8][9] ),
    .A2(_3640_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7660_ (.A1(_3406_),
    .A2(_3637_),
    .B(_3641_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7661_ (.A1(\reg_file.reg_storage[8][10] ),
    .A2(_3640_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7662_ (.A1(_3413_),
    .A2(_3637_),
    .B(_3642_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7663_ (.I(_3627_),
    .Z(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7664_ (.A1(\reg_file.reg_storage[8][11] ),
    .A2(_3640_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7665_ (.A1(_3420_),
    .A2(_3643_),
    .B(_3644_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7666_ (.I(_3622_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7667_ (.I0(\reg_file.reg_storage[8][12] ),
    .I1(_3430_),
    .S(_3645_),
    .Z(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7668_ (.I(_3646_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7669_ (.A1(\reg_file.reg_storage[8][13] ),
    .A2(_3640_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7670_ (.A1(_3439_),
    .A2(_3643_),
    .B(_3647_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7671_ (.I(_3626_),
    .Z(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7672_ (.A1(\reg_file.reg_storage[8][14] ),
    .A2(_3648_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7673_ (.A1(_3447_),
    .A2(_3643_),
    .B(_3649_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7674_ (.A1(\reg_file.reg_storage[8][15] ),
    .A2(_3648_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7675_ (.A1(_3453_),
    .A2(_3643_),
    .B(_3650_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7676_ (.I0(\reg_file.reg_storage[8][16] ),
    .I1(_3460_),
    .S(_3645_),
    .Z(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7677_ (.I(_3651_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7678_ (.I(_3627_),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7679_ (.A1(\reg_file.reg_storage[8][17] ),
    .A2(_3648_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7680_ (.A1(_3467_),
    .A2(_3652_),
    .B(_3653_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7681_ (.A1(\reg_file.reg_storage[8][18] ),
    .A2(_3648_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7682_ (.A1(_3475_),
    .A2(_3652_),
    .B(_3654_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7683_ (.I(_3626_),
    .Z(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7684_ (.A1(\reg_file.reg_storage[8][19] ),
    .A2(_3655_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7685_ (.A1(_3482_),
    .A2(_3652_),
    .B(_3656_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7686_ (.I0(\reg_file.reg_storage[8][20] ),
    .I1(_3490_),
    .S(_3645_),
    .Z(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7687_ (.I(_3657_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7688_ (.I0(\reg_file.reg_storage[8][21] ),
    .I1(_3497_),
    .S(_3645_),
    .Z(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7689_ (.I(_3658_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7690_ (.I0(\reg_file.reg_storage[8][22] ),
    .I1(_3504_),
    .S(_3629_),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7691_ (.I(_3659_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7692_ (.A1(\reg_file.reg_storage[8][23] ),
    .A2(_3655_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7693_ (.A1(_3510_),
    .A2(_3652_),
    .B(_3660_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7694_ (.I(_3623_),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7695_ (.A1(\reg_file.reg_storage[8][24] ),
    .A2(_3655_),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7696_ (.A1(_3516_),
    .A2(_3661_),
    .B(_3662_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7697_ (.A1(\reg_file.reg_storage[8][25] ),
    .A2(_3655_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7698_ (.A1(_3525_),
    .A2(_3661_),
    .B(_3663_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7699_ (.I(_3626_),
    .Z(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7700_ (.A1(\reg_file.reg_storage[8][26] ),
    .A2(_3664_),
    .ZN(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7701_ (.A1(_3531_),
    .A2(_3661_),
    .B(_3665_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7702_ (.A1(\reg_file.reg_storage[8][27] ),
    .A2(_3664_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7703_ (.A1(_3538_),
    .A2(_3661_),
    .B(_3666_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7704_ (.A1(\reg_file.reg_storage[8][28] ),
    .A2(_3664_),
    .ZN(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7705_ (.A1(_3544_),
    .A2(_3630_),
    .B(_3667_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7706_ (.I0(\reg_file.reg_storage[8][29] ),
    .I1(_3551_),
    .S(_3629_),
    .Z(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7707_ (.I(_3668_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7708_ (.I0(\reg_file.reg_storage[8][30] ),
    .I1(_3557_),
    .S(_3629_),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7709_ (.I(_3669_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7710_ (.A1(\reg_file.reg_storage[8][31] ),
    .A2(_3664_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7711_ (.A1(_3562_),
    .A2(_3630_),
    .B(_3670_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7712_ (.A1(_3564_),
    .A2(_3321_),
    .A3(_3619_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7713_ (.A1(_3618_),
    .A2(_3671_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7714_ (.I(_3672_),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7715_ (.I(_3673_),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7716_ (.I0(\reg_file.reg_storage[11][0] ),
    .I1(_3319_),
    .S(_3674_),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7717_ (.I(_3675_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7718_ (.I0(\reg_file.reg_storage[11][1] ),
    .I1(_3337_),
    .S(_3674_),
    .Z(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7719_ (.I(_3676_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7720_ (.I(_3672_),
    .Z(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7721_ (.I(_3677_),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7722_ (.I(_3678_),
    .Z(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7723_ (.I(_3672_),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7724_ (.I(_3680_),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7725_ (.A1(\reg_file.reg_storage[11][2] ),
    .A2(_3681_),
    .ZN(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7726_ (.A1(_3353_),
    .A2(_3679_),
    .B(_3682_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7727_ (.A1(\reg_file.reg_storage[11][3] ),
    .A2(_3681_),
    .ZN(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7728_ (.A1(_3363_),
    .A2(_3679_),
    .B(_3683_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7729_ (.I0(\reg_file.reg_storage[11][4] ),
    .I1(_3369_),
    .S(_3674_),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7730_ (.I(_3684_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7731_ (.I(_3673_),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7732_ (.A1(\reg_file.reg_storage[11][5] ),
    .A2(_3685_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7733_ (.A1(_3376_),
    .A2(_3679_),
    .B(_3686_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7734_ (.A1(\reg_file.reg_storage[11][6] ),
    .A2(_3685_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7735_ (.A1(_3385_),
    .A2(_3679_),
    .B(_3687_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7736_ (.I(_3678_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7737_ (.A1(\reg_file.reg_storage[11][7] ),
    .A2(_3685_),
    .ZN(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7738_ (.A1(_3395_),
    .A2(_3688_),
    .B(_3689_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7739_ (.A1(\reg_file.reg_storage[11][8] ),
    .A2(_3685_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7740_ (.A1(_3401_),
    .A2(_3688_),
    .B(_3690_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7741_ (.I(_3673_),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7742_ (.A1(\reg_file.reg_storage[11][9] ),
    .A2(_3691_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7743_ (.A1(_3406_),
    .A2(_3688_),
    .B(_3692_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7744_ (.A1(\reg_file.reg_storage[11][10] ),
    .A2(_3691_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7745_ (.A1(_3413_),
    .A2(_3688_),
    .B(_3693_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7746_ (.I(_3678_),
    .Z(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7747_ (.A1(\reg_file.reg_storage[11][11] ),
    .A2(_3691_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7748_ (.A1(_3420_),
    .A2(_3694_),
    .B(_3695_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7749_ (.I(_3673_),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7750_ (.I0(\reg_file.reg_storage[11][12] ),
    .I1(_3430_),
    .S(_3696_),
    .Z(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7751_ (.I(_3697_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7752_ (.A1(\reg_file.reg_storage[11][13] ),
    .A2(_3691_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7753_ (.A1(_3439_),
    .A2(_3694_),
    .B(_3698_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7754_ (.I(_3677_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7755_ (.A1(\reg_file.reg_storage[11][14] ),
    .A2(_3699_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7756_ (.A1(_3447_),
    .A2(_3694_),
    .B(_3700_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7757_ (.A1(\reg_file.reg_storage[11][15] ),
    .A2(_3699_),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7758_ (.A1(_3453_),
    .A2(_3694_),
    .B(_3701_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7759_ (.I0(\reg_file.reg_storage[11][16] ),
    .I1(_3460_),
    .S(_3696_),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7760_ (.I(_3702_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7761_ (.I(_3678_),
    .Z(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7762_ (.A1(\reg_file.reg_storage[11][17] ),
    .A2(_3699_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7763_ (.A1(_3467_),
    .A2(_3703_),
    .B(_3704_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7764_ (.A1(\reg_file.reg_storage[11][18] ),
    .A2(_3699_),
    .ZN(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7765_ (.A1(_3475_),
    .A2(_3703_),
    .B(_3705_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7766_ (.I(_3677_),
    .Z(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7767_ (.A1(\reg_file.reg_storage[11][19] ),
    .A2(_3706_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7768_ (.A1(_3482_),
    .A2(_3703_),
    .B(_3707_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7769_ (.I0(\reg_file.reg_storage[11][20] ),
    .I1(_3490_),
    .S(_3696_),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7770_ (.I(_3708_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7771_ (.I0(\reg_file.reg_storage[11][21] ),
    .I1(_3497_),
    .S(_3696_),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7772_ (.I(_3709_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7773_ (.I0(\reg_file.reg_storage[11][22] ),
    .I1(_3504_),
    .S(_3680_),
    .Z(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7774_ (.I(_3710_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7775_ (.A1(\reg_file.reg_storage[11][23] ),
    .A2(_3706_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7776_ (.A1(_3510_),
    .A2(_3703_),
    .B(_3711_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7777_ (.I(_3674_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7778_ (.A1(\reg_file.reg_storage[11][24] ),
    .A2(_3706_),
    .ZN(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7779_ (.A1(_3516_),
    .A2(_3712_),
    .B(_3713_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7780_ (.A1(\reg_file.reg_storage[11][25] ),
    .A2(_3706_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7781_ (.A1(_3525_),
    .A2(_3712_),
    .B(_3714_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7782_ (.I(_3677_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7783_ (.A1(\reg_file.reg_storage[11][26] ),
    .A2(_3715_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7784_ (.A1(_3531_),
    .A2(_3712_),
    .B(_3716_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7785_ (.A1(\reg_file.reg_storage[11][27] ),
    .A2(_3715_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7786_ (.A1(_3538_),
    .A2(_3712_),
    .B(_3717_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7787_ (.A1(\reg_file.reg_storage[11][28] ),
    .A2(_3715_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7788_ (.A1(_3544_),
    .A2(_3681_),
    .B(_3718_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7789_ (.I0(\reg_file.reg_storage[11][29] ),
    .I1(_3551_),
    .S(_3680_),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7790_ (.I(_3719_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7791_ (.I0(\reg_file.reg_storage[11][30] ),
    .I1(_3557_),
    .S(_3680_),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7792_ (.I(_3720_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7793_ (.A1(\reg_file.reg_storage[11][31] ),
    .A2(_3715_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7794_ (.A1(_3562_),
    .A2(_3681_),
    .B(_3721_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7795_ (.I(_3317_),
    .Z(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7796_ (.A1(_3320_),
    .A2(_3321_),
    .A3(_3619_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7797_ (.A1(_3618_),
    .A2(_3723_),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7798_ (.I(_3724_),
    .Z(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _7799_ (.I(_3725_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7800_ (.I0(\reg_file.reg_storage[9][0] ),
    .I1(_3722_),
    .S(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7801_ (.I(_3727_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7802_ (.I(_3335_),
    .Z(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7803_ (.I0(\reg_file.reg_storage[9][1] ),
    .I1(_3728_),
    .S(_3726_),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7804_ (.I(_3729_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7805_ (.I(_3352_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7806_ (.I(_3730_),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7807_ (.I(_3724_),
    .Z(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7808_ (.I(_3732_),
    .Z(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7809_ (.I(_3733_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7810_ (.I(_3724_),
    .Z(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7811_ (.I(_3735_),
    .Z(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7812_ (.A1(\reg_file.reg_storage[9][2] ),
    .A2(_3736_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7813_ (.A1(_3731_),
    .A2(_3734_),
    .B(_3737_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7814_ (.I(_3362_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7815_ (.I(_3738_),
    .Z(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7816_ (.A1(\reg_file.reg_storage[9][3] ),
    .A2(_3736_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7817_ (.A1(_3739_),
    .A2(_3734_),
    .B(_3740_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7818_ (.I(_3367_),
    .Z(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7819_ (.I0(\reg_file.reg_storage[9][4] ),
    .I1(_3741_),
    .S(_3726_),
    .Z(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7820_ (.I(_3742_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7821_ (.I(_3375_),
    .Z(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7822_ (.I(_3743_),
    .Z(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7823_ (.I(_3725_),
    .Z(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7824_ (.A1(\reg_file.reg_storage[9][5] ),
    .A2(_3745_),
    .ZN(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7825_ (.A1(_3744_),
    .A2(_3734_),
    .B(_3746_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7826_ (.I(_3384_),
    .Z(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7827_ (.I(_3747_),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7828_ (.A1(\reg_file.reg_storage[9][6] ),
    .A2(_3745_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7829_ (.A1(_3748_),
    .A2(_3734_),
    .B(_3749_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7830_ (.I(_3394_),
    .Z(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7831_ (.I(_3750_),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7832_ (.I(_3733_),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7833_ (.A1(\reg_file.reg_storage[9][7] ),
    .A2(_3745_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7834_ (.A1(_3751_),
    .A2(_3752_),
    .B(_3753_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7835_ (.I(_3400_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7836_ (.I(_3754_),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7837_ (.A1(\reg_file.reg_storage[9][8] ),
    .A2(_3745_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7838_ (.A1(_3755_),
    .A2(_3752_),
    .B(_3756_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7839_ (.I(_3405_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7840_ (.I(_3757_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7841_ (.I(_3725_),
    .Z(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7842_ (.A1(\reg_file.reg_storage[9][9] ),
    .A2(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7843_ (.A1(_3758_),
    .A2(_3752_),
    .B(_3760_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7844_ (.I(_3412_),
    .Z(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7845_ (.I(_3761_),
    .Z(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7846_ (.A1(\reg_file.reg_storage[9][10] ),
    .A2(_3759_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7847_ (.A1(_3762_),
    .A2(_3752_),
    .B(_3763_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7848_ (.I(_3419_),
    .Z(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7849_ (.I(_3764_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7850_ (.I(_3733_),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7851_ (.A1(\reg_file.reg_storage[9][11] ),
    .A2(_3759_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7852_ (.A1(_3765_),
    .A2(_3766_),
    .B(_3767_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7853_ (.I(_3428_),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7854_ (.I(_3725_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7855_ (.I0(\reg_file.reg_storage[9][12] ),
    .I1(_3768_),
    .S(_3769_),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7856_ (.I(_3770_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7857_ (.I(_3438_),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7858_ (.I(_3771_),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7859_ (.A1(\reg_file.reg_storage[9][13] ),
    .A2(_3759_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7860_ (.A1(_3772_),
    .A2(_3766_),
    .B(_3773_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7861_ (.I(_3446_),
    .Z(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7862_ (.I(_3774_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7863_ (.I(_3732_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7864_ (.A1(\reg_file.reg_storage[9][14] ),
    .A2(_3776_),
    .ZN(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7865_ (.A1(_3775_),
    .A2(_3766_),
    .B(_3777_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7866_ (.I(_3452_),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7867_ (.I(_3778_),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7868_ (.A1(\reg_file.reg_storage[9][15] ),
    .A2(_3776_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7869_ (.A1(_3779_),
    .A2(_3766_),
    .B(_3780_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7870_ (.I(_3458_),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7871_ (.I0(\reg_file.reg_storage[9][16] ),
    .I1(_3781_),
    .S(_3769_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7872_ (.I(_3782_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7873_ (.I(_3466_),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7874_ (.I(_3783_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7875_ (.I(_3733_),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7876_ (.A1(\reg_file.reg_storage[9][17] ),
    .A2(_3776_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7877_ (.A1(_3784_),
    .A2(_3785_),
    .B(_3786_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7878_ (.I(_3474_),
    .Z(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7879_ (.I(_3787_),
    .Z(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7880_ (.A1(\reg_file.reg_storage[9][18] ),
    .A2(_3776_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7881_ (.A1(_3788_),
    .A2(_3785_),
    .B(_3789_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7882_ (.I(_3481_),
    .Z(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7883_ (.I(_3790_),
    .Z(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7884_ (.I(_3732_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7885_ (.A1(\reg_file.reg_storage[9][19] ),
    .A2(_3792_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7886_ (.A1(_3791_),
    .A2(_3785_),
    .B(_3793_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7887_ (.I(_3488_),
    .Z(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7888_ (.I0(\reg_file.reg_storage[9][20] ),
    .I1(_3794_),
    .S(_3769_),
    .Z(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7889_ (.I(_3795_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7890_ (.I(_3495_),
    .Z(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7891_ (.I0(\reg_file.reg_storage[9][21] ),
    .I1(_3796_),
    .S(_3769_),
    .Z(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7892_ (.I(_3797_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7893_ (.I(_3502_),
    .Z(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7894_ (.I0(\reg_file.reg_storage[9][22] ),
    .I1(_3798_),
    .S(_3735_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7895_ (.I(_3799_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7896_ (.I(_3509_),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7897_ (.I(_3800_),
    .Z(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7898_ (.A1(\reg_file.reg_storage[9][23] ),
    .A2(_3792_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7899_ (.A1(_3801_),
    .A2(_3785_),
    .B(_3802_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7900_ (.I(_3515_),
    .Z(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7901_ (.I(_3803_),
    .Z(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7902_ (.I(_3726_),
    .Z(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7903_ (.A1(\reg_file.reg_storage[9][24] ),
    .A2(_3792_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7904_ (.A1(_3804_),
    .A2(_3805_),
    .B(_3806_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7905_ (.I(_3524_),
    .Z(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7906_ (.I(_3807_),
    .Z(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7907_ (.A1(\reg_file.reg_storage[9][25] ),
    .A2(_3792_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7908_ (.A1(_3808_),
    .A2(_3805_),
    .B(_3809_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7909_ (.I(_3530_),
    .Z(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7910_ (.I(_3810_),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7911_ (.I(_3732_),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7912_ (.A1(\reg_file.reg_storage[9][26] ),
    .A2(_3812_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7913_ (.A1(_3811_),
    .A2(_3805_),
    .B(_3813_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7914_ (.I(_3537_),
    .Z(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7915_ (.I(_3814_),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7916_ (.A1(\reg_file.reg_storage[9][27] ),
    .A2(_3812_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7917_ (.A1(_3815_),
    .A2(_3805_),
    .B(_3816_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7918_ (.I(_3543_),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7919_ (.I(_3817_),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7920_ (.A1(\reg_file.reg_storage[9][28] ),
    .A2(_3812_),
    .ZN(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7921_ (.A1(_3818_),
    .A2(_3736_),
    .B(_3819_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7922_ (.I(_3549_),
    .Z(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7923_ (.I0(\reg_file.reg_storage[9][29] ),
    .I1(_3820_),
    .S(_3735_),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7924_ (.I(_3821_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7925_ (.I(_3555_),
    .Z(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7926_ (.I0(\reg_file.reg_storage[9][30] ),
    .I1(_3822_),
    .S(_3735_),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7927_ (.I(_3823_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7928_ (.I(_3561_),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7929_ (.I(_3824_),
    .Z(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7930_ (.A1(\reg_file.reg_storage[9][31] ),
    .A2(_3812_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7931_ (.A1(_3825_),
    .A2(_3736_),
    .B(_3826_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7932_ (.A1(net2),
    .A2(_3617_),
    .Z(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7933_ (.A1(_3564_),
    .A2(_3565_),
    .A3(_3619_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7934_ (.A1(_3827_),
    .A2(_3828_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7935_ (.I(_3829_),
    .Z(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _7936_ (.I(_3830_),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7937_ (.I0(\reg_file.reg_storage[6][0] ),
    .I1(_3722_),
    .S(_3831_),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7938_ (.I(_3832_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7939_ (.I0(\reg_file.reg_storage[6][1] ),
    .I1(_3728_),
    .S(_3831_),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7940_ (.I(_3833_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7941_ (.I(_3829_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7942_ (.I(_3834_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7943_ (.I(_3835_),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7944_ (.I(_3829_),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7945_ (.I(_3837_),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7946_ (.A1(\reg_file.reg_storage[6][2] ),
    .A2(_3838_),
    .ZN(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7947_ (.A1(_3731_),
    .A2(_3836_),
    .B(_3839_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7948_ (.A1(\reg_file.reg_storage[6][3] ),
    .A2(_3838_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7949_ (.A1(_3739_),
    .A2(_3836_),
    .B(_3840_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7950_ (.I0(\reg_file.reg_storage[6][4] ),
    .I1(_3741_),
    .S(_3831_),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7951_ (.I(_3841_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7952_ (.I(_3830_),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7953_ (.A1(\reg_file.reg_storage[6][5] ),
    .A2(_3842_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7954_ (.A1(_3744_),
    .A2(_3836_),
    .B(_3843_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7955_ (.A1(\reg_file.reg_storage[6][6] ),
    .A2(_3842_),
    .ZN(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7956_ (.A1(_3748_),
    .A2(_3836_),
    .B(_3844_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7957_ (.I(_3835_),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7958_ (.A1(\reg_file.reg_storage[6][7] ),
    .A2(_3842_),
    .ZN(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7959_ (.A1(_3751_),
    .A2(_3845_),
    .B(_3846_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7960_ (.A1(\reg_file.reg_storage[6][8] ),
    .A2(_3842_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7961_ (.A1(_3755_),
    .A2(_3845_),
    .B(_3847_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7962_ (.I(_3830_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7963_ (.A1(\reg_file.reg_storage[6][9] ),
    .A2(_3848_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7964_ (.A1(_3758_),
    .A2(_3845_),
    .B(_3849_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7965_ (.A1(\reg_file.reg_storage[6][10] ),
    .A2(_3848_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7966_ (.A1(_3762_),
    .A2(_3845_),
    .B(_3850_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7967_ (.I(_3835_),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7968_ (.A1(\reg_file.reg_storage[6][11] ),
    .A2(_3848_),
    .ZN(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7969_ (.A1(_3765_),
    .A2(_3851_),
    .B(_3852_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7970_ (.I(_3830_),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7971_ (.I0(\reg_file.reg_storage[6][12] ),
    .I1(_3768_),
    .S(_3853_),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7972_ (.I(_3854_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7973_ (.A1(\reg_file.reg_storage[6][13] ),
    .A2(_3848_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7974_ (.A1(_3772_),
    .A2(_3851_),
    .B(_3855_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7975_ (.I(_3834_),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7976_ (.A1(\reg_file.reg_storage[6][14] ),
    .A2(_3856_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7977_ (.A1(_3775_),
    .A2(_3851_),
    .B(_3857_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7978_ (.A1(\reg_file.reg_storage[6][15] ),
    .A2(_3856_),
    .ZN(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7979_ (.A1(_3779_),
    .A2(_3851_),
    .B(_3858_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7980_ (.I0(\reg_file.reg_storage[6][16] ),
    .I1(_3781_),
    .S(_3853_),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7981_ (.I(_3859_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7982_ (.I(_3835_),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7983_ (.A1(\reg_file.reg_storage[6][17] ),
    .A2(_3856_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7984_ (.A1(_3784_),
    .A2(_3860_),
    .B(_3861_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7985_ (.A1(\reg_file.reg_storage[6][18] ),
    .A2(_3856_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7986_ (.A1(_3788_),
    .A2(_3860_),
    .B(_3862_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7987_ (.I(_3834_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7988_ (.A1(\reg_file.reg_storage[6][19] ),
    .A2(_3863_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7989_ (.A1(_3791_),
    .A2(_3860_),
    .B(_3864_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7990_ (.I0(\reg_file.reg_storage[6][20] ),
    .I1(_3794_),
    .S(_3853_),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7991_ (.I(_3865_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7992_ (.I0(\reg_file.reg_storage[6][21] ),
    .I1(_3796_),
    .S(_3853_),
    .Z(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7993_ (.I(_3866_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7994_ (.I0(\reg_file.reg_storage[6][22] ),
    .I1(_3798_),
    .S(_3837_),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7995_ (.I(_3867_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7996_ (.A1(\reg_file.reg_storage[6][23] ),
    .A2(_3863_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7997_ (.A1(_3801_),
    .A2(_3860_),
    .B(_3868_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7998_ (.I(_3831_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7999_ (.A1(\reg_file.reg_storage[6][24] ),
    .A2(_3863_),
    .ZN(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8000_ (.A1(_3804_),
    .A2(_3869_),
    .B(_3870_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8001_ (.A1(\reg_file.reg_storage[6][25] ),
    .A2(_3863_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8002_ (.A1(_3808_),
    .A2(_3869_),
    .B(_3871_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8003_ (.I(_3834_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8004_ (.A1(\reg_file.reg_storage[6][26] ),
    .A2(_3872_),
    .ZN(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8005_ (.A1(_3811_),
    .A2(_3869_),
    .B(_3873_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8006_ (.A1(\reg_file.reg_storage[6][27] ),
    .A2(_3872_),
    .ZN(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8007_ (.A1(_3815_),
    .A2(_3869_),
    .B(_3874_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8008_ (.A1(\reg_file.reg_storage[6][28] ),
    .A2(_3872_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8009_ (.A1(_3818_),
    .A2(_3838_),
    .B(_3875_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8010_ (.I0(\reg_file.reg_storage[6][29] ),
    .I1(_3820_),
    .S(_3837_),
    .Z(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8011_ (.I(_3876_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8012_ (.I0(\reg_file.reg_storage[6][30] ),
    .I1(_3822_),
    .S(_3837_),
    .Z(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8013_ (.I(_3877_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8014_ (.A1(\reg_file.reg_storage[6][31] ),
    .A2(_3872_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8015_ (.A1(_3825_),
    .A2(_3838_),
    .B(_3878_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8016_ (.A1(_3616_),
    .A2(_3322_),
    .A3(_3723_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8017_ (.I(_3879_),
    .Z(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8018_ (.I(_3880_),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8019_ (.I0(\reg_file.reg_storage[1][0] ),
    .I1(_3722_),
    .S(_3881_),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8020_ (.I(_3882_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8021_ (.I0(\reg_file.reg_storage[1][1] ),
    .I1(_3728_),
    .S(_3881_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8022_ (.I(_3883_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8023_ (.I(_3879_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8024_ (.I(_3884_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8025_ (.I(_3885_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8026_ (.I(_3879_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8027_ (.I(_3887_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8028_ (.A1(\reg_file.reg_storage[1][2] ),
    .A2(_3888_),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8029_ (.A1(_3731_),
    .A2(_3886_),
    .B(_3889_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8030_ (.A1(\reg_file.reg_storage[1][3] ),
    .A2(_3888_),
    .ZN(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8031_ (.A1(_3739_),
    .A2(_3886_),
    .B(_3890_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8032_ (.I0(\reg_file.reg_storage[1][4] ),
    .I1(_3741_),
    .S(_3881_),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8033_ (.I(_3891_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8034_ (.I(_3880_),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8035_ (.A1(\reg_file.reg_storage[1][5] ),
    .A2(_3892_),
    .ZN(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8036_ (.A1(_3744_),
    .A2(_3886_),
    .B(_3893_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8037_ (.A1(\reg_file.reg_storage[1][6] ),
    .A2(_3892_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8038_ (.A1(_3748_),
    .A2(_3886_),
    .B(_3894_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8039_ (.I(_3885_),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8040_ (.A1(\reg_file.reg_storage[1][7] ),
    .A2(_3892_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8041_ (.A1(_3751_),
    .A2(_3895_),
    .B(_3896_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8042_ (.A1(\reg_file.reg_storage[1][8] ),
    .A2(_3892_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8043_ (.A1(_3755_),
    .A2(_3895_),
    .B(_3897_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8044_ (.I(_3880_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8045_ (.A1(\reg_file.reg_storage[1][9] ),
    .A2(_3898_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8046_ (.A1(_3758_),
    .A2(_3895_),
    .B(_3899_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8047_ (.A1(\reg_file.reg_storage[1][10] ),
    .A2(_3898_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8048_ (.A1(_3762_),
    .A2(_3895_),
    .B(_3900_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8049_ (.I(_3885_),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8050_ (.A1(\reg_file.reg_storage[1][11] ),
    .A2(_3898_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8051_ (.A1(_3765_),
    .A2(_3901_),
    .B(_3902_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8052_ (.I(_3880_),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8053_ (.I0(\reg_file.reg_storage[1][12] ),
    .I1(_3768_),
    .S(_3903_),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8054_ (.I(_3904_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8055_ (.A1(\reg_file.reg_storage[1][13] ),
    .A2(_3898_),
    .ZN(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8056_ (.A1(_3772_),
    .A2(_3901_),
    .B(_3905_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8057_ (.I(_3884_),
    .Z(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8058_ (.A1(\reg_file.reg_storage[1][14] ),
    .A2(_3906_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8059_ (.A1(_3775_),
    .A2(_3901_),
    .B(_3907_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8060_ (.A1(\reg_file.reg_storage[1][15] ),
    .A2(_3906_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8061_ (.A1(_3779_),
    .A2(_3901_),
    .B(_3908_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8062_ (.I0(\reg_file.reg_storage[1][16] ),
    .I1(_3781_),
    .S(_3903_),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8063_ (.I(_3909_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8064_ (.I(_3885_),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8065_ (.A1(\reg_file.reg_storage[1][17] ),
    .A2(_3906_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8066_ (.A1(_3784_),
    .A2(_3910_),
    .B(_3911_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8067_ (.A1(\reg_file.reg_storage[1][18] ),
    .A2(_3906_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8068_ (.A1(_3788_),
    .A2(_3910_),
    .B(_3912_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8069_ (.I(_3884_),
    .Z(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8070_ (.A1(\reg_file.reg_storage[1][19] ),
    .A2(_3913_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8071_ (.A1(_3791_),
    .A2(_3910_),
    .B(_3914_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8072_ (.I0(\reg_file.reg_storage[1][20] ),
    .I1(_3794_),
    .S(_3903_),
    .Z(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8073_ (.I(_3915_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8074_ (.I0(\reg_file.reg_storage[1][21] ),
    .I1(_3796_),
    .S(_3903_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8075_ (.I(_3916_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8076_ (.I0(\reg_file.reg_storage[1][22] ),
    .I1(_3798_),
    .S(_3887_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8077_ (.I(_3917_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8078_ (.A1(\reg_file.reg_storage[1][23] ),
    .A2(_3913_),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8079_ (.A1(_3801_),
    .A2(_3910_),
    .B(_3918_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8080_ (.I(_3881_),
    .Z(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8081_ (.A1(\reg_file.reg_storage[1][24] ),
    .A2(_3913_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8082_ (.A1(_3804_),
    .A2(_3919_),
    .B(_3920_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8083_ (.A1(\reg_file.reg_storage[1][25] ),
    .A2(_3913_),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8084_ (.A1(_3808_),
    .A2(_3919_),
    .B(_3921_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8085_ (.I(_3884_),
    .Z(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8086_ (.A1(\reg_file.reg_storage[1][26] ),
    .A2(_3922_),
    .ZN(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8087_ (.A1(_3811_),
    .A2(_3919_),
    .B(_3923_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8088_ (.A1(\reg_file.reg_storage[1][27] ),
    .A2(_3922_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8089_ (.A1(_3815_),
    .A2(_3919_),
    .B(_3924_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8090_ (.A1(\reg_file.reg_storage[1][28] ),
    .A2(_3922_),
    .ZN(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8091_ (.A1(_3818_),
    .A2(_3888_),
    .B(_3925_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8092_ (.I0(\reg_file.reg_storage[1][29] ),
    .I1(_3820_),
    .S(_3887_),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8093_ (.I(_3926_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8094_ (.I0(\reg_file.reg_storage[1][30] ),
    .I1(_3822_),
    .S(_3887_),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8095_ (.I(_3927_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8096_ (.A1(\reg_file.reg_storage[1][31] ),
    .A2(_3922_),
    .ZN(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8097_ (.A1(_3825_),
    .A2(_3888_),
    .B(_3928_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8098_ (.A1(_3616_),
    .A2(_3322_),
    .A3(_3671_),
    .ZN(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8099_ (.I(_3929_),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8100_ (.I(_3930_),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8101_ (.I0(\reg_file.reg_storage[3][0] ),
    .I1(_3722_),
    .S(_3931_),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8102_ (.I(_3932_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8103_ (.I0(\reg_file.reg_storage[3][1] ),
    .I1(_3728_),
    .S(_3931_),
    .Z(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8104_ (.I(_3933_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8105_ (.I(_3929_),
    .Z(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8106_ (.I(_3934_),
    .Z(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8107_ (.I(_3935_),
    .Z(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8108_ (.I(_3929_),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8109_ (.I(_3937_),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8110_ (.A1(\reg_file.reg_storage[3][2] ),
    .A2(_3938_),
    .ZN(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8111_ (.A1(_3731_),
    .A2(_3936_),
    .B(_3939_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8112_ (.A1(\reg_file.reg_storage[3][3] ),
    .A2(_3938_),
    .ZN(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8113_ (.A1(_3739_),
    .A2(_3936_),
    .B(_3940_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8114_ (.I0(\reg_file.reg_storage[3][4] ),
    .I1(_3741_),
    .S(_3931_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8115_ (.I(_3941_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8116_ (.I(_3930_),
    .Z(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8117_ (.A1(\reg_file.reg_storage[3][5] ),
    .A2(_3942_),
    .ZN(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8118_ (.A1(_3744_),
    .A2(_3936_),
    .B(_3943_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8119_ (.A1(\reg_file.reg_storage[3][6] ),
    .A2(_3942_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8120_ (.A1(_3748_),
    .A2(_3936_),
    .B(_3944_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8121_ (.I(_3935_),
    .Z(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8122_ (.A1(\reg_file.reg_storage[3][7] ),
    .A2(_3942_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8123_ (.A1(_3751_),
    .A2(_3945_),
    .B(_3946_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8124_ (.A1(\reg_file.reg_storage[3][8] ),
    .A2(_3942_),
    .ZN(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8125_ (.A1(_3755_),
    .A2(_3945_),
    .B(_3947_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8126_ (.I(_3930_),
    .Z(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8127_ (.A1(\reg_file.reg_storage[3][9] ),
    .A2(_3948_),
    .ZN(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8128_ (.A1(_3758_),
    .A2(_3945_),
    .B(_3949_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8129_ (.A1(\reg_file.reg_storage[3][10] ),
    .A2(_3948_),
    .ZN(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8130_ (.A1(_3762_),
    .A2(_3945_),
    .B(_3950_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8131_ (.I(_3935_),
    .Z(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8132_ (.A1(\reg_file.reg_storage[3][11] ),
    .A2(_3948_),
    .ZN(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8133_ (.A1(_3765_),
    .A2(_3951_),
    .B(_3952_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8134_ (.I(_3930_),
    .Z(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8135_ (.I0(\reg_file.reg_storage[3][12] ),
    .I1(_3768_),
    .S(_3953_),
    .Z(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8136_ (.I(_3954_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8137_ (.A1(\reg_file.reg_storage[3][13] ),
    .A2(_3948_),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8138_ (.A1(_3772_),
    .A2(_3951_),
    .B(_3955_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8139_ (.I(_3934_),
    .Z(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8140_ (.A1(\reg_file.reg_storage[3][14] ),
    .A2(_3956_),
    .ZN(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8141_ (.A1(_3775_),
    .A2(_3951_),
    .B(_3957_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8142_ (.A1(\reg_file.reg_storage[3][15] ),
    .A2(_3956_),
    .ZN(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8143_ (.A1(_3779_),
    .A2(_3951_),
    .B(_3958_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8144_ (.I0(\reg_file.reg_storage[3][16] ),
    .I1(_3781_),
    .S(_3953_),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8145_ (.I(_3959_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8146_ (.I(_3935_),
    .Z(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8147_ (.A1(\reg_file.reg_storage[3][17] ),
    .A2(_3956_),
    .ZN(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8148_ (.A1(_3784_),
    .A2(_3960_),
    .B(_3961_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8149_ (.A1(\reg_file.reg_storage[3][18] ),
    .A2(_3956_),
    .ZN(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8150_ (.A1(_3788_),
    .A2(_3960_),
    .B(_3962_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8151_ (.I(_3934_),
    .Z(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8152_ (.A1(\reg_file.reg_storage[3][19] ),
    .A2(_3963_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8153_ (.A1(_3791_),
    .A2(_3960_),
    .B(_3964_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8154_ (.I0(\reg_file.reg_storage[3][20] ),
    .I1(_3794_),
    .S(_3953_),
    .Z(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8155_ (.I(_3965_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8156_ (.I0(\reg_file.reg_storage[3][21] ),
    .I1(_3796_),
    .S(_3953_),
    .Z(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8157_ (.I(_3966_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8158_ (.I0(\reg_file.reg_storage[3][22] ),
    .I1(_3798_),
    .S(_3937_),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8159_ (.I(_3967_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8160_ (.A1(\reg_file.reg_storage[3][23] ),
    .A2(_3963_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8161_ (.A1(_3801_),
    .A2(_3960_),
    .B(_3968_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8162_ (.I(_3931_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8163_ (.A1(\reg_file.reg_storage[3][24] ),
    .A2(_3963_),
    .ZN(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8164_ (.A1(_3804_),
    .A2(_3969_),
    .B(_3970_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8165_ (.A1(\reg_file.reg_storage[3][25] ),
    .A2(_3963_),
    .ZN(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8166_ (.A1(_3808_),
    .A2(_3969_),
    .B(_3971_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8167_ (.I(_3934_),
    .Z(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8168_ (.A1(\reg_file.reg_storage[3][26] ),
    .A2(_3972_),
    .ZN(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8169_ (.A1(_3811_),
    .A2(_3969_),
    .B(_3973_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8170_ (.A1(\reg_file.reg_storage[3][27] ),
    .A2(_3972_),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8171_ (.A1(_3815_),
    .A2(_3969_),
    .B(_3974_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8172_ (.A1(\reg_file.reg_storage[3][28] ),
    .A2(_3972_),
    .ZN(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8173_ (.A1(_3818_),
    .A2(_3938_),
    .B(_3975_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8174_ (.I0(\reg_file.reg_storage[3][29] ),
    .I1(_3820_),
    .S(_3937_),
    .Z(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8175_ (.I(_3976_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8176_ (.I0(\reg_file.reg_storage[3][30] ),
    .I1(_3822_),
    .S(_3937_),
    .Z(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8177_ (.I(_3977_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8178_ (.A1(\reg_file.reg_storage[3][31] ),
    .A2(_3972_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8179_ (.A1(_3825_),
    .A2(_3938_),
    .B(_3978_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8180_ (.I(_3317_),
    .Z(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _8181_ (.A1(_3320_),
    .A2(_3565_),
    .A3(_3325_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8182_ (.I(_3980_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _8183_ (.I(_3981_),
    .Z(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8184_ (.I0(\reg_file.reg_storage[15][0] ),
    .I1(_3979_),
    .S(_3982_),
    .Z(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8185_ (.I(_3983_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8186_ (.I(_3335_),
    .Z(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8187_ (.I0(\reg_file.reg_storage[15][1] ),
    .I1(_3984_),
    .S(_3982_),
    .Z(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8188_ (.I(_3985_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8189_ (.I(_3352_),
    .Z(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8190_ (.I(_3980_),
    .Z(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8191_ (.I(_3987_),
    .Z(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8192_ (.I(_3988_),
    .Z(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8193_ (.I(_3980_),
    .Z(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8194_ (.I(_3990_),
    .Z(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8195_ (.A1(\reg_file.reg_storage[15][2] ),
    .A2(_3991_),
    .ZN(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8196_ (.A1(_3986_),
    .A2(_3989_),
    .B(_3992_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8197_ (.I(_3362_),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8198_ (.A1(\reg_file.reg_storage[15][3] ),
    .A2(_3991_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8199_ (.A1(_3993_),
    .A2(_3989_),
    .B(_3994_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8200_ (.I(_3367_),
    .Z(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8201_ (.I0(\reg_file.reg_storage[15][4] ),
    .I1(_3995_),
    .S(_3982_),
    .Z(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8202_ (.I(_3996_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8203_ (.I(_3375_),
    .Z(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8204_ (.I(_3981_),
    .Z(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8205_ (.A1(\reg_file.reg_storage[15][5] ),
    .A2(_3998_),
    .ZN(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8206_ (.A1(_3997_),
    .A2(_3989_),
    .B(_3999_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8207_ (.I(_3384_),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8208_ (.A1(\reg_file.reg_storage[15][6] ),
    .A2(_3998_),
    .ZN(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8209_ (.A1(_4000_),
    .A2(_3989_),
    .B(_4001_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8210_ (.I(_3394_),
    .Z(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8211_ (.I(_3988_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8212_ (.A1(\reg_file.reg_storage[15][7] ),
    .A2(_3998_),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8213_ (.A1(_4002_),
    .A2(_4003_),
    .B(_4004_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8214_ (.I(_3400_),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8215_ (.A1(\reg_file.reg_storage[15][8] ),
    .A2(_3998_),
    .ZN(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8216_ (.A1(_4005_),
    .A2(_4003_),
    .B(_4006_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8217_ (.I(_3405_),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8218_ (.I(_3981_),
    .Z(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8219_ (.A1(\reg_file.reg_storage[15][9] ),
    .A2(_4008_),
    .ZN(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8220_ (.A1(_4007_),
    .A2(_4003_),
    .B(_4009_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8221_ (.I(_3412_),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8222_ (.A1(\reg_file.reg_storage[15][10] ),
    .A2(_4008_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8223_ (.A1(_4010_),
    .A2(_4003_),
    .B(_4011_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8224_ (.I(_3419_),
    .Z(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8225_ (.I(_3988_),
    .Z(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8226_ (.A1(\reg_file.reg_storage[15][11] ),
    .A2(_4008_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8227_ (.A1(_4012_),
    .A2(_4013_),
    .B(_4014_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8228_ (.I(_3428_),
    .Z(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8229_ (.I(_3981_),
    .Z(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8230_ (.I0(\reg_file.reg_storage[15][12] ),
    .I1(_4015_),
    .S(_4016_),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8231_ (.I(_4017_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8232_ (.I(_3438_),
    .Z(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8233_ (.A1(\reg_file.reg_storage[15][13] ),
    .A2(_4008_),
    .ZN(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8234_ (.A1(_4018_),
    .A2(_4013_),
    .B(_4019_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8235_ (.I(_3446_),
    .Z(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8236_ (.I(_3987_),
    .Z(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8237_ (.A1(\reg_file.reg_storage[15][14] ),
    .A2(_4021_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8238_ (.A1(_4020_),
    .A2(_4013_),
    .B(_4022_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8239_ (.I(_3452_),
    .Z(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8240_ (.A1(\reg_file.reg_storage[15][15] ),
    .A2(_4021_),
    .ZN(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8241_ (.A1(_4023_),
    .A2(_4013_),
    .B(_4024_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8242_ (.I(_3458_),
    .Z(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8243_ (.I0(\reg_file.reg_storage[15][16] ),
    .I1(_4025_),
    .S(_4016_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8244_ (.I(_4026_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8245_ (.I(_3466_),
    .Z(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8246_ (.I(_3988_),
    .Z(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8247_ (.A1(\reg_file.reg_storage[15][17] ),
    .A2(_4021_),
    .ZN(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8248_ (.A1(_4027_),
    .A2(_4028_),
    .B(_4029_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8249_ (.I(_3474_),
    .Z(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8250_ (.A1(\reg_file.reg_storage[15][18] ),
    .A2(_4021_),
    .ZN(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8251_ (.A1(_4030_),
    .A2(_4028_),
    .B(_4031_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8252_ (.I(_3481_),
    .Z(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8253_ (.I(_3987_),
    .Z(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8254_ (.A1(\reg_file.reg_storage[15][19] ),
    .A2(_4033_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8255_ (.A1(_4032_),
    .A2(_4028_),
    .B(_4034_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8256_ (.I(_3488_),
    .Z(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8257_ (.I0(\reg_file.reg_storage[15][20] ),
    .I1(_4035_),
    .S(_4016_),
    .Z(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8258_ (.I(_4036_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8259_ (.I(_3495_),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8260_ (.I0(\reg_file.reg_storage[15][21] ),
    .I1(_4037_),
    .S(_4016_),
    .Z(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8261_ (.I(_4038_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8262_ (.I(_3502_),
    .Z(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8263_ (.I0(\reg_file.reg_storage[15][22] ),
    .I1(_4039_),
    .S(_3990_),
    .Z(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8264_ (.I(_4040_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8265_ (.I(_3509_),
    .Z(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8266_ (.A1(\reg_file.reg_storage[15][23] ),
    .A2(_4033_),
    .ZN(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8267_ (.A1(_4041_),
    .A2(_4028_),
    .B(_4042_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8268_ (.I(_3515_),
    .Z(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8269_ (.I(_3982_),
    .Z(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8270_ (.A1(\reg_file.reg_storage[15][24] ),
    .A2(_4033_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8271_ (.A1(_4043_),
    .A2(_4044_),
    .B(_4045_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8272_ (.I(_3524_),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8273_ (.A1(\reg_file.reg_storage[15][25] ),
    .A2(_4033_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8274_ (.A1(_4046_),
    .A2(_4044_),
    .B(_4047_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8275_ (.I(_3530_),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8276_ (.I(_3987_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8277_ (.A1(\reg_file.reg_storage[15][26] ),
    .A2(_4049_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8278_ (.A1(_4048_),
    .A2(_4044_),
    .B(_4050_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8279_ (.I(_3537_),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8280_ (.A1(\reg_file.reg_storage[15][27] ),
    .A2(_4049_),
    .ZN(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8281_ (.A1(_4051_),
    .A2(_4044_),
    .B(_4052_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8282_ (.I(_3543_),
    .Z(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8283_ (.A1(\reg_file.reg_storage[15][28] ),
    .A2(_4049_),
    .ZN(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8284_ (.A1(_4053_),
    .A2(_3991_),
    .B(_4054_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8285_ (.I(_3549_),
    .Z(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8286_ (.I0(\reg_file.reg_storage[15][29] ),
    .I1(_4055_),
    .S(_3990_),
    .Z(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8287_ (.I(_4056_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8288_ (.I(_3555_),
    .Z(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8289_ (.I0(\reg_file.reg_storage[15][30] ),
    .I1(_4057_),
    .S(_3990_),
    .Z(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8290_ (.I(_4058_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8291_ (.I(_3561_),
    .Z(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8292_ (.A1(\reg_file.reg_storage[15][31] ),
    .A2(_4049_),
    .ZN(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8293_ (.A1(_4059_),
    .A2(_3991_),
    .B(_4060_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8294_ (.A1(_3620_),
    .A2(_3827_),
    .ZN(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8295_ (.I(_4061_),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _8296_ (.I(_4062_),
    .Z(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8297_ (.I0(\reg_file.reg_storage[4][0] ),
    .I1(_3979_),
    .S(_4063_),
    .Z(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8298_ (.I(_4064_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8299_ (.I0(\reg_file.reg_storage[4][1] ),
    .I1(_3984_),
    .S(_4063_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8300_ (.I(_4065_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8301_ (.I(_4061_),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8302_ (.I(_4066_),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8303_ (.I(_4067_),
    .Z(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8304_ (.I(_4061_),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8305_ (.I(_4069_),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8306_ (.A1(\reg_file.reg_storage[4][2] ),
    .A2(_4070_),
    .ZN(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8307_ (.A1(_3986_),
    .A2(_4068_),
    .B(_4071_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8308_ (.A1(\reg_file.reg_storage[4][3] ),
    .A2(_4070_),
    .ZN(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8309_ (.A1(_3993_),
    .A2(_4068_),
    .B(_4072_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8310_ (.I0(\reg_file.reg_storage[4][4] ),
    .I1(_3995_),
    .S(_4063_),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8311_ (.I(_4073_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8312_ (.I(_4062_),
    .Z(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8313_ (.A1(\reg_file.reg_storage[4][5] ),
    .A2(_4074_),
    .ZN(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8314_ (.A1(_3997_),
    .A2(_4068_),
    .B(_4075_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8315_ (.A1(\reg_file.reg_storage[4][6] ),
    .A2(_4074_),
    .ZN(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8316_ (.A1(_4000_),
    .A2(_4068_),
    .B(_4076_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8317_ (.I(_4067_),
    .Z(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8318_ (.A1(\reg_file.reg_storage[4][7] ),
    .A2(_4074_),
    .ZN(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8319_ (.A1(_4002_),
    .A2(_4077_),
    .B(_4078_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8320_ (.A1(\reg_file.reg_storage[4][8] ),
    .A2(_4074_),
    .ZN(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8321_ (.A1(_4005_),
    .A2(_4077_),
    .B(_4079_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8322_ (.I(_4062_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8323_ (.A1(\reg_file.reg_storage[4][9] ),
    .A2(_4080_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8324_ (.A1(_4007_),
    .A2(_4077_),
    .B(_4081_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8325_ (.A1(\reg_file.reg_storage[4][10] ),
    .A2(_4080_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8326_ (.A1(_4010_),
    .A2(_4077_),
    .B(_4082_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8327_ (.I(_4067_),
    .Z(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8328_ (.A1(\reg_file.reg_storage[4][11] ),
    .A2(_4080_),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8329_ (.A1(_4012_),
    .A2(_4083_),
    .B(_4084_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8330_ (.I(_4062_),
    .Z(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8331_ (.I0(\reg_file.reg_storage[4][12] ),
    .I1(_4015_),
    .S(_4085_),
    .Z(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8332_ (.I(_4086_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8333_ (.A1(\reg_file.reg_storage[4][13] ),
    .A2(_4080_),
    .ZN(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8334_ (.A1(_4018_),
    .A2(_4083_),
    .B(_4087_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8335_ (.I(_4066_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8336_ (.A1(\reg_file.reg_storage[4][14] ),
    .A2(_4088_),
    .ZN(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8337_ (.A1(_4020_),
    .A2(_4083_),
    .B(_4089_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8338_ (.A1(\reg_file.reg_storage[4][15] ),
    .A2(_4088_),
    .ZN(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8339_ (.A1(_4023_),
    .A2(_4083_),
    .B(_4090_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8340_ (.I0(\reg_file.reg_storage[4][16] ),
    .I1(_4025_),
    .S(_4085_),
    .Z(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8341_ (.I(_4091_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8342_ (.I(_4067_),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8343_ (.A1(\reg_file.reg_storage[4][17] ),
    .A2(_4088_),
    .ZN(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8344_ (.A1(_4027_),
    .A2(_4092_),
    .B(_4093_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8345_ (.A1(\reg_file.reg_storage[4][18] ),
    .A2(_4088_),
    .ZN(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8346_ (.A1(_4030_),
    .A2(_4092_),
    .B(_4094_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8347_ (.I(_4066_),
    .Z(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8348_ (.A1(\reg_file.reg_storage[4][19] ),
    .A2(_4095_),
    .ZN(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8349_ (.A1(_4032_),
    .A2(_4092_),
    .B(_4096_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8350_ (.I0(\reg_file.reg_storage[4][20] ),
    .I1(_4035_),
    .S(_4085_),
    .Z(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8351_ (.I(_4097_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8352_ (.I0(\reg_file.reg_storage[4][21] ),
    .I1(_4037_),
    .S(_4085_),
    .Z(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8353_ (.I(_4098_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8354_ (.I0(\reg_file.reg_storage[4][22] ),
    .I1(_4039_),
    .S(_4069_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8355_ (.I(_4099_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8356_ (.A1(\reg_file.reg_storage[4][23] ),
    .A2(_4095_),
    .ZN(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8357_ (.A1(_4041_),
    .A2(_4092_),
    .B(_4100_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8358_ (.I(_4063_),
    .Z(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8359_ (.A1(\reg_file.reg_storage[4][24] ),
    .A2(_4095_),
    .ZN(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8360_ (.A1(_4043_),
    .A2(_4101_),
    .B(_4102_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8361_ (.A1(\reg_file.reg_storage[4][25] ),
    .A2(_4095_),
    .ZN(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8362_ (.A1(_4046_),
    .A2(_4101_),
    .B(_4103_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8363_ (.I(_4066_),
    .Z(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8364_ (.A1(\reg_file.reg_storage[4][26] ),
    .A2(_4104_),
    .ZN(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8365_ (.A1(_4048_),
    .A2(_4101_),
    .B(_4105_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8366_ (.A1(\reg_file.reg_storage[4][27] ),
    .A2(_4104_),
    .ZN(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8367_ (.A1(_4051_),
    .A2(_4101_),
    .B(_4106_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8368_ (.A1(\reg_file.reg_storage[4][28] ),
    .A2(_4104_),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8369_ (.A1(_4053_),
    .A2(_4070_),
    .B(_4107_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8370_ (.I0(\reg_file.reg_storage[4][29] ),
    .I1(_4055_),
    .S(_4069_),
    .Z(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8371_ (.I(_4108_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8372_ (.I0(\reg_file.reg_storage[4][30] ),
    .I1(_4057_),
    .S(_4069_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8373_ (.I(_4109_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8374_ (.A1(\reg_file.reg_storage[4][31] ),
    .A2(_4104_),
    .ZN(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8375_ (.A1(_4059_),
    .A2(_4070_),
    .B(_4110_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8376_ (.A1(_3723_),
    .A2(_3827_),
    .ZN(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8377_ (.I(_4111_),
    .Z(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _8378_ (.I(_4112_),
    .Z(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8379_ (.I0(\reg_file.reg_storage[5][0] ),
    .I1(_3979_),
    .S(_4113_),
    .Z(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8380_ (.I(_4114_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8381_ (.I0(\reg_file.reg_storage[5][1] ),
    .I1(_3984_),
    .S(_4113_),
    .Z(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8382_ (.I(_4115_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8383_ (.I(_4111_),
    .Z(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8384_ (.I(_4116_),
    .Z(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8385_ (.I(_4117_),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8386_ (.I(_4111_),
    .Z(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8387_ (.I(_4119_),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8388_ (.A1(\reg_file.reg_storage[5][2] ),
    .A2(_4120_),
    .ZN(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8389_ (.A1(_3986_),
    .A2(_4118_),
    .B(_4121_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8390_ (.A1(\reg_file.reg_storage[5][3] ),
    .A2(_4120_),
    .ZN(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8391_ (.A1(_3993_),
    .A2(_4118_),
    .B(_4122_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8392_ (.I0(\reg_file.reg_storage[5][4] ),
    .I1(_3995_),
    .S(_4113_),
    .Z(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8393_ (.I(_4123_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8394_ (.I(_4112_),
    .Z(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8395_ (.A1(\reg_file.reg_storage[5][5] ),
    .A2(_4124_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8396_ (.A1(_3997_),
    .A2(_4118_),
    .B(_4125_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8397_ (.A1(\reg_file.reg_storage[5][6] ),
    .A2(_4124_),
    .ZN(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8398_ (.A1(_4000_),
    .A2(_4118_),
    .B(_4126_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8399_ (.I(_4117_),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8400_ (.A1(\reg_file.reg_storage[5][7] ),
    .A2(_4124_),
    .ZN(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8401_ (.A1(_4002_),
    .A2(_4127_),
    .B(_4128_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8402_ (.A1(\reg_file.reg_storage[5][8] ),
    .A2(_4124_),
    .ZN(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8403_ (.A1(_4005_),
    .A2(_4127_),
    .B(_4129_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8404_ (.I(_4112_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8405_ (.A1(\reg_file.reg_storage[5][9] ),
    .A2(_4130_),
    .ZN(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8406_ (.A1(_4007_),
    .A2(_4127_),
    .B(_4131_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8407_ (.A1(\reg_file.reg_storage[5][10] ),
    .A2(_4130_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8408_ (.A1(_4010_),
    .A2(_4127_),
    .B(_4132_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8409_ (.I(_4117_),
    .Z(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8410_ (.A1(\reg_file.reg_storage[5][11] ),
    .A2(_4130_),
    .ZN(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8411_ (.A1(_4012_),
    .A2(_4133_),
    .B(_4134_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8412_ (.I(_4112_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8413_ (.I0(\reg_file.reg_storage[5][12] ),
    .I1(_4015_),
    .S(_4135_),
    .Z(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8414_ (.I(_4136_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8415_ (.A1(\reg_file.reg_storage[5][13] ),
    .A2(_4130_),
    .ZN(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8416_ (.A1(_4018_),
    .A2(_4133_),
    .B(_4137_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8417_ (.I(_4116_),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8418_ (.A1(\reg_file.reg_storage[5][14] ),
    .A2(_4138_),
    .ZN(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8419_ (.A1(_4020_),
    .A2(_4133_),
    .B(_4139_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8420_ (.A1(\reg_file.reg_storage[5][15] ),
    .A2(_4138_),
    .ZN(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8421_ (.A1(_4023_),
    .A2(_4133_),
    .B(_4140_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8422_ (.I0(\reg_file.reg_storage[5][16] ),
    .I1(_4025_),
    .S(_4135_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8423_ (.I(_4141_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8424_ (.I(_4117_),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8425_ (.A1(\reg_file.reg_storage[5][17] ),
    .A2(_4138_),
    .ZN(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8426_ (.A1(_4027_),
    .A2(_4142_),
    .B(_4143_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8427_ (.A1(\reg_file.reg_storage[5][18] ),
    .A2(_4138_),
    .ZN(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8428_ (.A1(_4030_),
    .A2(_4142_),
    .B(_4144_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8429_ (.I(_4116_),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8430_ (.A1(\reg_file.reg_storage[5][19] ),
    .A2(_4145_),
    .ZN(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8431_ (.A1(_4032_),
    .A2(_4142_),
    .B(_4146_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8432_ (.I0(\reg_file.reg_storage[5][20] ),
    .I1(_4035_),
    .S(_4135_),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8433_ (.I(_4147_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8434_ (.I0(\reg_file.reg_storage[5][21] ),
    .I1(_4037_),
    .S(_4135_),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8435_ (.I(_4148_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8436_ (.I0(\reg_file.reg_storage[5][22] ),
    .I1(_4039_),
    .S(_4119_),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8437_ (.I(_4149_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8438_ (.A1(\reg_file.reg_storage[5][23] ),
    .A2(_4145_),
    .ZN(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8439_ (.A1(_4041_),
    .A2(_4142_),
    .B(_4150_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8440_ (.I(_4113_),
    .Z(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8441_ (.A1(\reg_file.reg_storage[5][24] ),
    .A2(_4145_),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8442_ (.A1(_4043_),
    .A2(_4151_),
    .B(_4152_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8443_ (.A1(\reg_file.reg_storage[5][25] ),
    .A2(_4145_),
    .ZN(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8444_ (.A1(_4046_),
    .A2(_4151_),
    .B(_4153_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8445_ (.I(_4116_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8446_ (.A1(\reg_file.reg_storage[5][26] ),
    .A2(_4154_),
    .ZN(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8447_ (.A1(_4048_),
    .A2(_4151_),
    .B(_4155_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8448_ (.A1(\reg_file.reg_storage[5][27] ),
    .A2(_4154_),
    .ZN(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8449_ (.A1(_4051_),
    .A2(_4151_),
    .B(_4156_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8450_ (.A1(\reg_file.reg_storage[5][28] ),
    .A2(_4154_),
    .ZN(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8451_ (.A1(_4053_),
    .A2(_4120_),
    .B(_4157_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8452_ (.I0(\reg_file.reg_storage[5][29] ),
    .I1(_4055_),
    .S(_4119_),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8453_ (.I(_4158_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8454_ (.I0(\reg_file.reg_storage[5][30] ),
    .I1(_4057_),
    .S(_4119_),
    .Z(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8455_ (.I(_4159_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8456_ (.A1(\reg_file.reg_storage[5][31] ),
    .A2(_4154_),
    .ZN(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8457_ (.A1(_4059_),
    .A2(_4120_),
    .B(_4160_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _8458_ (.A1(_3564_),
    .A2(_3321_),
    .A3(_3325_),
    .ZN(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8459_ (.I(_4161_),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _8460_ (.I(_4162_),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8461_ (.I0(\reg_file.reg_storage[12][0] ),
    .I1(_3979_),
    .S(_4163_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8462_ (.I(_4164_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8463_ (.I0(\reg_file.reg_storage[12][1] ),
    .I1(_3984_),
    .S(_4163_),
    .Z(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8464_ (.I(_4165_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8465_ (.I(_4161_),
    .Z(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8466_ (.I(_4166_),
    .Z(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8467_ (.I(_4167_),
    .Z(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8468_ (.I(_4161_),
    .Z(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8469_ (.I(_4169_),
    .Z(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8470_ (.A1(\reg_file.reg_storage[12][2] ),
    .A2(_4170_),
    .ZN(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8471_ (.A1(_3986_),
    .A2(_4168_),
    .B(_4171_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8472_ (.A1(\reg_file.reg_storage[12][3] ),
    .A2(_4170_),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8473_ (.A1(_3993_),
    .A2(_4168_),
    .B(_4172_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8474_ (.I0(\reg_file.reg_storage[12][4] ),
    .I1(_3995_),
    .S(_4163_),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8475_ (.I(_4173_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8476_ (.I(_4162_),
    .Z(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8477_ (.A1(\reg_file.reg_storage[12][5] ),
    .A2(_4174_),
    .ZN(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8478_ (.A1(_3997_),
    .A2(_4168_),
    .B(_4175_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8479_ (.A1(\reg_file.reg_storage[12][6] ),
    .A2(_4174_),
    .ZN(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8480_ (.A1(_4000_),
    .A2(_4168_),
    .B(_4176_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8481_ (.I(_4167_),
    .Z(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8482_ (.A1(\reg_file.reg_storage[12][7] ),
    .A2(_4174_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8483_ (.A1(_4002_),
    .A2(_4177_),
    .B(_4178_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8484_ (.A1(\reg_file.reg_storage[12][8] ),
    .A2(_4174_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8485_ (.A1(_4005_),
    .A2(_4177_),
    .B(_4179_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8486_ (.I(_4162_),
    .Z(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8487_ (.A1(\reg_file.reg_storage[12][9] ),
    .A2(_4180_),
    .ZN(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8488_ (.A1(_4007_),
    .A2(_4177_),
    .B(_4181_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8489_ (.A1(\reg_file.reg_storage[12][10] ),
    .A2(_4180_),
    .ZN(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8490_ (.A1(_4010_),
    .A2(_4177_),
    .B(_4182_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8491_ (.I(_4167_),
    .Z(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8492_ (.A1(\reg_file.reg_storage[12][11] ),
    .A2(_4180_),
    .ZN(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8493_ (.A1(_4012_),
    .A2(_4183_),
    .B(_4184_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8494_ (.I(_4162_),
    .Z(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8495_ (.I0(\reg_file.reg_storage[12][12] ),
    .I1(_4015_),
    .S(_4185_),
    .Z(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8496_ (.I(_4186_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8497_ (.A1(\reg_file.reg_storage[12][13] ),
    .A2(_4180_),
    .ZN(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8498_ (.A1(_4018_),
    .A2(_4183_),
    .B(_4187_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8499_ (.I(_4166_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8500_ (.A1(\reg_file.reg_storage[12][14] ),
    .A2(_4188_),
    .ZN(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8501_ (.A1(_4020_),
    .A2(_4183_),
    .B(_4189_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8502_ (.A1(\reg_file.reg_storage[12][15] ),
    .A2(_4188_),
    .ZN(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8503_ (.A1(_4023_),
    .A2(_4183_),
    .B(_4190_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8504_ (.I0(\reg_file.reg_storage[12][16] ),
    .I1(_4025_),
    .S(_4185_),
    .Z(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8505_ (.I(_4191_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8506_ (.I(_4167_),
    .Z(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8507_ (.A1(\reg_file.reg_storage[12][17] ),
    .A2(_4188_),
    .ZN(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8508_ (.A1(_4027_),
    .A2(_4192_),
    .B(_4193_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8509_ (.A1(\reg_file.reg_storage[12][18] ),
    .A2(_4188_),
    .ZN(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8510_ (.A1(_4030_),
    .A2(_4192_),
    .B(_4194_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8511_ (.I(_4166_),
    .Z(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8512_ (.A1(\reg_file.reg_storage[12][19] ),
    .A2(_4195_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8513_ (.A1(_4032_),
    .A2(_4192_),
    .B(_4196_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8514_ (.I0(\reg_file.reg_storage[12][20] ),
    .I1(_4035_),
    .S(_4185_),
    .Z(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8515_ (.I(_4197_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8516_ (.I0(\reg_file.reg_storage[12][21] ),
    .I1(_4037_),
    .S(_4185_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8517_ (.I(_4198_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8518_ (.I0(\reg_file.reg_storage[12][22] ),
    .I1(_4039_),
    .S(_4169_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8519_ (.I(_4199_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8520_ (.A1(\reg_file.reg_storage[12][23] ),
    .A2(_4195_),
    .ZN(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8521_ (.A1(_4041_),
    .A2(_4192_),
    .B(_4200_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8522_ (.I(_4163_),
    .Z(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8523_ (.A1(\reg_file.reg_storage[12][24] ),
    .A2(_4195_),
    .ZN(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8524_ (.A1(_4043_),
    .A2(_4201_),
    .B(_4202_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8525_ (.A1(\reg_file.reg_storage[12][25] ),
    .A2(_4195_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8526_ (.A1(_4046_),
    .A2(_4201_),
    .B(_4203_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8527_ (.I(_4166_),
    .Z(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8528_ (.A1(\reg_file.reg_storage[12][26] ),
    .A2(_4204_),
    .ZN(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8529_ (.A1(_4048_),
    .A2(_4201_),
    .B(_4205_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8530_ (.A1(\reg_file.reg_storage[12][27] ),
    .A2(_4204_),
    .ZN(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8531_ (.A1(_4051_),
    .A2(_4201_),
    .B(_4206_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8532_ (.A1(\reg_file.reg_storage[12][28] ),
    .A2(_4204_),
    .ZN(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8533_ (.A1(_4053_),
    .A2(_4170_),
    .B(_4207_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8534_ (.I0(\reg_file.reg_storage[12][29] ),
    .I1(_4055_),
    .S(_4169_),
    .Z(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8535_ (.I(_4208_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8536_ (.I0(\reg_file.reg_storage[12][30] ),
    .I1(_4057_),
    .S(_4169_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8537_ (.I(_4209_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8538_ (.A1(\reg_file.reg_storage[12][31] ),
    .A2(_4204_),
    .ZN(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8539_ (.A1(_4059_),
    .A2(_4170_),
    .B(_4210_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8540_ (.A1(_3618_),
    .A2(_3828_),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8541_ (.I(_4211_),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _8542_ (.I(_4212_),
    .Z(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8543_ (.I0(\reg_file.reg_storage[10][0] ),
    .I1(_3318_),
    .S(_4213_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8544_ (.I(_4214_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8545_ (.I0(\reg_file.reg_storage[10][1] ),
    .I1(_3336_),
    .S(_4213_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8546_ (.I(_4215_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8547_ (.I(_4211_),
    .Z(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8548_ (.I(_4216_),
    .Z(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8549_ (.I(_4217_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8550_ (.I(_4211_),
    .Z(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8551_ (.I(_4219_),
    .Z(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8552_ (.A1(\reg_file.reg_storage[10][2] ),
    .A2(_4220_),
    .ZN(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8553_ (.A1(_3730_),
    .A2(_4218_),
    .B(_4221_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8554_ (.A1(\reg_file.reg_storage[10][3] ),
    .A2(_4220_),
    .ZN(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8555_ (.A1(_3738_),
    .A2(_4218_),
    .B(_4222_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8556_ (.I0(\reg_file.reg_storage[10][4] ),
    .I1(_3368_),
    .S(_4213_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8557_ (.I(_4223_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8558_ (.I(_4212_),
    .Z(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8559_ (.A1(\reg_file.reg_storage[10][5] ),
    .A2(_4224_),
    .ZN(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8560_ (.A1(_3743_),
    .A2(_4218_),
    .B(_4225_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8561_ (.A1(\reg_file.reg_storage[10][6] ),
    .A2(_4224_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8562_ (.A1(_3747_),
    .A2(_4218_),
    .B(_4226_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8563_ (.I(_4217_),
    .Z(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8564_ (.A1(\reg_file.reg_storage[10][7] ),
    .A2(_4224_),
    .ZN(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8565_ (.A1(_3750_),
    .A2(_4227_),
    .B(_4228_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8566_ (.A1(\reg_file.reg_storage[10][8] ),
    .A2(_4224_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8567_ (.A1(_3754_),
    .A2(_4227_),
    .B(_4229_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8568_ (.I(_4212_),
    .Z(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8569_ (.A1(\reg_file.reg_storage[10][9] ),
    .A2(_4230_),
    .ZN(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8570_ (.A1(_3757_),
    .A2(_4227_),
    .B(_4231_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8571_ (.A1(\reg_file.reg_storage[10][10] ),
    .A2(_4230_),
    .ZN(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8572_ (.A1(_3761_),
    .A2(_4227_),
    .B(_4232_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8573_ (.I(_4217_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8574_ (.A1(\reg_file.reg_storage[10][11] ),
    .A2(_4230_),
    .ZN(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8575_ (.A1(_3764_),
    .A2(_4233_),
    .B(_4234_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8576_ (.I(_4212_),
    .Z(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8577_ (.I0(\reg_file.reg_storage[10][12] ),
    .I1(_3429_),
    .S(_4235_),
    .Z(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8578_ (.I(_4236_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8579_ (.A1(\reg_file.reg_storage[10][13] ),
    .A2(_4230_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8580_ (.A1(_3771_),
    .A2(_4233_),
    .B(_4237_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8581_ (.I(_4216_),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8582_ (.A1(\reg_file.reg_storage[10][14] ),
    .A2(_4238_),
    .ZN(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8583_ (.A1(_3774_),
    .A2(_4233_),
    .B(_4239_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8584_ (.A1(\reg_file.reg_storage[10][15] ),
    .A2(_4238_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8585_ (.A1(_3778_),
    .A2(_4233_),
    .B(_4240_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8586_ (.I0(\reg_file.reg_storage[10][16] ),
    .I1(_3459_),
    .S(_4235_),
    .Z(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8587_ (.I(_4241_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8588_ (.I(_4217_),
    .Z(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8589_ (.A1(\reg_file.reg_storage[10][17] ),
    .A2(_4238_),
    .ZN(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8590_ (.A1(_3783_),
    .A2(_4242_),
    .B(_4243_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8591_ (.A1(\reg_file.reg_storage[10][18] ),
    .A2(_4238_),
    .ZN(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8592_ (.A1(_3787_),
    .A2(_4242_),
    .B(_4244_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8593_ (.I(_4216_),
    .Z(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8594_ (.A1(\reg_file.reg_storage[10][19] ),
    .A2(_4245_),
    .ZN(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8595_ (.A1(_3790_),
    .A2(_4242_),
    .B(_4246_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8596_ (.I0(\reg_file.reg_storage[10][20] ),
    .I1(_3489_),
    .S(_4235_),
    .Z(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8597_ (.I(_4247_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8598_ (.I0(\reg_file.reg_storage[10][21] ),
    .I1(_3496_),
    .S(_4235_),
    .Z(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8599_ (.I(_4248_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8600_ (.I0(\reg_file.reg_storage[10][22] ),
    .I1(_3503_),
    .S(_4219_),
    .Z(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8601_ (.I(_4249_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8602_ (.A1(\reg_file.reg_storage[10][23] ),
    .A2(_4245_),
    .ZN(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8603_ (.A1(_3800_),
    .A2(_4242_),
    .B(_4250_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8604_ (.I(_4213_),
    .Z(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8605_ (.A1(\reg_file.reg_storage[10][24] ),
    .A2(_4245_),
    .ZN(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8606_ (.A1(_3803_),
    .A2(_4251_),
    .B(_4252_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8607_ (.A1(\reg_file.reg_storage[10][25] ),
    .A2(_4245_),
    .ZN(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8608_ (.A1(_3807_),
    .A2(_4251_),
    .B(_4253_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8609_ (.I(_4216_),
    .Z(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8610_ (.A1(\reg_file.reg_storage[10][26] ),
    .A2(_4254_),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8611_ (.A1(_3810_),
    .A2(_4251_),
    .B(_4255_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8612_ (.A1(\reg_file.reg_storage[10][27] ),
    .A2(_4254_),
    .ZN(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8613_ (.A1(_3814_),
    .A2(_4251_),
    .B(_4256_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8614_ (.A1(\reg_file.reg_storage[10][28] ),
    .A2(_4254_),
    .ZN(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8615_ (.A1(_3817_),
    .A2(_4220_),
    .B(_4257_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8616_ (.I0(\reg_file.reg_storage[10][29] ),
    .I1(_3550_),
    .S(_4219_),
    .Z(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8617_ (.I(_4258_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8618_ (.I0(\reg_file.reg_storage[10][30] ),
    .I1(_3556_),
    .S(_4219_),
    .Z(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8619_ (.I(_4259_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8620_ (.A1(\reg_file.reg_storage[10][31] ),
    .A2(_4254_),
    .ZN(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8621_ (.A1(_3824_),
    .A2(_4220_),
    .B(_4260_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8622_ (.A1(_3616_),
    .A2(_3322_),
    .A3(_3828_),
    .ZN(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8623_ (.I(_4261_),
    .Z(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _8624_ (.I(_4262_),
    .Z(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8625_ (.I0(\reg_file.reg_storage[2][0] ),
    .I1(_3318_),
    .S(_4263_),
    .Z(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8626_ (.I(_4264_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8627_ (.I0(\reg_file.reg_storage[2][1] ),
    .I1(_3336_),
    .S(_4263_),
    .Z(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8628_ (.I(_4265_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8629_ (.I(_4261_),
    .Z(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8630_ (.I(_4266_),
    .Z(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8631_ (.I(_4267_),
    .Z(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8632_ (.I(_4261_),
    .Z(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8633_ (.I(_4269_),
    .Z(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8634_ (.A1(\reg_file.reg_storage[2][2] ),
    .A2(_4270_),
    .ZN(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8635_ (.A1(_3730_),
    .A2(_4268_),
    .B(_4271_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8636_ (.A1(\reg_file.reg_storage[2][3] ),
    .A2(_4270_),
    .ZN(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8637_ (.A1(_3738_),
    .A2(_4268_),
    .B(_4272_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8638_ (.I0(\reg_file.reg_storage[2][4] ),
    .I1(_3368_),
    .S(_4263_),
    .Z(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8639_ (.I(_4273_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8640_ (.I(_4262_),
    .Z(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8641_ (.A1(\reg_file.reg_storage[2][5] ),
    .A2(_4274_),
    .ZN(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8642_ (.A1(_3743_),
    .A2(_4268_),
    .B(_4275_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8643_ (.A1(\reg_file.reg_storage[2][6] ),
    .A2(_4274_),
    .ZN(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8644_ (.A1(_3747_),
    .A2(_4268_),
    .B(_4276_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8645_ (.I(_4267_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8646_ (.A1(\reg_file.reg_storage[2][7] ),
    .A2(_4274_),
    .ZN(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8647_ (.A1(_3750_),
    .A2(_4277_),
    .B(_4278_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8648_ (.A1(\reg_file.reg_storage[2][8] ),
    .A2(_4274_),
    .ZN(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8649_ (.A1(_3754_),
    .A2(_4277_),
    .B(_4279_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8650_ (.I(_4262_),
    .Z(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8651_ (.A1(\reg_file.reg_storage[2][9] ),
    .A2(_4280_),
    .ZN(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8652_ (.A1(_3757_),
    .A2(_4277_),
    .B(_4281_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8653_ (.A1(\reg_file.reg_storage[2][10] ),
    .A2(_4280_),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8654_ (.A1(_3761_),
    .A2(_4277_),
    .B(_4282_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8655_ (.I(_4267_),
    .Z(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8656_ (.A1(\reg_file.reg_storage[2][11] ),
    .A2(_4280_),
    .ZN(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8657_ (.A1(_3764_),
    .A2(_4283_),
    .B(_4284_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8658_ (.I(_4262_),
    .Z(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8659_ (.I0(\reg_file.reg_storage[2][12] ),
    .I1(_3429_),
    .S(_4285_),
    .Z(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8660_ (.I(_4286_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8661_ (.A1(\reg_file.reg_storage[2][13] ),
    .A2(_4280_),
    .ZN(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8662_ (.A1(_3771_),
    .A2(_4283_),
    .B(_4287_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8663_ (.I(_4266_),
    .Z(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8664_ (.A1(\reg_file.reg_storage[2][14] ),
    .A2(_4288_),
    .ZN(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8665_ (.A1(_3774_),
    .A2(_4283_),
    .B(_4289_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8666_ (.A1(\reg_file.reg_storage[2][15] ),
    .A2(_4288_),
    .ZN(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8667_ (.A1(_3778_),
    .A2(_4283_),
    .B(_4290_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8668_ (.I0(\reg_file.reg_storage[2][16] ),
    .I1(_3459_),
    .S(_4285_),
    .Z(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8669_ (.I(_4291_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8670_ (.I(_4267_),
    .Z(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8671_ (.A1(\reg_file.reg_storage[2][17] ),
    .A2(_4288_),
    .ZN(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8672_ (.A1(_3783_),
    .A2(_4292_),
    .B(_4293_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8673_ (.A1(\reg_file.reg_storage[2][18] ),
    .A2(_4288_),
    .ZN(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8674_ (.A1(_3787_),
    .A2(_4292_),
    .B(_4294_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8675_ (.I(_4266_),
    .Z(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8676_ (.A1(\reg_file.reg_storage[2][19] ),
    .A2(_4295_),
    .ZN(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8677_ (.A1(_3790_),
    .A2(_4292_),
    .B(_4296_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8678_ (.I0(\reg_file.reg_storage[2][20] ),
    .I1(_3489_),
    .S(_4285_),
    .Z(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8679_ (.I(_4297_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8680_ (.I0(\reg_file.reg_storage[2][21] ),
    .I1(_3496_),
    .S(_4285_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8681_ (.I(_4298_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8682_ (.I0(\reg_file.reg_storage[2][22] ),
    .I1(_3503_),
    .S(_4269_),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8683_ (.I(_4299_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8684_ (.A1(\reg_file.reg_storage[2][23] ),
    .A2(_4295_),
    .ZN(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8685_ (.A1(_3800_),
    .A2(_4292_),
    .B(_4300_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8686_ (.I(_4263_),
    .Z(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8687_ (.A1(\reg_file.reg_storage[2][24] ),
    .A2(_4295_),
    .ZN(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8688_ (.A1(_3803_),
    .A2(_4301_),
    .B(_4302_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8689_ (.A1(\reg_file.reg_storage[2][25] ),
    .A2(_4295_),
    .ZN(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8690_ (.A1(_3807_),
    .A2(_4301_),
    .B(_4303_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8691_ (.I(_4266_),
    .Z(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8692_ (.A1(\reg_file.reg_storage[2][26] ),
    .A2(_4304_),
    .ZN(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8693_ (.A1(_3810_),
    .A2(_4301_),
    .B(_4305_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8694_ (.A1(\reg_file.reg_storage[2][27] ),
    .A2(_4304_),
    .ZN(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8695_ (.A1(_3814_),
    .A2(_4301_),
    .B(_4306_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8696_ (.A1(\reg_file.reg_storage[2][28] ),
    .A2(_4304_),
    .ZN(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8697_ (.A1(_3817_),
    .A2(_4270_),
    .B(_4307_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8698_ (.I0(\reg_file.reg_storage[2][29] ),
    .I1(_3550_),
    .S(_4269_),
    .Z(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8699_ (.I(_4308_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8700_ (.I0(\reg_file.reg_storage[2][30] ),
    .I1(_3556_),
    .S(_4269_),
    .Z(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8701_ (.I(_4309_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8702_ (.A1(\reg_file.reg_storage[2][31] ),
    .A2(_4304_),
    .ZN(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8703_ (.A1(_3824_),
    .A2(_4270_),
    .B(_4310_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8704_ (.A1(_3671_),
    .A2(_3827_),
    .ZN(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8705_ (.I(_4311_),
    .Z(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _8706_ (.I(_4312_),
    .Z(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8707_ (.I0(\reg_file.reg_storage[7][0] ),
    .I1(_3318_),
    .S(_4313_),
    .Z(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8708_ (.I(_4314_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8709_ (.I0(\reg_file.reg_storage[7][1] ),
    .I1(_3336_),
    .S(_4313_),
    .Z(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8710_ (.I(_4315_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8711_ (.I(_4311_),
    .Z(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8712_ (.I(_4316_),
    .Z(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8713_ (.I(_4317_),
    .Z(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8714_ (.I(_4311_),
    .Z(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8715_ (.I(_4319_),
    .Z(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8716_ (.A1(\reg_file.reg_storage[7][2] ),
    .A2(_4320_),
    .ZN(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8717_ (.A1(_3730_),
    .A2(_4318_),
    .B(_4321_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8718_ (.A1(\reg_file.reg_storage[7][3] ),
    .A2(_4320_),
    .ZN(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8719_ (.A1(_3738_),
    .A2(_4318_),
    .B(_4322_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8720_ (.I0(\reg_file.reg_storage[7][4] ),
    .I1(_3368_),
    .S(_4313_),
    .Z(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8721_ (.I(_4323_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8722_ (.I(_4312_),
    .Z(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8723_ (.A1(\reg_file.reg_storage[7][5] ),
    .A2(_4324_),
    .ZN(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8724_ (.A1(_3743_),
    .A2(_4318_),
    .B(_4325_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8725_ (.A1(\reg_file.reg_storage[7][6] ),
    .A2(_4324_),
    .ZN(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8726_ (.A1(_3747_),
    .A2(_4318_),
    .B(_4326_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8727_ (.I(_4317_),
    .Z(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8728_ (.A1(\reg_file.reg_storage[7][7] ),
    .A2(_4324_),
    .ZN(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8729_ (.A1(_3750_),
    .A2(_4327_),
    .B(_4328_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8730_ (.A1(\reg_file.reg_storage[7][8] ),
    .A2(_4324_),
    .ZN(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8731_ (.A1(_3754_),
    .A2(_4327_),
    .B(_4329_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8732_ (.I(_4312_),
    .Z(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8733_ (.A1(\reg_file.reg_storage[7][9] ),
    .A2(_4330_),
    .ZN(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8734_ (.A1(_3757_),
    .A2(_4327_),
    .B(_4331_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8735_ (.A1(\reg_file.reg_storage[7][10] ),
    .A2(_4330_),
    .ZN(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8736_ (.A1(_3761_),
    .A2(_4327_),
    .B(_4332_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8737_ (.I(_4317_),
    .Z(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8738_ (.A1(\reg_file.reg_storage[7][11] ),
    .A2(_4330_),
    .ZN(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8739_ (.A1(_3764_),
    .A2(_4333_),
    .B(_4334_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _8740_ (.I(_4312_),
    .Z(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8741_ (.I0(\reg_file.reg_storage[7][12] ),
    .I1(_3429_),
    .S(_4335_),
    .Z(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8742_ (.I(_4336_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8743_ (.A1(\reg_file.reg_storage[7][13] ),
    .A2(_4330_),
    .ZN(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8744_ (.A1(_3771_),
    .A2(_4333_),
    .B(_4337_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8745_ (.I(_4316_),
    .Z(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8746_ (.A1(\reg_file.reg_storage[7][14] ),
    .A2(_4338_),
    .ZN(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8747_ (.A1(_3774_),
    .A2(_4333_),
    .B(_4339_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8748_ (.A1(\reg_file.reg_storage[7][15] ),
    .A2(_4338_),
    .ZN(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8749_ (.A1(_3778_),
    .A2(_4333_),
    .B(_4340_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8750_ (.I0(\reg_file.reg_storage[7][16] ),
    .I1(_3459_),
    .S(_4335_),
    .Z(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8751_ (.I(_4341_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8752_ (.I(_4317_),
    .Z(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8753_ (.A1(\reg_file.reg_storage[7][17] ),
    .A2(_4338_),
    .ZN(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8754_ (.A1(_3783_),
    .A2(_4342_),
    .B(_4343_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8755_ (.A1(\reg_file.reg_storage[7][18] ),
    .A2(_4338_),
    .ZN(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8756_ (.A1(_3787_),
    .A2(_4342_),
    .B(_4344_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8757_ (.I(_4316_),
    .Z(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8758_ (.A1(\reg_file.reg_storage[7][19] ),
    .A2(_4345_),
    .ZN(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8759_ (.A1(_3790_),
    .A2(_4342_),
    .B(_4346_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8760_ (.I0(\reg_file.reg_storage[7][20] ),
    .I1(_3489_),
    .S(_4335_),
    .Z(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8761_ (.I(_4347_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8762_ (.I0(\reg_file.reg_storage[7][21] ),
    .I1(_3496_),
    .S(_4335_),
    .Z(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8763_ (.I(_4348_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8764_ (.I0(\reg_file.reg_storage[7][22] ),
    .I1(_3503_),
    .S(_4319_),
    .Z(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8765_ (.I(_4349_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8766_ (.A1(\reg_file.reg_storage[7][23] ),
    .A2(_4345_),
    .ZN(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8767_ (.A1(_3800_),
    .A2(_4342_),
    .B(_4350_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8768_ (.I(_4313_),
    .Z(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8769_ (.A1(\reg_file.reg_storage[7][24] ),
    .A2(_4345_),
    .ZN(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8770_ (.A1(_3803_),
    .A2(_4351_),
    .B(_4352_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8771_ (.A1(\reg_file.reg_storage[7][25] ),
    .A2(_4345_),
    .ZN(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8772_ (.A1(_3807_),
    .A2(_4351_),
    .B(_4353_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8773_ (.I(_4316_),
    .Z(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8774_ (.A1(\reg_file.reg_storage[7][26] ),
    .A2(_4354_),
    .ZN(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8775_ (.A1(_3810_),
    .A2(_4351_),
    .B(_4355_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8776_ (.A1(\reg_file.reg_storage[7][27] ),
    .A2(_4354_),
    .ZN(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8777_ (.A1(_3814_),
    .A2(_4351_),
    .B(_4356_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8778_ (.A1(\reg_file.reg_storage[7][28] ),
    .A2(_4354_),
    .ZN(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8779_ (.A1(_3817_),
    .A2(_4320_),
    .B(_4357_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8780_ (.I0(\reg_file.reg_storage[7][29] ),
    .I1(_3550_),
    .S(_4319_),
    .Z(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8781_ (.I(_4358_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8782_ (.I0(\reg_file.reg_storage[7][30] ),
    .I1(_3556_),
    .S(_4319_),
    .Z(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8783_ (.I(_4359_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8784_ (.A1(\reg_file.reg_storage[7][31] ),
    .A2(_4354_),
    .ZN(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8785_ (.A1(_3824_),
    .A2(_4320_),
    .B(_4360_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8786_ (.D(_0000_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8787_ (.D(_0001_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8788_ (.D(_0002_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8789_ (.D(_0003_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8790_ (.D(_0004_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8791_ (.D(_0005_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8792_ (.D(_0006_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8793_ (.D(_0007_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8794_ (.D(_0008_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8795_ (.D(_0009_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8796_ (.D(_0010_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8797_ (.D(_0011_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8798_ (.D(_0012_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8799_ (.D(_0013_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8800_ (.D(_0014_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8801_ (.D(_0015_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8802_ (.D(_0016_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[14][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _8803_ (.D(_0017_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8804_ (.D(_0018_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8805_ (.D(_0019_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8806_ (.D(_0020_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8807_ (.D(_0021_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8808_ (.D(_0022_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8809_ (.D(_0023_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8810_ (.D(_0024_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8811_ (.D(_0025_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8812_ (.D(_0026_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8813_ (.D(_0027_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8814_ (.D(_0028_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8815_ (.D(_0029_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[14][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8816_ (.D(_0030_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[14][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8817_ (.D(_0031_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[14][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8818_ (.D(_0032_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8819_ (.D(_0033_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8820_ (.D(_0034_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8821_ (.D(_0035_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8822_ (.D(_0036_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8823_ (.D(_0037_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8824_ (.D(_0038_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8825_ (.D(_0039_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8826_ (.D(_0040_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8827_ (.D(_0041_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8828_ (.D(_0042_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8829_ (.D(_0043_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8830_ (.D(_0044_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8831_ (.D(_0045_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8832_ (.D(_0046_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8833_ (.D(_0047_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8834_ (.D(_0048_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8835_ (.D(_0049_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8836_ (.D(_0050_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8837_ (.D(_0051_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8838_ (.D(_0052_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8839_ (.D(_0053_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8840_ (.D(_0054_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8841_ (.D(_0055_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8842_ (.D(_0056_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8843_ (.D(_0057_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8844_ (.D(_0058_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8845_ (.D(_0059_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8846_ (.D(_0060_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8847_ (.D(_0061_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[13][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8848_ (.D(_0062_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[13][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8849_ (.D(_0063_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[13][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8850_ (.D(_0064_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8851_ (.D(_0065_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8852_ (.D(_0066_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8853_ (.D(_0067_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8854_ (.D(_0068_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8855_ (.D(_0069_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8856_ (.D(_0070_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8857_ (.D(_0071_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8858_ (.D(_0072_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8859_ (.D(_0073_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8860_ (.D(_0074_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8861_ (.D(_0075_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8862_ (.D(_0076_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8863_ (.D(_0077_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8864_ (.D(_0078_),
    .CLK(clknet_leaf_78_clk),
    .Q(\reg_file.reg_storage[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8865_ (.D(_0079_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8866_ (.D(_0080_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8867_ (.D(_0081_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8868_ (.D(_0082_),
    .CLK(clknet_leaf_77_clk),
    .Q(\reg_file.reg_storage[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8869_ (.D(_0083_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8870_ (.D(_0084_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8871_ (.D(_0085_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8872_ (.D(_0086_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8873_ (.D(_0087_),
    .CLK(clknet_leaf_75_clk),
    .Q(\reg_file.reg_storage[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8874_ (.D(_0088_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8875_ (.D(_0089_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8876_ (.D(_0090_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8877_ (.D(_0091_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8878_ (.D(_0092_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8879_ (.D(_0093_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[8][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8880_ (.D(_0094_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[8][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8881_ (.D(_0095_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[8][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8882_ (.D(_0096_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8883_ (.D(_0097_),
    .CLK(clknet_leaf_107_clk),
    .Q(\reg_file.reg_storage[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8884_ (.D(_0098_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8885_ (.D(_0099_),
    .CLK(clknet_leaf_8_clk),
    .Q(\reg_file.reg_storage[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8886_ (.D(_0100_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8887_ (.D(_0101_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8888_ (.D(_0102_),
    .CLK(clknet_leaf_6_clk),
    .Q(\reg_file.reg_storage[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8889_ (.D(_0103_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8890_ (.D(_0104_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8891_ (.D(_0105_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8892_ (.D(_0106_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8893_ (.D(_0107_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8894_ (.D(_0108_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8895_ (.D(_0109_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8896_ (.D(_0110_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8897_ (.D(_0111_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8898_ (.D(_0112_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[11][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8899_ (.D(_0113_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8900_ (.D(_0114_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8901_ (.D(_0115_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[11][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8902_ (.D(_0116_),
    .CLK(clknet_leaf_98_clk),
    .Q(\reg_file.reg_storage[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8903_ (.D(_0117_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[11][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8904_ (.D(_0118_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8905_ (.D(_0119_),
    .CLK(clknet_leaf_76_clk),
    .Q(\reg_file.reg_storage[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8906_ (.D(_0120_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8907_ (.D(_0121_),
    .CLK(clknet_leaf_74_clk),
    .Q(\reg_file.reg_storage[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8908_ (.D(_0122_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[11][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8909_ (.D(_0123_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8910_ (.D(_0124_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8911_ (.D(_0125_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[11][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8912_ (.D(_0126_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[11][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8913_ (.D(_0127_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[11][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8914_ (.D(_0128_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8915_ (.D(_0129_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8916_ (.D(_0130_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8917_ (.D(_0131_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8918_ (.D(_0132_),
    .CLK(clknet_leaf_0_clk),
    .Q(\reg_file.reg_storage[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8919_ (.D(_0133_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8920_ (.D(_0134_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8921_ (.D(_0135_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8922_ (.D(_0136_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8923_ (.D(_0137_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8924_ (.D(_0138_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8925_ (.D(_0139_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8926_ (.D(_0140_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8927_ (.D(_0141_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8928_ (.D(_0142_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8929_ (.D(_0143_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8930_ (.D(_0144_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[9][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8931_ (.D(_0145_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8932_ (.D(_0146_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8933_ (.D(_0147_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8934_ (.D(_0148_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8935_ (.D(_0149_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8936_ (.D(_0150_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8937_ (.D(_0151_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8938_ (.D(_0152_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8939_ (.D(_0153_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8940_ (.D(_0154_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8941_ (.D(_0155_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8942_ (.D(_0156_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[9][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8943_ (.D(_0157_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[9][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8944_ (.D(_0158_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[9][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8945_ (.D(_0159_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[9][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8946_ (.D(_0160_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8947_ (.D(_0161_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8948_ (.D(_0162_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8949_ (.D(_0163_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8950_ (.D(_0164_),
    .CLK(clknet_leaf_2_clk),
    .Q(\reg_file.reg_storage[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8951_ (.D(_0165_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8952_ (.D(_0166_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8953_ (.D(_0167_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8954_ (.D(_0168_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8955_ (.D(_0169_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8956_ (.D(_0170_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8957_ (.D(_0171_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8958_ (.D(_0172_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8959_ (.D(_0173_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8960_ (.D(_0174_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8961_ (.D(_0175_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8962_ (.D(_0176_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[6][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8963_ (.D(_0177_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[6][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8964_ (.D(_0178_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8965_ (.D(_0179_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[6][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8966_ (.D(_0180_),
    .CLK(clknet_leaf_90_clk),
    .Q(\reg_file.reg_storage[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8967_ (.D(_0181_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8968_ (.D(_0182_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8969_ (.D(_0183_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8970_ (.D(_0184_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8971_ (.D(_0185_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8972_ (.D(_0186_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8973_ (.D(_0187_),
    .CLK(clknet_leaf_63_clk),
    .Q(\reg_file.reg_storage[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8974_ (.D(_0188_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8975_ (.D(_0189_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[6][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8976_ (.D(_0190_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[6][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8977_ (.D(_0191_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[6][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8978_ (.D(_0192_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8979_ (.D(_0193_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _8980_ (.D(_0194_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8981_ (.D(_0195_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8982_ (.D(_0196_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8983_ (.D(_0197_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8984_ (.D(_0198_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8985_ (.D(_0199_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8986_ (.D(_0200_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8987_ (.D(_0201_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8988_ (.D(_0202_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8989_ (.D(_0203_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8990_ (.D(_0204_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8991_ (.D(_0205_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8992_ (.D(_0206_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8993_ (.D(_0207_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8994_ (.D(_0208_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8995_ (.D(_0209_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8996_ (.D(_0210_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8997_ (.D(_0211_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8998_ (.D(_0212_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8999_ (.D(_0213_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9000_ (.D(_0214_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9001_ (.D(_0215_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9002_ (.D(_0216_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9003_ (.D(_0217_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9004_ (.D(_0218_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9005_ (.D(_0219_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9006_ (.D(_0220_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[1][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9007_ (.D(_0221_),
    .CLK(clknet_leaf_39_clk),
    .Q(\reg_file.reg_storage[1][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9008_ (.D(_0222_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[1][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9009_ (.D(_0223_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[1][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9010_ (.D(_0224_),
    .CLK(clknet_leaf_4_clk),
    .Q(\reg_file.reg_storage[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9011_ (.D(_0225_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9012_ (.D(_0226_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9013_ (.D(_0227_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9014_ (.D(_0228_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9015_ (.D(_0229_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9016_ (.D(_0230_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9017_ (.D(_0231_),
    .CLK(clknet_leaf_20_clk),
    .Q(\reg_file.reg_storage[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9018_ (.D(_0232_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9019_ (.D(_0233_),
    .CLK(clknet_leaf_19_clk),
    .Q(\reg_file.reg_storage[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9020_ (.D(_0234_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9021_ (.D(_0235_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9022_ (.D(_0236_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9023_ (.D(_0237_),
    .CLK(clknet_leaf_54_clk),
    .Q(\reg_file.reg_storage[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9024_ (.D(_0238_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9025_ (.D(_0239_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9026_ (.D(_0240_),
    .CLK(clknet_leaf_88_clk),
    .Q(\reg_file.reg_storage[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9027_ (.D(_0241_),
    .CLK(clknet_leaf_53_clk),
    .Q(\reg_file.reg_storage[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9028_ (.D(_0242_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9029_ (.D(_0243_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9030_ (.D(_0244_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9031_ (.D(_0245_),
    .CLK(clknet_leaf_92_clk),
    .Q(\reg_file.reg_storage[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9032_ (.D(_0246_),
    .CLK(clknet_leaf_31_clk),
    .Q(\reg_file.reg_storage[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9033_ (.D(_0247_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9034_ (.D(_0248_),
    .CLK(clknet_leaf_63_clk),
    .Q(\reg_file.reg_storage[3][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9035_ (.D(_0249_),
    .CLK(clknet_leaf_57_clk),
    .Q(\reg_file.reg_storage[3][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9036_ (.D(_0250_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[3][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9037_ (.D(_0251_),
    .CLK(clknet_leaf_52_clk),
    .Q(\reg_file.reg_storage[3][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9038_ (.D(_0252_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9039_ (.D(_0253_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[3][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9040_ (.D(_0254_),
    .CLK(clknet_leaf_40_clk),
    .Q(\reg_file.reg_storage[3][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9041_ (.D(_0255_),
    .CLK(clknet_leaf_50_clk),
    .Q(\reg_file.reg_storage[3][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9042_ (.D(_0256_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9043_ (.D(_0257_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9044_ (.D(_0258_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9045_ (.D(_0259_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9046_ (.D(_0260_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9047_ (.D(_0261_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9048_ (.D(_0262_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9049_ (.D(_0263_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9050_ (.D(_0264_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9051_ (.D(_0265_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9052_ (.D(_0266_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9053_ (.D(_0267_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9054_ (.D(_0268_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9055_ (.D(_0269_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9056_ (.D(_0270_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9057_ (.D(_0271_),
    .CLK(clknet_leaf_82_clk),
    .Q(\reg_file.reg_storage[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9058_ (.D(_0272_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[15][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9059_ (.D(_0273_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9060_ (.D(_0274_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[15][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9061_ (.D(_0275_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[15][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9062_ (.D(_0276_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9063_ (.D(_0277_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9064_ (.D(_0278_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9065_ (.D(_0279_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9066_ (.D(_0280_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9067_ (.D(_0281_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9068_ (.D(_0282_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9069_ (.D(_0283_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9070_ (.D(_0284_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9071_ (.D(_0285_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[15][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9072_ (.D(_0286_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[15][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9073_ (.D(_0287_),
    .CLK(clknet_leaf_43_clk),
    .Q(\reg_file.reg_storage[15][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9074_ (.D(_0288_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9075_ (.D(_0289_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9076_ (.D(_0290_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9077_ (.D(_0291_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9078_ (.D(_0292_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9079_ (.D(_0293_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9080_ (.D(_0294_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9081_ (.D(_0295_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9082_ (.D(_0296_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9083_ (.D(_0297_),
    .CLK(clknet_leaf_14_clk),
    .Q(\reg_file.reg_storage[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9084_ (.D(_0298_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9085_ (.D(_0299_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9086_ (.D(_0300_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9087_ (.D(_0301_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9088_ (.D(_0302_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9089_ (.D(_0303_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9090_ (.D(_0304_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9091_ (.D(_0305_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9092_ (.D(_0306_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9093_ (.D(_0307_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9094_ (.D(_0308_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[4][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9095_ (.D(_0309_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9096_ (.D(_0310_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[4][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9097_ (.D(_0311_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9098_ (.D(_0312_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9099_ (.D(_0313_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9100_ (.D(_0314_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9101_ (.D(_0315_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[4][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9102_ (.D(_0316_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9103_ (.D(_0317_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[4][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9104_ (.D(_0318_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[4][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9105_ (.D(_0319_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[4][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9106_ (.D(_0320_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9107_ (.D(_0321_),
    .CLK(clknet_leaf_106_clk),
    .Q(\reg_file.reg_storage[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9108_ (.D(_0322_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9109_ (.D(_0323_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9110_ (.D(_0324_),
    .CLK(clknet_leaf_104_clk),
    .Q(\reg_file.reg_storage[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9111_ (.D(_0325_),
    .CLK(clknet_leaf_10_clk),
    .Q(\reg_file.reg_storage[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9112_ (.D(_0326_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9113_ (.D(_0327_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9114_ (.D(_0328_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9115_ (.D(_0329_),
    .CLK(clknet_leaf_12_clk),
    .Q(\reg_file.reg_storage[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9116_ (.D(_0330_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9117_ (.D(_0331_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9118_ (.D(_0332_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9119_ (.D(_0333_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9120_ (.D(_0334_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9121_ (.D(_0335_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9122_ (.D(_0336_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9123_ (.D(_0337_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9124_ (.D(_0338_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9125_ (.D(_0339_),
    .CLK(clknet_leaf_71_clk),
    .Q(\reg_file.reg_storage[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9126_ (.D(_0340_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9127_ (.D(_0341_),
    .CLK(clknet_leaf_100_clk),
    .Q(\reg_file.reg_storage[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9128_ (.D(_0342_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9129_ (.D(_0343_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9130_ (.D(_0344_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9131_ (.D(_0345_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9132_ (.D(_0346_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9133_ (.D(_0347_),
    .CLK(clknet_leaf_66_clk),
    .Q(\reg_file.reg_storage[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9134_ (.D(_0348_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9135_ (.D(_0349_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[5][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9136_ (.D(_0350_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[5][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9137_ (.D(_0351_),
    .CLK(clknet_leaf_45_clk),
    .Q(\reg_file.reg_storage[5][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9138_ (.D(_0352_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9139_ (.D(_0353_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9140_ (.D(_0354_),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\reg_file.reg_storage[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9141_ (.D(_0355_),
    .CLK(clknet_leaf_7_clk),
    .Q(\reg_file.reg_storage[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9142_ (.D(_0356_),
    .CLK(clknet_leaf_105_clk),
    .Q(\reg_file.reg_storage[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9143_ (.D(_0357_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9144_ (.D(_0358_),
    .CLK(clknet_leaf_9_clk),
    .Q(\reg_file.reg_storage[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9145_ (.D(_0359_),
    .CLK(clknet_leaf_11_clk),
    .Q(\reg_file.reg_storage[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9146_ (.D(_0360_),
    .CLK(clknet_leaf_15_clk),
    .Q(\reg_file.reg_storage[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9147_ (.D(_0361_),
    .CLK(clknet_leaf_91_clk),
    .Q(\reg_file.reg_storage[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9148_ (.D(_0362_),
    .CLK(clknet_leaf_89_clk),
    .Q(\reg_file.reg_storage[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9149_ (.D(_0363_),
    .CLK(clknet_leaf_86_clk),
    .Q(\reg_file.reg_storage[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9150_ (.D(_0364_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9151_ (.D(_0365_),
    .CLK(clknet_leaf_87_clk),
    .Q(\reg_file.reg_storage[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9152_ (.D(_0366_),
    .CLK(clknet_leaf_81_clk),
    .Q(\reg_file.reg_storage[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9153_ (.D(_0367_),
    .CLK(clknet_leaf_80_clk),
    .Q(\reg_file.reg_storage[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9154_ (.D(_0368_),
    .CLK(clknet_leaf_96_clk),
    .Q(\reg_file.reg_storage[12][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9155_ (.D(_0369_),
    .CLK(clknet_leaf_79_clk),
    .Q(\reg_file.reg_storage[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9156_ (.D(_0370_),
    .CLK(clknet_leaf_70_clk),
    .Q(\reg_file.reg_storage[12][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9157_ (.D(_0371_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[12][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9158_ (.D(_0372_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[12][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9159_ (.D(_0373_),
    .CLK(clknet_leaf_99_clk),
    .Q(\reg_file.reg_storage[12][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9160_ (.D(_0374_),
    .CLK(clknet_leaf_30_clk),
    .Q(\reg_file.reg_storage[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9161_ (.D(_0375_),
    .CLK(clknet_leaf_73_clk),
    .Q(\reg_file.reg_storage[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9162_ (.D(_0376_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[12][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9163_ (.D(_0377_),
    .CLK(clknet_leaf_72_clk),
    .Q(\reg_file.reg_storage[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9164_ (.D(_0378_),
    .CLK(clknet_leaf_46_clk),
    .Q(\reg_file.reg_storage[12][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9165_ (.D(_0379_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9166_ (.D(_0380_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9167_ (.D(_0381_),
    .CLK(clknet_leaf_38_clk),
    .Q(\reg_file.reg_storage[12][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9168_ (.D(_0382_),
    .CLK(clknet_leaf_37_clk),
    .Q(\reg_file.reg_storage[12][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9169_ (.D(_0383_),
    .CLK(clknet_leaf_44_clk),
    .Q(\reg_file.reg_storage[12][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9170_ (.D(_0384_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9171_ (.D(_0385_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9172_ (.D(_0386_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9173_ (.D(_0387_),
    .CLK(clknet_leaf_28_clk),
    .Q(\reg_file.reg_storage[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9174_ (.D(_0388_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9175_ (.D(_0389_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9176_ (.D(_0390_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9177_ (.D(_0391_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9178_ (.D(_0392_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9179_ (.D(_0393_),
    .CLK(clknet_leaf_13_clk),
    .Q(\reg_file.reg_storage[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9180_ (.D(_0394_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9181_ (.D(_0395_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9182_ (.D(_0396_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9183_ (.D(_0397_),
    .CLK(clknet_leaf_85_clk),
    .Q(\reg_file.reg_storage[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9184_ (.D(_0398_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9185_ (.D(_0399_),
    .CLK(clknet_leaf_83_clk),
    .Q(\reg_file.reg_storage[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9186_ (.D(_0400_),
    .CLK(clknet_leaf_97_clk),
    .Q(\reg_file.reg_storage[10][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9187_ (.D(_0401_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9188_ (.D(_0402_),
    .CLK(clknet_leaf_60_clk),
    .Q(\reg_file.reg_storage[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9189_ (.D(_0403_),
    .CLK(clknet_leaf_69_clk),
    .Q(\reg_file.reg_storage[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9190_ (.D(_0404_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[10][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9191_ (.D(_0405_),
    .CLK(clknet_leaf_103_clk),
    .Q(\reg_file.reg_storage[10][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9192_ (.D(_0406_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[10][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9193_ (.D(_0407_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[10][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9194_ (.D(_0408_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9195_ (.D(_0409_),
    .CLK(clknet_leaf_68_clk),
    .Q(\reg_file.reg_storage[10][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9196_ (.D(_0410_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[10][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9197_ (.D(_0411_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9198_ (.D(_0412_),
    .CLK(clknet_leaf_41_clk),
    .Q(\reg_file.reg_storage[10][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9199_ (.D(_0413_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[10][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9200_ (.D(_0414_),
    .CLK(clknet_leaf_35_clk),
    .Q(\reg_file.reg_storage[10][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9201_ (.D(_0415_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[10][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9202_ (.D(_0416_),
    .CLK(clknet_leaf_3_clk),
    .Q(\reg_file.reg_storage[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9203_ (.D(_0417_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9204_ (.D(_0418_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9205_ (.D(_0419_),
    .CLK(clknet_leaf_26_clk),
    .Q(\reg_file.reg_storage[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9206_ (.D(_0420_),
    .CLK(clknet_leaf_5_clk),
    .Q(\reg_file.reg_storage[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9207_ (.D(_0421_),
    .CLK(clknet_leaf_27_clk),
    .Q(\reg_file.reg_storage[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9208_ (.D(_0422_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9209_ (.D(_0423_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9210_ (.D(_0424_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9211_ (.D(_0425_),
    .CLK(clknet_leaf_18_clk),
    .Q(\reg_file.reg_storage[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9212_ (.D(_0426_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9213_ (.D(_0427_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9214_ (.D(_0428_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9215_ (.D(_0429_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9216_ (.D(_0430_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9217_ (.D(_0431_),
    .CLK(clknet_leaf_56_clk),
    .Q(\reg_file.reg_storage[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9218_ (.D(_0432_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9219_ (.D(_0433_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9220_ (.D(_0434_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9221_ (.D(_0435_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9222_ (.D(_0436_),
    .CLK(clknet_leaf_94_clk),
    .Q(\reg_file.reg_storage[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9223_ (.D(_0437_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9224_ (.D(_0438_),
    .CLK(clknet_leaf_29_clk),
    .Q(\reg_file.reg_storage[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9225_ (.D(_0439_),
    .CLK(clknet_leaf_62_clk),
    .Q(\reg_file.reg_storage[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9226_ (.D(_0440_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9227_ (.D(_0441_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9228_ (.D(_0442_),
    .CLK(clknet_leaf_47_clk),
    .Q(\reg_file.reg_storage[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9229_ (.D(_0443_),
    .CLK(clknet_leaf_48_clk),
    .Q(\reg_file.reg_storage[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9230_ (.D(_0444_),
    .CLK(clknet_leaf_51_clk),
    .Q(\reg_file.reg_storage[2][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9231_ (.D(_0445_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[2][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9232_ (.D(_0446_),
    .CLK(clknet_leaf_32_clk),
    .Q(\reg_file.reg_storage[2][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9233_ (.D(_0447_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[2][31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9234_ (.D(_0448_),
    .CLK(clknet_leaf_102_clk),
    .Q(\reg_file.reg_storage[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9235_ (.D(_0449_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9236_ (.D(_0450_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9237_ (.D(_0451_),
    .CLK(clknet_leaf_25_clk),
    .Q(\reg_file.reg_storage[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9238_ (.D(_0452_),
    .CLK(clknet_leaf_1_clk),
    .Q(\reg_file.reg_storage[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9239_ (.D(_0453_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9240_ (.D(_0454_),
    .CLK(clknet_leaf_23_clk),
    .Q(\reg_file.reg_storage[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9241_ (.D(_0455_),
    .CLK(clknet_leaf_21_clk),
    .Q(\reg_file.reg_storage[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9242_ (.D(_0456_),
    .CLK(clknet_leaf_22_clk),
    .Q(\reg_file.reg_storage[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9243_ (.D(_0457_),
    .CLK(clknet_leaf_17_clk),
    .Q(\reg_file.reg_storage[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9244_ (.D(_0458_),
    .CLK(clknet_leaf_16_clk),
    .Q(\reg_file.reg_storage[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9245_ (.D(_0459_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9246_ (.D(_0460_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9247_ (.D(_0461_),
    .CLK(clknet_leaf_55_clk),
    .Q(\reg_file.reg_storage[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9248_ (.D(_0462_),
    .CLK(clknet_leaf_84_clk),
    .Q(\reg_file.reg_storage[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9249_ (.D(_0463_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9250_ (.D(_0464_),
    .CLK(clknet_leaf_95_clk),
    .Q(\reg_file.reg_storage[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9251_ (.D(_0465_),
    .CLK(clknet_leaf_58_clk),
    .Q(\reg_file.reg_storage[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9252_ (.D(_0466_),
    .CLK(clknet_leaf_59_clk),
    .Q(\reg_file.reg_storage[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9253_ (.D(_0467_),
    .CLK(clknet_leaf_64_clk),
    .Q(\reg_file.reg_storage[7][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9254_ (.D(_0468_),
    .CLK(clknet_leaf_93_clk),
    .Q(\reg_file.reg_storage[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9255_ (.D(_0469_),
    .CLK(clknet_leaf_101_clk),
    .Q(\reg_file.reg_storage[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9256_ (.D(_0470_),
    .CLK(clknet_leaf_33_clk),
    .Q(\reg_file.reg_storage[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9257_ (.D(_0471_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9258_ (.D(_0472_),
    .CLK(clknet_leaf_67_clk),
    .Q(\reg_file.reg_storage[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9259_ (.D(_0473_),
    .CLK(clknet_leaf_61_clk),
    .Q(\reg_file.reg_storage[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9260_ (.D(_0474_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9261_ (.D(_0475_),
    .CLK(clknet_leaf_65_clk),
    .Q(\reg_file.reg_storage[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9262_ (.D(_0476_),
    .CLK(clknet_leaf_49_clk),
    .Q(\reg_file.reg_storage[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9263_ (.D(_0477_),
    .CLK(clknet_leaf_36_clk),
    .Q(\reg_file.reg_storage[7][29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9264_ (.D(_0478_),
    .CLK(clknet_leaf_34_clk),
    .Q(\reg_file.reg_storage[7][30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9265_ (.D(_0479_),
    .CLK(clknet_leaf_42_clk),
    .Q(\reg_file.reg_storage[7][31] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(inst[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(inst[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(inst[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(inst[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input13 (.I(inst[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(inst[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(inst[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(inst[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input17 (.I(inst[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(inst[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(inst[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input2 (.I(inst[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(inst[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(inst[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(inst[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(inst[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input24 (.I(inst[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input25 (.I(inst[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input26 (.I(inst[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input27 (.I(inst[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input28 (.I(inst[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input29 (.I(inst[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input3 (.I(inst[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input30 (.I(inst[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input31 (.I(inst[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(inst[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input33 (.I(mem_load_out[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(mem_load_out[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input35 (.I(mem_load_out[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input36 (.I(mem_load_out[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input37 (.I(mem_load_out[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input38 (.I(mem_load_out[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input39 (.I(mem_load_out[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input4 (.I(inst[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input40 (.I(mem_load_out[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input41 (.I(mem_load_out[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input42 (.I(mem_load_out[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(mem_load_out[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input44 (.I(mem_load_out[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input45 (.I(mem_load_out[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(mem_load_out[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(mem_load_out[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input48 (.I(mem_load_out[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input49 (.I(mem_load_out[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input5 (.I(inst[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input50 (.I(mem_load_out[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input51 (.I(mem_load_out[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input52 (.I(mem_load_out[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input53 (.I(mem_load_out[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input54 (.I(mem_load_out[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input55 (.I(mem_load_out[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input56 (.I(mem_load_out[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input57 (.I(mem_load_out[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input58 (.I(mem_load_out[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input59 (.I(mem_load_out[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(inst[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input60 (.I(mem_load_out[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input61 (.I(mem_load_out[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(mem_load_out[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input63 (.I(mem_load_out[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input64 (.I(mem_load_out[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input65 (.I(pc[0]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input66 (.I(pc[10]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input67 (.I(pc[11]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(pc[12]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input69 (.I(pc[13]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input7 (.I(inst[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input70 (.I(pc[14]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input71 (.I(pc[15]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input72 (.I(pc[16]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input73 (.I(pc[17]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input74 (.I(pc[18]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input75 (.I(pc[19]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input76 (.I(pc[1]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input77 (.I(pc[20]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input78 (.I(pc[21]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input79 (.I(pc[22]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(inst[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input80 (.I(pc[23]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input81 (.I(pc[24]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input82 (.I(pc[25]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input83 (.I(pc[26]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input84 (.I(pc[27]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input85 (.I(pc[28]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input86 (.I(pc[29]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input87 (.I(pc[2]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input88 (.I(pc[30]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input89 (.I(pc[31]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(inst[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input90 (.I(pc[3]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input91 (.I(pc[4]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input92 (.I(pc[5]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input93 (.I(pc[6]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input94 (.I(pc[7]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input95 (.I(pc[8]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input96 (.I(pc[9]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap161 (.I(net121),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap162 (.I(_2222_),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap163 (.I(net118),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap164 (.I(_2181_),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap165 (.I(_1935_),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 max_cap166 (.I(_2799_),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output100 (.I(net100),
    .Z(alu_out_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output101 (.I(net101),
    .Z(alu_out_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output102 (.I(net102),
    .Z(alu_out_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output103 (.I(net103),
    .Z(alu_out_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output104 (.I(net104),
    .Z(alu_out_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output105 (.I(net105),
    .Z(alu_out_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output106 (.I(net106),
    .Z(alu_out_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output107 (.I(net107),
    .Z(alu_out_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output108 (.I(net108),
    .Z(alu_out_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output109 (.I(net109),
    .Z(alu_out_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output110 (.I(net110),
    .Z(alu_out_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output111 (.I(net111),
    .Z(alu_out_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output112 (.I(net112),
    .Z(alu_out_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output113 (.I(net113),
    .Z(alu_out_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output114 (.I(net114),
    .Z(alu_out_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output115 (.I(net115),
    .Z(alu_out_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output116 (.I(net116),
    .Z(alu_out_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output117 (.I(net117),
    .Z(alu_out_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output118 (.I(net163),
    .Z(alu_out_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output119 (.I(net119),
    .Z(alu_out_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output120 (.I(net120),
    .Z(alu_out_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output121 (.I(net161),
    .Z(alu_out_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output122 (.I(net122),
    .Z(alu_out_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output123 (.I(net123),
    .Z(alu_out_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output124 (.I(net124),
    .Z(alu_out_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output125 (.I(net125),
    .Z(alu_out_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output126 (.I(net126),
    .Z(alu_out_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output127 (.I(net127),
    .Z(alu_out_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output128 (.I(net128),
    .Z(alu_out_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output129 (.I(net129),
    .Z(pc_next[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output130 (.I(net130),
    .Z(pc_next[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output131 (.I(net131),
    .Z(pc_next[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output132 (.I(net132),
    .Z(pc_next[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output133 (.I(net133),
    .Z(pc_next[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output134 (.I(net134),
    .Z(pc_next[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output135 (.I(net135),
    .Z(pc_next[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output136 (.I(net136),
    .Z(pc_next[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output137 (.I(net137),
    .Z(pc_next[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output138 (.I(net138),
    .Z(pc_next[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output139 (.I(net139),
    .Z(pc_next[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output140 (.I(net140),
    .Z(pc_next[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output141 (.I(net141),
    .Z(pc_next[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output142 (.I(net142),
    .Z(pc_next[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output143 (.I(net143),
    .Z(pc_next[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output144 (.I(net144),
    .Z(pc_next[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output145 (.I(net145),
    .Z(pc_next[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output146 (.I(net146),
    .Z(pc_next[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output147 (.I(net147),
    .Z(pc_next[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output148 (.I(net148),
    .Z(pc_next[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output149 (.I(net149),
    .Z(pc_next[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output150 (.I(net150),
    .Z(pc_next[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output151 (.I(net151),
    .Z(pc_next[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output152 (.I(net152),
    .Z(pc_next[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output153 (.I(net153),
    .Z(pc_next[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output154 (.I(net154),
    .Z(pc_next[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output155 (.I(net155),
    .Z(pc_next[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output156 (.I(net156),
    .Z(pc_next[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output157 (.I(net157),
    .Z(pc_next[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output158 (.I(net158),
    .Z(pc_next[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output159 (.I(net159),
    .Z(pc_next[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output160 (.I(net160),
    .Z(pc_next[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output97 (.I(net97),
    .Z(alu_out_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output98 (.I(net98),
    .Z(alu_out_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output99 (.I(net99),
    .Z(alu_out_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer1 (.I(_2336_),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(net175),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_1529_),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(net177),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer13 (.I(_2281_),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer14 (.I(net181),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(_0963_),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer16 (.I(_1202_),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer17 (.I(_1196_),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer18 (.I(_0744_),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer19 (.I(_0762_),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(_1428_),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer20 (.I(_1483_),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer21 (.I(net201),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer22 (.I(_0963_),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer23 (.I(_2283_),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer24 (.I(net189),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer25 (.I(net228),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer26 (.I(_1097_),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer27 (.I(_2138_),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer28 (.I(net193),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer29 (.I(_2025_),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer3 (.I(_2428_),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer30 (.I(net195),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer31 (.I(_1049_),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer32 (.I(_1049_),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer33 (.I(_1178_),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer34 (.I(_1278_),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer35 (.I(net214),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer36 (.I(_2346_),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer37 (.I(_2190_),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer38 (.I(_1880_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer39 (.I(_1046_),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_1879_),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer40 (.I(net205),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer41 (.I(_0935_),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer42 (.I(_0967_),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer43 (.I(net208),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer44 (.I(_1628_),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer45 (.I(_1720_),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer46 (.I(_1434_),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer47 (.I(net229),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer48 (.I(_1110_),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer49 (.I(_2675_),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_1851_),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer50 (.I(_1213_),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer51 (.I(_1871_),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer52 (.I(net121),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer53 (.I(_1518_),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer54 (.I(net219),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer55 (.I(_1210_),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer56 (.I(_1643_),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer57 (.I(net222),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer58 (.I(_0537_),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer59 (.I(_2222_),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(net191),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer60 (.I(_0964_),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer61 (.I(net226),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer62 (.I(_1097_),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer63 (.I(_1674_),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(net226),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer8 (.I(_1388_),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(net174),
    .Z(net175));
endmodule

