magic
tech gf180mcuD
magscale 1 5
timestamp 1699637964
<< obsm1 >>
rect 672 1538 39392 18454
<< metal2 >>
rect 784 19600 840 20000
rect 2016 19600 2072 20000
rect 3248 19600 3304 20000
rect 4480 19600 4536 20000
rect 5712 19600 5768 20000
rect 6944 19600 7000 20000
rect 8176 19600 8232 20000
rect 9408 19600 9464 20000
rect 10640 19600 10696 20000
rect 11872 19600 11928 20000
rect 13104 19600 13160 20000
rect 14336 19600 14392 20000
rect 15568 19600 15624 20000
rect 16800 19600 16856 20000
rect 18032 19600 18088 20000
rect 19264 19600 19320 20000
rect 20496 19600 20552 20000
rect 21728 19600 21784 20000
rect 22960 19600 23016 20000
rect 24192 19600 24248 20000
rect 25424 19600 25480 20000
rect 26656 19600 26712 20000
rect 27888 19600 27944 20000
rect 29120 19600 29176 20000
rect 30352 19600 30408 20000
rect 31584 19600 31640 20000
rect 32816 19600 32872 20000
rect 34048 19600 34104 20000
rect 35280 19600 35336 20000
rect 36512 19600 36568 20000
rect 37744 19600 37800 20000
rect 38976 19600 39032 20000
rect 1792 0 1848 400
rect 3808 0 3864 400
rect 5824 0 5880 400
rect 7840 0 7896 400
rect 9856 0 9912 400
rect 11872 0 11928 400
rect 13888 0 13944 400
rect 15904 0 15960 400
rect 17920 0 17976 400
rect 19936 0 19992 400
rect 21952 0 22008 400
rect 23968 0 24024 400
rect 25984 0 26040 400
rect 28000 0 28056 400
rect 30016 0 30072 400
rect 32032 0 32088 400
rect 34048 0 34104 400
rect 36064 0 36120 400
rect 38080 0 38136 400
<< obsm2 >>
rect 870 19570 1986 19642
rect 2102 19570 3218 19642
rect 3334 19570 4450 19642
rect 4566 19570 5682 19642
rect 5798 19570 6914 19642
rect 7030 19570 8146 19642
rect 8262 19570 9378 19642
rect 9494 19570 10610 19642
rect 10726 19570 11842 19642
rect 11958 19570 13074 19642
rect 13190 19570 14306 19642
rect 14422 19570 15538 19642
rect 15654 19570 16770 19642
rect 16886 19570 18002 19642
rect 18118 19570 19234 19642
rect 19350 19570 20466 19642
rect 20582 19570 21698 19642
rect 21814 19570 22930 19642
rect 23046 19570 24162 19642
rect 24278 19570 25394 19642
rect 25510 19570 26626 19642
rect 26742 19570 27858 19642
rect 27974 19570 29090 19642
rect 29206 19570 30322 19642
rect 30438 19570 31554 19642
rect 31670 19570 32786 19642
rect 32902 19570 34018 19642
rect 34134 19570 35250 19642
rect 35366 19570 36482 19642
rect 36598 19570 37714 19642
rect 37830 19570 38946 19642
rect 39062 19570 39378 19642
rect 798 430 39378 19570
rect 798 350 1762 430
rect 1878 350 3778 430
rect 3894 350 5794 430
rect 5910 350 7810 430
rect 7926 350 9826 430
rect 9942 350 11842 430
rect 11958 350 13858 430
rect 13974 350 15874 430
rect 15990 350 17890 430
rect 18006 350 19906 430
rect 20022 350 21922 430
rect 22038 350 23938 430
rect 24054 350 25954 430
rect 26070 350 27970 430
rect 28086 350 29986 430
rect 30102 350 32002 430
rect 32118 350 34018 430
rect 34134 350 36034 430
rect 36150 350 38050 430
rect 38166 350 39378 430
<< metal3 >>
rect 0 19152 400 19208
rect 39600 19152 40000 19208
rect 0 17920 400 17976
rect 39600 17920 40000 17976
rect 0 16688 400 16744
rect 39600 16688 40000 16744
rect 0 15456 400 15512
rect 39600 15456 40000 15512
rect 0 14224 400 14280
rect 39600 14224 40000 14280
rect 0 12992 400 13048
rect 39600 12992 40000 13048
rect 0 11760 400 11816
rect 39600 11760 40000 11816
rect 0 10528 400 10584
rect 39600 10528 40000 10584
rect 0 9296 400 9352
rect 39600 9296 40000 9352
rect 0 8064 400 8120
rect 39600 8064 40000 8120
rect 0 6832 400 6888
rect 39600 6832 40000 6888
rect 0 5600 400 5656
rect 39600 5600 40000 5656
rect 0 4368 400 4424
rect 39600 4368 40000 4424
rect 0 3136 400 3192
rect 39600 3136 40000 3192
rect 0 1904 400 1960
rect 39600 1904 40000 1960
rect 0 672 400 728
rect 39600 672 40000 728
<< obsm3 >>
rect 430 19122 39570 19194
rect 400 18006 39600 19122
rect 430 17890 39570 18006
rect 400 16774 39600 17890
rect 430 16658 39570 16774
rect 400 15542 39600 16658
rect 430 15426 39570 15542
rect 400 14310 39600 15426
rect 430 14194 39570 14310
rect 400 13078 39600 14194
rect 430 12962 39570 13078
rect 400 11846 39600 12962
rect 430 11730 39570 11846
rect 400 10614 39600 11730
rect 430 10498 39570 10614
rect 400 9382 39600 10498
rect 430 9266 39570 9382
rect 400 8150 39600 9266
rect 430 8034 39570 8150
rect 400 6918 39600 8034
rect 430 6802 39570 6918
rect 400 5686 39600 6802
rect 430 5570 39570 5686
rect 400 4454 39600 5570
rect 430 4338 39570 4454
rect 400 3222 39600 4338
rect 430 3106 39570 3222
rect 400 1990 39600 3106
rect 430 1874 39570 1990
rect 400 758 39600 1874
rect 430 686 39570 758
<< metal4 >>
rect 5422 1538 5582 18454
rect 10252 1538 10412 18454
rect 15082 1538 15242 18454
rect 19912 1538 20072 18454
rect 24742 1538 24902 18454
rect 29572 1538 29732 18454
rect 34402 1538 34562 18454
rect 39232 1538 39392 18454
<< labels >>
rlabel metal2 s 36064 0 36120 400 6 clk
port 1 nsew signal input
rlabel metal3 s 0 19152 400 19208 6 dmem_addr[0]
port 2 nsew signal output
rlabel metal3 s 0 6832 400 6888 6 dmem_addr[10]
port 3 nsew signal output
rlabel metal3 s 0 5600 400 5656 6 dmem_addr[11]
port 4 nsew signal output
rlabel metal3 s 0 4368 400 4424 6 dmem_addr[12]
port 5 nsew signal output
rlabel metal3 s 0 3136 400 3192 6 dmem_addr[13]
port 6 nsew signal output
rlabel metal3 s 0 1904 400 1960 6 dmem_addr[14]
port 7 nsew signal output
rlabel metal3 s 0 672 400 728 6 dmem_addr[15]
port 8 nsew signal output
rlabel metal3 s 0 17920 400 17976 6 dmem_addr[1]
port 9 nsew signal output
rlabel metal3 s 0 16688 400 16744 6 dmem_addr[2]
port 10 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 dmem_addr[3]
port 11 nsew signal output
rlabel metal3 s 0 14224 400 14280 6 dmem_addr[4]
port 12 nsew signal output
rlabel metal3 s 0 12992 400 13048 6 dmem_addr[5]
port 13 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 dmem_addr[6]
port 14 nsew signal output
rlabel metal3 s 0 10528 400 10584 6 dmem_addr[7]
port 15 nsew signal output
rlabel metal3 s 0 9296 400 9352 6 dmem_addr[8]
port 16 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 dmem_addr[9]
port 17 nsew signal output
rlabel metal3 s 39600 672 40000 728 6 dmem_data_in[0]
port 18 nsew signal output
rlabel metal3 s 39600 12992 40000 13048 6 dmem_data_in[10]
port 19 nsew signal output
rlabel metal3 s 39600 14224 40000 14280 6 dmem_data_in[11]
port 20 nsew signal output
rlabel metal3 s 39600 15456 40000 15512 6 dmem_data_in[12]
port 21 nsew signal output
rlabel metal3 s 39600 16688 40000 16744 6 dmem_data_in[13]
port 22 nsew signal output
rlabel metal3 s 39600 17920 40000 17976 6 dmem_data_in[14]
port 23 nsew signal output
rlabel metal3 s 39600 19152 40000 19208 6 dmem_data_in[15]
port 24 nsew signal output
rlabel metal3 s 39600 1904 40000 1960 6 dmem_data_in[1]
port 25 nsew signal output
rlabel metal3 s 39600 3136 40000 3192 6 dmem_data_in[2]
port 26 nsew signal output
rlabel metal3 s 39600 4368 40000 4424 6 dmem_data_in[3]
port 27 nsew signal output
rlabel metal3 s 39600 5600 40000 5656 6 dmem_data_in[4]
port 28 nsew signal output
rlabel metal3 s 39600 6832 40000 6888 6 dmem_data_in[5]
port 29 nsew signal output
rlabel metal3 s 39600 8064 40000 8120 6 dmem_data_in[6]
port 30 nsew signal output
rlabel metal3 s 39600 9296 40000 9352 6 dmem_data_in[7]
port 31 nsew signal output
rlabel metal3 s 39600 10528 40000 10584 6 dmem_data_in[8]
port 32 nsew signal output
rlabel metal3 s 39600 11760 40000 11816 6 dmem_data_in[9]
port 33 nsew signal output
rlabel metal2 s 1792 0 1848 400 6 dmem_data_out[0]
port 34 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 dmem_data_out[10]
port 35 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 dmem_data_out[11]
port 36 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 dmem_data_out[12]
port 37 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 dmem_data_out[13]
port 38 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 dmem_data_out[14]
port 39 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 dmem_data_out[15]
port 40 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 dmem_data_out[1]
port 41 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 dmem_data_out[2]
port 42 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 dmem_data_out[3]
port 43 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 dmem_data_out[4]
port 44 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 dmem_data_out[5]
port 45 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 dmem_data_out[6]
port 46 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 dmem_data_out[7]
port 47 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 dmem_data_out[8]
port 48 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 dmem_data_out[9]
port 49 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 dmem_we
port 50 nsew signal output
rlabel metal2 s 19264 19600 19320 20000 6 instr[0]
port 51 nsew signal input
rlabel metal2 s 6944 19600 7000 20000 6 instr[10]
port 52 nsew signal input
rlabel metal2 s 5712 19600 5768 20000 6 instr[11]
port 53 nsew signal input
rlabel metal2 s 4480 19600 4536 20000 6 instr[12]
port 54 nsew signal input
rlabel metal2 s 3248 19600 3304 20000 6 instr[13]
port 55 nsew signal input
rlabel metal2 s 2016 19600 2072 20000 6 instr[14]
port 56 nsew signal input
rlabel metal2 s 784 19600 840 20000 6 instr[15]
port 57 nsew signal input
rlabel metal2 s 18032 19600 18088 20000 6 instr[1]
port 58 nsew signal input
rlabel metal2 s 16800 19600 16856 20000 6 instr[2]
port 59 nsew signal input
rlabel metal2 s 15568 19600 15624 20000 6 instr[3]
port 60 nsew signal input
rlabel metal2 s 14336 19600 14392 20000 6 instr[4]
port 61 nsew signal input
rlabel metal2 s 13104 19600 13160 20000 6 instr[5]
port 62 nsew signal input
rlabel metal2 s 11872 19600 11928 20000 6 instr[6]
port 63 nsew signal input
rlabel metal2 s 10640 19600 10696 20000 6 instr[7]
port 64 nsew signal input
rlabel metal2 s 9408 19600 9464 20000 6 instr[8]
port 65 nsew signal input
rlabel metal2 s 8176 19600 8232 20000 6 instr[9]
port 66 nsew signal input
rlabel metal2 s 38976 19600 39032 20000 6 pc[0]
port 67 nsew signal output
rlabel metal2 s 26656 19600 26712 20000 6 pc[10]
port 68 nsew signal output
rlabel metal2 s 25424 19600 25480 20000 6 pc[11]
port 69 nsew signal output
rlabel metal2 s 24192 19600 24248 20000 6 pc[12]
port 70 nsew signal output
rlabel metal2 s 22960 19600 23016 20000 6 pc[13]
port 71 nsew signal output
rlabel metal2 s 21728 19600 21784 20000 6 pc[14]
port 72 nsew signal output
rlabel metal2 s 20496 19600 20552 20000 6 pc[15]
port 73 nsew signal output
rlabel metal2 s 37744 19600 37800 20000 6 pc[1]
port 74 nsew signal output
rlabel metal2 s 36512 19600 36568 20000 6 pc[2]
port 75 nsew signal output
rlabel metal2 s 35280 19600 35336 20000 6 pc[3]
port 76 nsew signal output
rlabel metal2 s 34048 19600 34104 20000 6 pc[4]
port 77 nsew signal output
rlabel metal2 s 32816 19600 32872 20000 6 pc[5]
port 78 nsew signal output
rlabel metal2 s 31584 19600 31640 20000 6 pc[6]
port 79 nsew signal output
rlabel metal2 s 30352 19600 30408 20000 6 pc[7]
port 80 nsew signal output
rlabel metal2 s 29120 19600 29176 20000 6 pc[8]
port 81 nsew signal output
rlabel metal2 s 27888 19600 27944 20000 6 pc[9]
port 82 nsew signal output
rlabel metal2 s 38080 0 38136 400 6 rst_n
port 83 nsew signal input
rlabel metal4 s 5422 1538 5582 18454 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 15082 1538 15242 18454 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 24742 1538 24902 18454 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 34402 1538 34562 18454 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 10252 1538 10412 18454 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 19912 1538 20072 18454 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 29572 1538 29732 18454 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 39232 1538 39392 18454 6 vss
port 85 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2805766
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/risc16/runs/23_11_10_12_35/results/signoff/risc16.magic.gds
string GDS_START 410372
<< end >>

