VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tjrpu
  CLASS BLOCK ;
  FOREIGN tjrpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 800.000 ;
  PIN gpu_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2760.800 796.000 2761.360 800.000 ;
    END
  END gpu_clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 99.680 2800.000 100.240 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 692.160 4.000 692.720 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.800 4.000 689.360 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 685.440 4.000 686.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.720 4.000 679.280 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.360 4.000 675.920 ;
    END
  END io_in[15]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 103.040 2800.000 103.600 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 106.400 2800.000 106.960 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 109.760 2800.000 110.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 113.120 2800.000 113.680 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 116.480 2800.000 117.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 119.840 2800.000 120.400 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 123.200 2800.000 123.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 698.880 4.000 699.440 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 695.520 4.000 696.080 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 101.920 2800.000 102.480 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 689.920 4.000 690.480 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 686.560 4.000 687.120 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 683.200 4.000 683.760 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 679.840 4.000 680.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 676.480 4.000 677.040 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 673.120 4.000 673.680 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 105.280 2800.000 105.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 108.640 2800.000 109.200 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 112.000 2800.000 112.560 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 115.360 2800.000 115.920 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 118.720 2800.000 119.280 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 122.080 2800.000 122.640 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 125.440 2800.000 126.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 696.640 4.000 697.200 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 693.280 4.000 693.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 100.800 2800.000 101.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 691.040 4.000 691.600 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 687.680 4.000 688.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 684.320 4.000 684.880 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 680.960 4.000 681.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 677.600 4.000 678.160 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 674.240 4.000 674.800 ;
    END
  END io_out[15]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 104.160 2800.000 104.720 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 107.520 2800.000 108.080 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 110.880 2800.000 111.440 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 114.240 2800.000 114.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 117.600 2800.000 118.160 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 120.960 2800.000 121.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 124.320 2800.000 124.880 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 697.760 4.000 698.320 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1036.000 0.000 1036.560 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1039.360 0.000 1039.920 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1042.720 0.000 1043.280 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.680 0.000 492.240 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 0.000 502.320 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 0.000 512.400 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 0.000 522.480 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 0.000 542.640 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 0.000 552.720 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 0.000 562.800 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 572.320 0.000 572.880 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 0.000 582.960 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 0.000 593.040 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 612.640 0.000 613.200 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 0.000 623.280 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 0.000 633.360 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 642.880 0.000 643.440 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 652.960 0.000 653.520 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 663.040 0.000 663.600 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 0.000 673.680 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 0.000 683.760 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 0.000 411.600 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 0.000 693.840 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 703.360 0.000 703.920 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 713.440 0.000 714.000 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 0.000 724.080 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 733.600 0.000 734.160 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 0.000 744.240 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 753.760 0.000 754.320 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 773.920 0.000 774.480 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 784.000 0.000 784.560 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 0.000 421.680 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 0.000 794.640 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 804.160 0.000 804.720 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.240 0.000 814.800 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 0.000 824.880 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 834.400 0.000 834.960 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 844.480 0.000 845.040 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 854.560 0.000 855.120 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 864.640 0.000 865.200 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 874.720 0.000 875.280 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 0.000 885.360 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 0.000 431.760 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.880 0.000 895.440 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 904.960 0.000 905.520 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 915.040 0.000 915.600 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 925.120 0.000 925.680 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 935.200 0.000 935.760 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 945.280 0.000 945.840 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 955.360 0.000 955.920 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 965.440 0.000 966.000 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 975.520 0.000 976.080 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 985.600 0.000 986.160 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 995.680 0.000 996.240 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1005.760 0.000 1006.320 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1015.840 0.000 1016.400 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1025.920 0.000 1026.480 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 0.000 472.080 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 0.000 394.800 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 0.000 495.600 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 0.000 505.680 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 0.000 525.840 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 0.000 535.920 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 545.440 0.000 546.000 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 0.000 556.080 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 0.000 566.160 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 585.760 0.000 586.320 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 0.000 404.880 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 595.840 0.000 596.400 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 0.000 606.480 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 0.000 616.560 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 0.000 626.640 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 636.160 0.000 636.720 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 0.000 646.800 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 0.000 656.880 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 0.000 666.960 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 676.480 0.000 677.040 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 686.560 0.000 687.120 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 0.000 707.280 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 716.800 0.000 717.360 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 726.880 0.000 727.440 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 0.000 737.520 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 747.040 0.000 747.600 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 757.120 0.000 757.680 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 777.280 0.000 777.840 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 787.360 0.000 787.920 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 797.440 0.000 798.000 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 807.520 0.000 808.080 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 0.000 818.160 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 0.000 828.240 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 0.000 838.320 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 847.840 0.000 848.400 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 0.000 858.480 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 868.000 0.000 868.560 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 878.080 0.000 878.640 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 888.160 0.000 888.720 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 0.000 435.120 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 898.240 0.000 898.800 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 908.320 0.000 908.880 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 918.400 0.000 918.960 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 928.480 0.000 929.040 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 0.000 939.120 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 948.640 0.000 949.200 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 958.720 0.000 959.280 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 968.800 0.000 969.360 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 978.880 0.000 979.440 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 988.960 0.000 989.520 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 0.000 445.200 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 999.040 0.000 999.600 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1009.120 0.000 1009.680 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1019.200 0.000 1019.760 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1029.280 0.000 1029.840 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 0.000 455.280 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 0.000 465.360 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 0.000 475.440 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 0.000 485.520 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 0.000 398.160 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 0.000 498.960 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 0.000 519.120 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 0.000 529.200 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 0.000 539.280 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 0.000 559.440 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.960 0.000 569.520 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 0.000 589.680 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 0.000 408.240 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 0.000 599.760 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.280 0.000 609.840 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 0.000 619.920 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 0.000 630.000 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 0.000 640.080 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 0.000 660.240 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 0.000 670.320 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 679.840 0.000 680.400 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 0.000 690.480 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 0.000 418.320 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 700.000 0.000 700.560 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 0.000 710.640 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 0.000 720.720 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 730.240 0.000 730.800 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 0.000 740.880 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 750.400 0.000 750.960 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 0.000 761.040 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 770.560 0.000 771.120 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 780.640 0.000 781.200 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 0.000 791.280 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 0.000 428.400 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 0.000 801.360 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 810.880 0.000 811.440 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 0.000 821.520 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 831.040 0.000 831.600 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 0.000 841.680 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 851.200 0.000 851.760 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 871.360 0.000 871.920 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 0.000 882.000 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 891.520 0.000 892.080 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 0.000 438.480 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 0.000 902.160 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 911.680 0.000 912.240 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 921.760 0.000 922.320 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 931.840 0.000 932.400 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 941.920 0.000 942.480 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 0.000 952.560 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 0.000 962.640 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 972.160 0.000 972.720 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 982.240 0.000 982.800 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 992.320 0.000 992.880 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 0.000 448.560 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1002.400 0.000 1002.960 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1012.480 0.000 1013.040 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1022.560 0.000 1023.120 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1032.640 0.000 1033.200 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 0.000 468.720 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 0.000 478.800 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 0.000 488.880 4.000 ;
    END
  END la_oenb[9]
  PIN tri_wbs_ack_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1377.600 796.000 1378.160 800.000 ;
    END
  END tri_wbs_ack_o[0]
  PIN tri_wbs_ack_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1164.800 796.000 1165.360 800.000 ;
    END
  END tri_wbs_ack_o[10]
  PIN tri_wbs_ack_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1143.520 796.000 1144.080 800.000 ;
    END
  END tri_wbs_ack_o[11]
  PIN tri_wbs_ack_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1122.240 796.000 1122.800 800.000 ;
    END
  END tri_wbs_ack_o[12]
  PIN tri_wbs_ack_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1100.960 796.000 1101.520 800.000 ;
    END
  END tri_wbs_ack_o[13]
  PIN tri_wbs_ack_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1079.680 796.000 1080.240 800.000 ;
    END
  END tri_wbs_ack_o[14]
  PIN tri_wbs_ack_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 796.000 1058.960 800.000 ;
    END
  END tri_wbs_ack_o[15]
  PIN tri_wbs_ack_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1037.120 796.000 1037.680 800.000 ;
    END
  END tri_wbs_ack_o[16]
  PIN tri_wbs_ack_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1015.840 796.000 1016.400 800.000 ;
    END
  END tri_wbs_ack_o[17]
  PIN tri_wbs_ack_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 796.000 995.120 800.000 ;
    END
  END tri_wbs_ack_o[18]
  PIN tri_wbs_ack_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 796.000 973.840 800.000 ;
    END
  END tri_wbs_ack_o[19]
  PIN tri_wbs_ack_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1356.320 796.000 1356.880 800.000 ;
    END
  END tri_wbs_ack_o[1]
  PIN tri_wbs_ack_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 796.000 952.560 800.000 ;
    END
  END tri_wbs_ack_o[20]
  PIN tri_wbs_ack_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 796.000 931.280 800.000 ;
    END
  END tri_wbs_ack_o[21]
  PIN tri_wbs_ack_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 909.440 796.000 910.000 800.000 ;
    END
  END tri_wbs_ack_o[22]
  PIN tri_wbs_ack_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 888.160 796.000 888.720 800.000 ;
    END
  END tri_wbs_ack_o[23]
  PIN tri_wbs_ack_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 796.000 867.440 800.000 ;
    END
  END tri_wbs_ack_o[24]
  PIN tri_wbs_ack_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 845.600 796.000 846.160 800.000 ;
    END
  END tri_wbs_ack_o[25]
  PIN tri_wbs_ack_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 796.000 824.880 800.000 ;
    END
  END tri_wbs_ack_o[26]
  PIN tri_wbs_ack_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 796.000 803.600 800.000 ;
    END
  END tri_wbs_ack_o[27]
  PIN tri_wbs_ack_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 796.000 782.320 800.000 ;
    END
  END tri_wbs_ack_o[28]
  PIN tri_wbs_ack_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 796.000 761.040 800.000 ;
    END
  END tri_wbs_ack_o[29]
  PIN tri_wbs_ack_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1335.040 796.000 1335.600 800.000 ;
    END
  END tri_wbs_ack_o[2]
  PIN tri_wbs_ack_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 796.000 739.760 800.000 ;
    END
  END tri_wbs_ack_o[30]
  PIN tri_wbs_ack_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 717.920 796.000 718.480 800.000 ;
    END
  END tri_wbs_ack_o[31]
  PIN tri_wbs_ack_o[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 796.000 697.200 800.000 ;
    END
  END tri_wbs_ack_o[32]
  PIN tri_wbs_ack_o[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 796.000 675.920 800.000 ;
    END
  END tri_wbs_ack_o[33]
  PIN tri_wbs_ack_o[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 654.080 796.000 654.640 800.000 ;
    END
  END tri_wbs_ack_o[34]
  PIN tri_wbs_ack_o[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 796.000 633.360 800.000 ;
    END
  END tri_wbs_ack_o[35]
  PIN tri_wbs_ack_o[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 796.000 612.080 800.000 ;
    END
  END tri_wbs_ack_o[36]
  PIN tri_wbs_ack_o[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 796.000 590.800 800.000 ;
    END
  END tri_wbs_ack_o[37]
  PIN tri_wbs_ack_o[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 568.960 796.000 569.520 800.000 ;
    END
  END tri_wbs_ack_o[38]
  PIN tri_wbs_ack_o[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 796.000 548.240 800.000 ;
    END
  END tri_wbs_ack_o[39]
  PIN tri_wbs_ack_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1313.760 796.000 1314.320 800.000 ;
    END
  END tri_wbs_ack_o[3]
  PIN tri_wbs_ack_o[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 796.000 526.960 800.000 ;
    END
  END tri_wbs_ack_o[40]
  PIN tri_wbs_ack_o[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 796.000 505.680 800.000 ;
    END
  END tri_wbs_ack_o[41]
  PIN tri_wbs_ack_o[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 796.000 484.400 800.000 ;
    END
  END tri_wbs_ack_o[42]
  PIN tri_wbs_ack_o[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 796.000 463.120 800.000 ;
    END
  END tri_wbs_ack_o[43]
  PIN tri_wbs_ack_o[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 796.000 441.840 800.000 ;
    END
  END tri_wbs_ack_o[44]
  PIN tri_wbs_ack_o[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 796.000 420.560 800.000 ;
    END
  END tri_wbs_ack_o[45]
  PIN tri_wbs_ack_o[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 796.000 399.280 800.000 ;
    END
  END tri_wbs_ack_o[46]
  PIN tri_wbs_ack_o[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 796.000 378.000 800.000 ;
    END
  END tri_wbs_ack_o[47]
  PIN tri_wbs_ack_o[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 796.000 356.720 800.000 ;
    END
  END tri_wbs_ack_o[48]
  PIN tri_wbs_ack_o[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 796.000 335.440 800.000 ;
    END
  END tri_wbs_ack_o[49]
  PIN tri_wbs_ack_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1292.480 796.000 1293.040 800.000 ;
    END
  END tri_wbs_ack_o[4]
  PIN tri_wbs_ack_o[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 796.000 314.160 800.000 ;
    END
  END tri_wbs_ack_o[50]
  PIN tri_wbs_ack_o[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 796.000 292.880 800.000 ;
    END
  END tri_wbs_ack_o[51]
  PIN tri_wbs_ack_o[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 796.000 271.600 800.000 ;
    END
  END tri_wbs_ack_o[52]
  PIN tri_wbs_ack_o[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 796.000 250.320 800.000 ;
    END
  END tri_wbs_ack_o[53]
  PIN tri_wbs_ack_o[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 796.000 229.040 800.000 ;
    END
  END tri_wbs_ack_o[54]
  PIN tri_wbs_ack_o[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 796.000 207.760 800.000 ;
    END
  END tri_wbs_ack_o[55]
  PIN tri_wbs_ack_o[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 796.000 186.480 800.000 ;
    END
  END tri_wbs_ack_o[56]
  PIN tri_wbs_ack_o[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 796.000 165.200 800.000 ;
    END
  END tri_wbs_ack_o[57]
  PIN tri_wbs_ack_o[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 796.000 143.920 800.000 ;
    END
  END tri_wbs_ack_o[58]
  PIN tri_wbs_ack_o[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 796.000 122.640 800.000 ;
    END
  END tri_wbs_ack_o[59]
  PIN tri_wbs_ack_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1271.200 796.000 1271.760 800.000 ;
    END
  END tri_wbs_ack_o[5]
  PIN tri_wbs_ack_o[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 796.000 101.360 800.000 ;
    END
  END tri_wbs_ack_o[60]
  PIN tri_wbs_ack_o[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 796.000 80.080 800.000 ;
    END
  END tri_wbs_ack_o[61]
  PIN tri_wbs_ack_o[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 796.000 58.800 800.000 ;
    END
  END tri_wbs_ack_o[62]
  PIN tri_wbs_ack_o[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 796.000 37.520 800.000 ;
    END
  END tri_wbs_ack_o[63]
  PIN tri_wbs_ack_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1249.920 796.000 1250.480 800.000 ;
    END
  END tri_wbs_ack_o[6]
  PIN tri_wbs_ack_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1228.640 796.000 1229.200 800.000 ;
    END
  END tri_wbs_ack_o[7]
  PIN tri_wbs_ack_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1207.360 796.000 1207.920 800.000 ;
    END
  END tri_wbs_ack_o[8]
  PIN tri_wbs_ack_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1186.080 796.000 1186.640 800.000 ;
    END
  END tri_wbs_ack_o[9]
  PIN tri_wbs_stb_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2739.520 796.000 2740.080 800.000 ;
    END
  END tri_wbs_stb_i[0]
  PIN tri_wbs_stb_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2526.720 796.000 2527.280 800.000 ;
    END
  END tri_wbs_stb_i[10]
  PIN tri_wbs_stb_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2505.440 796.000 2506.000 800.000 ;
    END
  END tri_wbs_stb_i[11]
  PIN tri_wbs_stb_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2484.160 796.000 2484.720 800.000 ;
    END
  END tri_wbs_stb_i[12]
  PIN tri_wbs_stb_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2462.880 796.000 2463.440 800.000 ;
    END
  END tri_wbs_stb_i[13]
  PIN tri_wbs_stb_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2441.600 796.000 2442.160 800.000 ;
    END
  END tri_wbs_stb_i[14]
  PIN tri_wbs_stb_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2420.320 796.000 2420.880 800.000 ;
    END
  END tri_wbs_stb_i[15]
  PIN tri_wbs_stb_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2399.040 796.000 2399.600 800.000 ;
    END
  END tri_wbs_stb_i[16]
  PIN tri_wbs_stb_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2377.760 796.000 2378.320 800.000 ;
    END
  END tri_wbs_stb_i[17]
  PIN tri_wbs_stb_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2356.480 796.000 2357.040 800.000 ;
    END
  END tri_wbs_stb_i[18]
  PIN tri_wbs_stb_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2335.200 796.000 2335.760 800.000 ;
    END
  END tri_wbs_stb_i[19]
  PIN tri_wbs_stb_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2718.240 796.000 2718.800 800.000 ;
    END
  END tri_wbs_stb_i[1]
  PIN tri_wbs_stb_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2313.920 796.000 2314.480 800.000 ;
    END
  END tri_wbs_stb_i[20]
  PIN tri_wbs_stb_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2292.640 796.000 2293.200 800.000 ;
    END
  END tri_wbs_stb_i[21]
  PIN tri_wbs_stb_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2271.360 796.000 2271.920 800.000 ;
    END
  END tri_wbs_stb_i[22]
  PIN tri_wbs_stb_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2250.080 796.000 2250.640 800.000 ;
    END
  END tri_wbs_stb_i[23]
  PIN tri_wbs_stb_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2228.800 796.000 2229.360 800.000 ;
    END
  END tri_wbs_stb_i[24]
  PIN tri_wbs_stb_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2207.520 796.000 2208.080 800.000 ;
    END
  END tri_wbs_stb_i[25]
  PIN tri_wbs_stb_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2186.240 796.000 2186.800 800.000 ;
    END
  END tri_wbs_stb_i[26]
  PIN tri_wbs_stb_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2164.960 796.000 2165.520 800.000 ;
    END
  END tri_wbs_stb_i[27]
  PIN tri_wbs_stb_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2143.680 796.000 2144.240 800.000 ;
    END
  END tri_wbs_stb_i[28]
  PIN tri_wbs_stb_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2122.400 796.000 2122.960 800.000 ;
    END
  END tri_wbs_stb_i[29]
  PIN tri_wbs_stb_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2696.960 796.000 2697.520 800.000 ;
    END
  END tri_wbs_stb_i[2]
  PIN tri_wbs_stb_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2101.120 796.000 2101.680 800.000 ;
    END
  END tri_wbs_stb_i[30]
  PIN tri_wbs_stb_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2079.840 796.000 2080.400 800.000 ;
    END
  END tri_wbs_stb_i[31]
  PIN tri_wbs_stb_i[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2058.560 796.000 2059.120 800.000 ;
    END
  END tri_wbs_stb_i[32]
  PIN tri_wbs_stb_i[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2037.280 796.000 2037.840 800.000 ;
    END
  END tri_wbs_stb_i[33]
  PIN tri_wbs_stb_i[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2016.000 796.000 2016.560 800.000 ;
    END
  END tri_wbs_stb_i[34]
  PIN tri_wbs_stb_i[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1994.720 796.000 1995.280 800.000 ;
    END
  END tri_wbs_stb_i[35]
  PIN tri_wbs_stb_i[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1973.440 796.000 1974.000 800.000 ;
    END
  END tri_wbs_stb_i[36]
  PIN tri_wbs_stb_i[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1952.160 796.000 1952.720 800.000 ;
    END
  END tri_wbs_stb_i[37]
  PIN tri_wbs_stb_i[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1930.880 796.000 1931.440 800.000 ;
    END
  END tri_wbs_stb_i[38]
  PIN tri_wbs_stb_i[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1909.600 796.000 1910.160 800.000 ;
    END
  END tri_wbs_stb_i[39]
  PIN tri_wbs_stb_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2675.680 796.000 2676.240 800.000 ;
    END
  END tri_wbs_stb_i[3]
  PIN tri_wbs_stb_i[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1888.320 796.000 1888.880 800.000 ;
    END
  END tri_wbs_stb_i[40]
  PIN tri_wbs_stb_i[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1867.040 796.000 1867.600 800.000 ;
    END
  END tri_wbs_stb_i[41]
  PIN tri_wbs_stb_i[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1845.760 796.000 1846.320 800.000 ;
    END
  END tri_wbs_stb_i[42]
  PIN tri_wbs_stb_i[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1824.480 796.000 1825.040 800.000 ;
    END
  END tri_wbs_stb_i[43]
  PIN tri_wbs_stb_i[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1803.200 796.000 1803.760 800.000 ;
    END
  END tri_wbs_stb_i[44]
  PIN tri_wbs_stb_i[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1781.920 796.000 1782.480 800.000 ;
    END
  END tri_wbs_stb_i[45]
  PIN tri_wbs_stb_i[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1760.640 796.000 1761.200 800.000 ;
    END
  END tri_wbs_stb_i[46]
  PIN tri_wbs_stb_i[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1739.360 796.000 1739.920 800.000 ;
    END
  END tri_wbs_stb_i[47]
  PIN tri_wbs_stb_i[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1718.080 796.000 1718.640 800.000 ;
    END
  END tri_wbs_stb_i[48]
  PIN tri_wbs_stb_i[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1696.800 796.000 1697.360 800.000 ;
    END
  END tri_wbs_stb_i[49]
  PIN tri_wbs_stb_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2654.400 796.000 2654.960 800.000 ;
    END
  END tri_wbs_stb_i[4]
  PIN tri_wbs_stb_i[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1675.520 796.000 1676.080 800.000 ;
    END
  END tri_wbs_stb_i[50]
  PIN tri_wbs_stb_i[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1654.240 796.000 1654.800 800.000 ;
    END
  END tri_wbs_stb_i[51]
  PIN tri_wbs_stb_i[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1632.960 796.000 1633.520 800.000 ;
    END
  END tri_wbs_stb_i[52]
  PIN tri_wbs_stb_i[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1611.680 796.000 1612.240 800.000 ;
    END
  END tri_wbs_stb_i[53]
  PIN tri_wbs_stb_i[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1590.400 796.000 1590.960 800.000 ;
    END
  END tri_wbs_stb_i[54]
  PIN tri_wbs_stb_i[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1569.120 796.000 1569.680 800.000 ;
    END
  END tri_wbs_stb_i[55]
  PIN tri_wbs_stb_i[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1547.840 796.000 1548.400 800.000 ;
    END
  END tri_wbs_stb_i[56]
  PIN tri_wbs_stb_i[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1526.560 796.000 1527.120 800.000 ;
    END
  END tri_wbs_stb_i[57]
  PIN tri_wbs_stb_i[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1505.280 796.000 1505.840 800.000 ;
    END
  END tri_wbs_stb_i[58]
  PIN tri_wbs_stb_i[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1484.000 796.000 1484.560 800.000 ;
    END
  END tri_wbs_stb_i[59]
  PIN tri_wbs_stb_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2633.120 796.000 2633.680 800.000 ;
    END
  END tri_wbs_stb_i[5]
  PIN tri_wbs_stb_i[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1462.720 796.000 1463.280 800.000 ;
    END
  END tri_wbs_stb_i[60]
  PIN tri_wbs_stb_i[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1441.440 796.000 1442.000 800.000 ;
    END
  END tri_wbs_stb_i[61]
  PIN tri_wbs_stb_i[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1420.160 796.000 1420.720 800.000 ;
    END
  END tri_wbs_stb_i[62]
  PIN tri_wbs_stb_i[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1398.880 796.000 1399.440 800.000 ;
    END
  END tri_wbs_stb_i[63]
  PIN tri_wbs_stb_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2611.840 796.000 2612.400 800.000 ;
    END
  END tri_wbs_stb_i[6]
  PIN tri_wbs_stb_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2590.560 796.000 2591.120 800.000 ;
    END
  END tri_wbs_stb_i[7]
  PIN tri_wbs_stb_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2569.280 796.000 2569.840 800.000 ;
    END
  END tri_wbs_stb_i[8]
  PIN tri_wbs_stb_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2548.000 796.000 2548.560 800.000 ;
    END
  END tri_wbs_stb_i[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.120 0.000 169.680 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 0.000 220.080 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 0.000 300.720 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 0.000 310.800 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 0.000 330.960 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 0.000 351.120 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 0.000 371.280 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 0.000 129.360 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 0.000 223.440 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 0.000 233.520 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 0.000 243.600 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 0.000 263.760 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 0.000 283.920 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 303.520 0.000 304.080 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 0.000 344.400 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 0.000 354.480 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.160 0.000 384.720 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 0.000 196.560 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 0.000 206.640 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 0.000 216.720 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 0.000 236.880 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 0.000 267.120 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 0.000 75.600 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 0.000 277.200 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 0.000 317.520 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 0.000 327.600 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 0.000 337.680 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 88.480 0.000 89.040 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 0.000 378.000 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 0.000 102.480 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 0.000 166.320 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.555000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END wbs_we_i
  PIN x_end[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 672.000 4.000 672.560 ;
    END
  END x_end[0]
  PIN x_end[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END x_end[100]
  PIN x_end[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 4.000 559.440 ;
    END
  END x_end[101]
  PIN x_end[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.760 4.000 558.320 ;
    END
  END x_end[102]
  PIN x_end[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 556.640 4.000 557.200 ;
    END
  END x_end[103]
  PIN x_end[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 555.520 4.000 556.080 ;
    END
  END x_end[104]
  PIN x_end[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END x_end[105]
  PIN x_end[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 553.280 4.000 553.840 ;
    END
  END x_end[106]
  PIN x_end[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.160 4.000 552.720 ;
    END
  END x_end[107]
  PIN x_end[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 551.040 4.000 551.600 ;
    END
  END x_end[108]
  PIN x_end[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 549.920 4.000 550.480 ;
    END
  END x_end[109]
  PIN x_end[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 660.800 4.000 661.360 ;
    END
  END x_end[10]
  PIN x_end[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END x_end[110]
  PIN x_end[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END x_end[111]
  PIN x_end[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.560 4.000 547.120 ;
    END
  END x_end[112]
  PIN x_end[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 545.440 4.000 546.000 ;
    END
  END x_end[113]
  PIN x_end[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END x_end[114]
  PIN x_end[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.200 4.000 543.760 ;
    END
  END x_end[115]
  PIN x_end[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 542.080 4.000 542.640 ;
    END
  END x_end[116]
  PIN x_end[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.960 4.000 541.520 ;
    END
  END x_end[117]
  PIN x_end[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 539.840 4.000 540.400 ;
    END
  END x_end[118]
  PIN x_end[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 538.720 4.000 539.280 ;
    END
  END x_end[119]
  PIN x_end[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 659.680 4.000 660.240 ;
    END
  END x_end[11]
  PIN x_end[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END x_end[120]
  PIN x_end[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 536.480 4.000 537.040 ;
    END
  END x_end[121]
  PIN x_end[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 535.360 4.000 535.920 ;
    END
  END x_end[122]
  PIN x_end[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END x_end[123]
  PIN x_end[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 533.120 4.000 533.680 ;
    END
  END x_end[124]
  PIN x_end[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 532.000 4.000 532.560 ;
    END
  END x_end[125]
  PIN x_end[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 530.880 4.000 531.440 ;
    END
  END x_end[126]
  PIN x_end[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 529.760 4.000 530.320 ;
    END
  END x_end[127]
  PIN x_end[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.640 4.000 529.200 ;
    END
  END x_end[128]
  PIN x_end[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 527.520 4.000 528.080 ;
    END
  END x_end[129]
  PIN x_end[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 658.560 4.000 659.120 ;
    END
  END x_end[12]
  PIN x_end[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 526.400 4.000 526.960 ;
    END
  END x_end[130]
  PIN x_end[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 525.280 4.000 525.840 ;
    END
  END x_end[131]
  PIN x_end[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END x_end[132]
  PIN x_end[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 523.040 4.000 523.600 ;
    END
  END x_end[133]
  PIN x_end[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END x_end[134]
  PIN x_end[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END x_end[135]
  PIN x_end[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 519.680 4.000 520.240 ;
    END
  END x_end[136]
  PIN x_end[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 518.560 4.000 519.120 ;
    END
  END x_end[137]
  PIN x_end[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 517.440 4.000 518.000 ;
    END
  END x_end[138]
  PIN x_end[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 516.320 4.000 516.880 ;
    END
  END x_end[139]
  PIN x_end[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 657.440 4.000 658.000 ;
    END
  END x_end[13]
  PIN x_end[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.200 4.000 515.760 ;
    END
  END x_end[140]
  PIN x_end[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END x_end[141]
  PIN x_end[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 512.960 4.000 513.520 ;
    END
  END x_end[142]
  PIN x_end[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 511.840 4.000 512.400 ;
    END
  END x_end[143]
  PIN x_end[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.720 4.000 511.280 ;
    END
  END x_end[144]
  PIN x_end[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END x_end[145]
  PIN x_end[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 508.480 4.000 509.040 ;
    END
  END x_end[146]
  PIN x_end[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 507.360 4.000 507.920 ;
    END
  END x_end[147]
  PIN x_end[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 506.240 4.000 506.800 ;
    END
  END x_end[148]
  PIN x_end[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 505.120 4.000 505.680 ;
    END
  END x_end[149]
  PIN x_end[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 656.320 4.000 656.880 ;
    END
  END x_end[14]
  PIN x_end[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END x_end[150]
  PIN x_end[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 502.880 4.000 503.440 ;
    END
  END x_end[151]
  PIN x_end[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 501.760 4.000 502.320 ;
    END
  END x_end[152]
  PIN x_end[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 500.640 4.000 501.200 ;
    END
  END x_end[153]
  PIN x_end[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 499.520 4.000 500.080 ;
    END
  END x_end[154]
  PIN x_end[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 498.400 4.000 498.960 ;
    END
  END x_end[155]
  PIN x_end[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END x_end[156]
  PIN x_end[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 496.160 4.000 496.720 ;
    END
  END x_end[157]
  PIN x_end[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 495.040 4.000 495.600 ;
    END
  END x_end[158]
  PIN x_end[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 493.920 4.000 494.480 ;
    END
  END x_end[159]
  PIN x_end[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 655.200 4.000 655.760 ;
    END
  END x_end[15]
  PIN x_end[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 492.800 4.000 493.360 ;
    END
  END x_end[160]
  PIN x_end[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.680 4.000 492.240 ;
    END
  END x_end[161]
  PIN x_end[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.560 4.000 491.120 ;
    END
  END x_end[162]
  PIN x_end[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 489.440 4.000 490.000 ;
    END
  END x_end[163]
  PIN x_end[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END x_end[164]
  PIN x_end[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END x_end[165]
  PIN x_end[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 486.080 4.000 486.640 ;
    END
  END x_end[166]
  PIN x_end[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 484.960 4.000 485.520 ;
    END
  END x_end[167]
  PIN x_end[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.840 4.000 484.400 ;
    END
  END x_end[168]
  PIN x_end[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 482.720 4.000 483.280 ;
    END
  END x_end[169]
  PIN x_end[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 654.080 4.000 654.640 ;
    END
  END x_end[16]
  PIN x_end[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.600 4.000 482.160 ;
    END
  END x_end[170]
  PIN x_end[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END x_end[171]
  PIN x_end[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 479.360 4.000 479.920 ;
    END
  END x_end[172]
  PIN x_end[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.240 4.000 478.800 ;
    END
  END x_end[173]
  PIN x_end[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 477.120 4.000 477.680 ;
    END
  END x_end[174]
  PIN x_end[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END x_end[175]
  PIN x_end[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 474.880 4.000 475.440 ;
    END
  END x_end[176]
  PIN x_end[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.760 4.000 474.320 ;
    END
  END x_end[177]
  PIN x_end[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 472.640 4.000 473.200 ;
    END
  END x_end[178]
  PIN x_end[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 471.520 4.000 472.080 ;
    END
  END x_end[179]
  PIN x_end[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 652.960 4.000 653.520 ;
    END
  END x_end[17]
  PIN x_end[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END x_end[180]
  PIN x_end[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.280 4.000 469.840 ;
    END
  END x_end[181]
  PIN x_end[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 468.160 4.000 468.720 ;
    END
  END x_end[182]
  PIN x_end[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 467.040 4.000 467.600 ;
    END
  END x_end[183]
  PIN x_end[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 465.920 4.000 466.480 ;
    END
  END x_end[184]
  PIN x_end[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 464.800 4.000 465.360 ;
    END
  END x_end[185]
  PIN x_end[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.680 4.000 464.240 ;
    END
  END x_end[186]
  PIN x_end[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 462.560 4.000 463.120 ;
    END
  END x_end[187]
  PIN x_end[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 461.440 4.000 462.000 ;
    END
  END x_end[188]
  PIN x_end[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END x_end[189]
  PIN x_end[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.840 4.000 652.400 ;
    END
  END x_end[18]
  PIN x_end[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 459.200 4.000 459.760 ;
    END
  END x_end[190]
  PIN x_end[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 458.080 4.000 458.640 ;
    END
  END x_end[191]
  PIN x_end[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 456.960 4.000 457.520 ;
    END
  END x_end[192]
  PIN x_end[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 455.840 4.000 456.400 ;
    END
  END x_end[193]
  PIN x_end[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.720 4.000 455.280 ;
    END
  END x_end[194]
  PIN x_end[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END x_end[195]
  PIN x_end[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 452.480 4.000 453.040 ;
    END
  END x_end[196]
  PIN x_end[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 451.360 4.000 451.920 ;
    END
  END x_end[197]
  PIN x_end[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 450.240 4.000 450.800 ;
    END
  END x_end[198]
  PIN x_end[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 449.120 4.000 449.680 ;
    END
  END x_end[199]
  PIN x_end[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 650.720 4.000 651.280 ;
    END
  END x_end[19]
  PIN x_end[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 670.880 4.000 671.440 ;
    END
  END x_end[1]
  PIN x_end[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END x_end[200]
  PIN x_end[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 446.880 4.000 447.440 ;
    END
  END x_end[201]
  PIN x_end[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 445.760 4.000 446.320 ;
    END
  END x_end[202]
  PIN x_end[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 444.640 4.000 445.200 ;
    END
  END x_end[203]
  PIN x_end[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 443.520 4.000 444.080 ;
    END
  END x_end[204]
  PIN x_end[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END x_end[205]
  PIN x_end[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 441.280 4.000 441.840 ;
    END
  END x_end[206]
  PIN x_end[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 440.160 4.000 440.720 ;
    END
  END x_end[207]
  PIN x_end[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 439.040 4.000 439.600 ;
    END
  END x_end[208]
  PIN x_end[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 437.920 4.000 438.480 ;
    END
  END x_end[209]
  PIN x_end[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 649.600 4.000 650.160 ;
    END
  END x_end[20]
  PIN x_end[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.800 4.000 437.360 ;
    END
  END x_end[210]
  PIN x_end[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END x_end[211]
  PIN x_end[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 434.560 4.000 435.120 ;
    END
  END x_end[212]
  PIN x_end[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 433.440 4.000 434.000 ;
    END
  END x_end[213]
  PIN x_end[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 432.320 4.000 432.880 ;
    END
  END x_end[214]
  PIN x_end[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 431.200 4.000 431.760 ;
    END
  END x_end[215]
  PIN x_end[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 430.080 4.000 430.640 ;
    END
  END x_end[216]
  PIN x_end[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 428.960 4.000 429.520 ;
    END
  END x_end[217]
  PIN x_end[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 427.840 4.000 428.400 ;
    END
  END x_end[218]
  PIN x_end[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 426.720 4.000 427.280 ;
    END
  END x_end[219]
  PIN x_end[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 648.480 4.000 649.040 ;
    END
  END x_end[21]
  PIN x_end[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END x_end[220]
  PIN x_end[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 424.480 4.000 425.040 ;
    END
  END x_end[221]
  PIN x_end[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END x_end[222]
  PIN x_end[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 422.240 4.000 422.800 ;
    END
  END x_end[223]
  PIN x_end[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 421.120 4.000 421.680 ;
    END
  END x_end[224]
  PIN x_end[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 4.000 420.560 ;
    END
  END x_end[225]
  PIN x_end[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 418.880 4.000 419.440 ;
    END
  END x_end[226]
  PIN x_end[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.760 4.000 418.320 ;
    END
  END x_end[227]
  PIN x_end[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.640 4.000 417.200 ;
    END
  END x_end[228]
  PIN x_end[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 415.520 4.000 416.080 ;
    END
  END x_end[229]
  PIN x_end[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 647.360 4.000 647.920 ;
    END
  END x_end[22]
  PIN x_end[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END x_end[230]
  PIN x_end[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 413.280 4.000 413.840 ;
    END
  END x_end[231]
  PIN x_end[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 412.160 4.000 412.720 ;
    END
  END x_end[232]
  PIN x_end[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.040 4.000 411.600 ;
    END
  END x_end[233]
  PIN x_end[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 409.920 4.000 410.480 ;
    END
  END x_end[234]
  PIN x_end[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END x_end[235]
  PIN x_end[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 407.680 4.000 408.240 ;
    END
  END x_end[236]
  PIN x_end[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 406.560 4.000 407.120 ;
    END
  END x_end[237]
  PIN x_end[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 405.440 4.000 406.000 ;
    END
  END x_end[238]
  PIN x_end[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.320 4.000 404.880 ;
    END
  END x_end[239]
  PIN x_end[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 646.240 4.000 646.800 ;
    END
  END x_end[23]
  PIN x_end[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END x_end[240]
  PIN x_end[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 402.080 4.000 402.640 ;
    END
  END x_end[241]
  PIN x_end[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.960 4.000 401.520 ;
    END
  END x_end[242]
  PIN x_end[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 399.840 4.000 400.400 ;
    END
  END x_end[243]
  PIN x_end[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END x_end[244]
  PIN x_end[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.600 4.000 398.160 ;
    END
  END x_end[245]
  PIN x_end[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 396.480 4.000 397.040 ;
    END
  END x_end[246]
  PIN x_end[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 395.360 4.000 395.920 ;
    END
  END x_end[247]
  PIN x_end[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 394.240 4.000 394.800 ;
    END
  END x_end[248]
  PIN x_end[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.120 4.000 393.680 ;
    END
  END x_end[249]
  PIN x_end[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END x_end[24]
  PIN x_end[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.000 4.000 392.560 ;
    END
  END x_end[250]
  PIN x_end[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 390.880 4.000 391.440 ;
    END
  END x_end[251]
  PIN x_end[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.760 4.000 390.320 ;
    END
  END x_end[252]
  PIN x_end[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 388.640 4.000 389.200 ;
    END
  END x_end[253]
  PIN x_end[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 387.520 4.000 388.080 ;
    END
  END x_end[254]
  PIN x_end[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END x_end[255]
  PIN x_end[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 385.280 4.000 385.840 ;
    END
  END x_end[256]
  PIN x_end[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 384.160 4.000 384.720 ;
    END
  END x_end[257]
  PIN x_end[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 383.040 4.000 383.600 ;
    END
  END x_end[258]
  PIN x_end[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 381.920 4.000 382.480 ;
    END
  END x_end[259]
  PIN x_end[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 644.000 4.000 644.560 ;
    END
  END x_end[25]
  PIN x_end[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END x_end[260]
  PIN x_end[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.680 4.000 380.240 ;
    END
  END x_end[261]
  PIN x_end[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 378.560 4.000 379.120 ;
    END
  END x_end[262]
  PIN x_end[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.440 4.000 378.000 ;
    END
  END x_end[263]
  PIN x_end[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 376.320 4.000 376.880 ;
    END
  END x_end[264]
  PIN x_end[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 4.000 375.760 ;
    END
  END x_end[265]
  PIN x_end[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END x_end[266]
  PIN x_end[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.960 4.000 373.520 ;
    END
  END x_end[267]
  PIN x_end[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 371.840 4.000 372.400 ;
    END
  END x_end[268]
  PIN x_end[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 370.720 4.000 371.280 ;
    END
  END x_end[269]
  PIN x_end[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 642.880 4.000 643.440 ;
    END
  END x_end[26]
  PIN x_end[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.600 4.000 370.160 ;
    END
  END x_end[270]
  PIN x_end[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.480 4.000 369.040 ;
    END
  END x_end[271]
  PIN x_end[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 367.360 4.000 367.920 ;
    END
  END x_end[272]
  PIN x_end[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 366.240 4.000 366.800 ;
    END
  END x_end[273]
  PIN x_end[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.120 4.000 365.680 ;
    END
  END x_end[274]
  PIN x_end[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END x_end[275]
  PIN x_end[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.880 4.000 363.440 ;
    END
  END x_end[276]
  PIN x_end[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 361.760 4.000 362.320 ;
    END
  END x_end[277]
  PIN x_end[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 360.640 4.000 361.200 ;
    END
  END x_end[278]
  PIN x_end[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 359.520 4.000 360.080 ;
    END
  END x_end[279]
  PIN x_end[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 641.760 4.000 642.320 ;
    END
  END x_end[27]
  PIN x_end[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END x_end[280]
  PIN x_end[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 357.280 4.000 357.840 ;
    END
  END x_end[281]
  PIN x_end[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 356.160 4.000 356.720 ;
    END
  END x_end[282]
  PIN x_end[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.040 4.000 355.600 ;
    END
  END x_end[283]
  PIN x_end[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.920 4.000 354.480 ;
    END
  END x_end[284]
  PIN x_end[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END x_end[285]
  PIN x_end[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 351.680 4.000 352.240 ;
    END
  END x_end[286]
  PIN x_end[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 350.560 4.000 351.120 ;
    END
  END x_end[287]
  PIN x_end[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.440 4.000 350.000 ;
    END
  END x_end[288]
  PIN x_end[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 348.320 4.000 348.880 ;
    END
  END x_end[289]
  PIN x_end[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 640.640 4.000 641.200 ;
    END
  END x_end[28]
  PIN x_end[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END x_end[290]
  PIN x_end[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.080 4.000 346.640 ;
    END
  END x_end[291]
  PIN x_end[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.960 4.000 345.520 ;
    END
  END x_end[292]
  PIN x_end[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 343.840 4.000 344.400 ;
    END
  END x_end[293]
  PIN x_end[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.720 4.000 343.280 ;
    END
  END x_end[294]
  PIN x_end[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END x_end[295]
  PIN x_end[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 340.480 4.000 341.040 ;
    END
  END x_end[296]
  PIN x_end[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.360 4.000 339.920 ;
    END
  END x_end[297]
  PIN x_end[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 338.240 4.000 338.800 ;
    END
  END x_end[298]
  PIN x_end[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.120 4.000 337.680 ;
    END
  END x_end[299]
  PIN x_end[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 639.520 4.000 640.080 ;
    END
  END x_end[29]
  PIN x_end[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 669.760 4.000 670.320 ;
    END
  END x_end[2]
  PIN x_end[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END x_end[300]
  PIN x_end[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.880 4.000 335.440 ;
    END
  END x_end[301]
  PIN x_end[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 333.760 4.000 334.320 ;
    END
  END x_end[302]
  PIN x_end[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.640 4.000 333.200 ;
    END
  END x_end[303]
  PIN x_end[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 331.520 4.000 332.080 ;
    END
  END x_end[304]
  PIN x_end[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.400 4.000 330.960 ;
    END
  END x_end[305]
  PIN x_end[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 329.280 4.000 329.840 ;
    END
  END x_end[306]
  PIN x_end[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.160 4.000 328.720 ;
    END
  END x_end[307]
  PIN x_end[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 327.040 4.000 327.600 ;
    END
  END x_end[308]
  PIN x_end[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.920 4.000 326.480 ;
    END
  END x_end[309]
  PIN x_end[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.400 4.000 638.960 ;
    END
  END x_end[30]
  PIN x_end[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END x_end[310]
  PIN x_end[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 323.680 4.000 324.240 ;
    END
  END x_end[311]
  PIN x_end[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.560 4.000 323.120 ;
    END
  END x_end[312]
  PIN x_end[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 321.440 4.000 322.000 ;
    END
  END x_end[313]
  PIN x_end[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.320 4.000 320.880 ;
    END
  END x_end[314]
  PIN x_end[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END x_end[315]
  PIN x_end[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.080 4.000 318.640 ;
    END
  END x_end[316]
  PIN x_end[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.960 4.000 317.520 ;
    END
  END x_end[317]
  PIN x_end[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.840 4.000 316.400 ;
    END
  END x_end[318]
  PIN x_end[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 314.720 4.000 315.280 ;
    END
  END x_end[319]
  PIN x_end[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 637.280 4.000 637.840 ;
    END
  END x_end[31]
  PIN x_end[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END x_end[320]
  PIN x_end[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END x_end[321]
  PIN x_end[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.360 4.000 311.920 ;
    END
  END x_end[322]
  PIN x_end[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.240 4.000 310.800 ;
    END
  END x_end[323]
  PIN x_end[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END x_end[324]
  PIN x_end[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.000 4.000 308.560 ;
    END
  END x_end[325]
  PIN x_end[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.880 4.000 307.440 ;
    END
  END x_end[326]
  PIN x_end[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 305.760 4.000 306.320 ;
    END
  END x_end[327]
  PIN x_end[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 304.640 4.000 305.200 ;
    END
  END x_end[328]
  PIN x_end[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 303.520 4.000 304.080 ;
    END
  END x_end[329]
  PIN x_end[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 636.160 4.000 636.720 ;
    END
  END x_end[32]
  PIN x_end[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END x_end[330]
  PIN x_end[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.280 4.000 301.840 ;
    END
  END x_end[331]
  PIN x_end[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 300.160 4.000 300.720 ;
    END
  END x_end[332]
  PIN x_end[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.040 4.000 299.600 ;
    END
  END x_end[333]
  PIN x_end[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 297.920 4.000 298.480 ;
    END
  END x_end[334]
  PIN x_end[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.800 4.000 297.360 ;
    END
  END x_end[335]
  PIN x_end[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.680 4.000 296.240 ;
    END
  END x_end[336]
  PIN x_end[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.560 4.000 295.120 ;
    END
  END x_end[337]
  PIN x_end[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 293.440 4.000 294.000 ;
    END
  END x_end[338]
  PIN x_end[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.320 4.000 292.880 ;
    END
  END x_end[339]
  PIN x_end[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END x_end[33]
  PIN x_end[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END x_end[340]
  PIN x_end[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.080 4.000 290.640 ;
    END
  END x_end[341]
  PIN x_end[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.960 4.000 289.520 ;
    END
  END x_end[342]
  PIN x_end[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END x_end[343]
  PIN x_end[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END x_end[344]
  PIN x_end[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END x_end[345]
  PIN x_end[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 284.480 4.000 285.040 ;
    END
  END x_end[346]
  PIN x_end[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.360 4.000 283.920 ;
    END
  END x_end[347]
  PIN x_end[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 282.240 4.000 282.800 ;
    END
  END x_end[348]
  PIN x_end[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.120 4.000 281.680 ;
    END
  END x_end[349]
  PIN x_end[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 633.920 4.000 634.480 ;
    END
  END x_end[34]
  PIN x_end[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END x_end[350]
  PIN x_end[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END x_end[351]
  PIN x_end[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 277.760 4.000 278.320 ;
    END
  END x_end[352]
  PIN x_end[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.640 4.000 277.200 ;
    END
  END x_end[353]
  PIN x_end[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END x_end[354]
  PIN x_end[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END x_end[355]
  PIN x_end[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.280 4.000 273.840 ;
    END
  END x_end[356]
  PIN x_end[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END x_end[357]
  PIN x_end[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.040 4.000 271.600 ;
    END
  END x_end[358]
  PIN x_end[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 4.000 270.480 ;
    END
  END x_end[359]
  PIN x_end[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END x_end[35]
  PIN x_end[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END x_end[360]
  PIN x_end[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.680 4.000 268.240 ;
    END
  END x_end[361]
  PIN x_end[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END x_end[362]
  PIN x_end[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 4.000 266.000 ;
    END
  END x_end[363]
  PIN x_end[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.320 4.000 264.880 ;
    END
  END x_end[364]
  PIN x_end[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END x_end[365]
  PIN x_end[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.080 4.000 262.640 ;
    END
  END x_end[366]
  PIN x_end[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END x_end[367]
  PIN x_end[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 259.840 4.000 260.400 ;
    END
  END x_end[368]
  PIN x_end[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 4.000 259.280 ;
    END
  END x_end[369]
  PIN x_end[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END x_end[36]
  PIN x_end[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END x_end[370]
  PIN x_end[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 4.000 257.040 ;
    END
  END x_end[371]
  PIN x_end[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END x_end[372]
  PIN x_end[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.240 4.000 254.800 ;
    END
  END x_end[373]
  PIN x_end[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 4.000 253.680 ;
    END
  END x_end[374]
  PIN x_end[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END x_end[375]
  PIN x_end[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.880 4.000 251.440 ;
    END
  END x_end[376]
  PIN x_end[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.760 4.000 250.320 ;
    END
  END x_end[377]
  PIN x_end[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.640 4.000 249.200 ;
    END
  END x_end[378]
  PIN x_end[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 247.520 4.000 248.080 ;
    END
  END x_end[379]
  PIN x_end[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 630.560 4.000 631.120 ;
    END
  END x_end[37]
  PIN x_end[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END x_end[380]
  PIN x_end[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 4.000 245.840 ;
    END
  END x_end[381]
  PIN x_end[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.160 4.000 244.720 ;
    END
  END x_end[382]
  PIN x_end[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.040 4.000 243.600 ;
    END
  END x_end[383]
  PIN x_end[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END x_end[384]
  PIN x_end[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END x_end[385]
  PIN x_end[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 239.680 4.000 240.240 ;
    END
  END x_end[386]
  PIN x_end[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END x_end[387]
  PIN x_end[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.440 4.000 238.000 ;
    END
  END x_end[388]
  PIN x_end[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 236.320 4.000 236.880 ;
    END
  END x_end[389]
  PIN x_end[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 629.440 4.000 630.000 ;
    END
  END x_end[38]
  PIN x_end[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 4.000 235.760 ;
    END
  END x_end[390]
  PIN x_end[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 4.000 234.640 ;
    END
  END x_end[391]
  PIN x_end[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END x_end[392]
  PIN x_end[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.840 4.000 232.400 ;
    END
  END x_end[393]
  PIN x_end[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.720 4.000 231.280 ;
    END
  END x_end[394]
  PIN x_end[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END x_end[395]
  PIN x_end[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.480 4.000 229.040 ;
    END
  END x_end[396]
  PIN x_end[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.360 4.000 227.920 ;
    END
  END x_end[397]
  PIN x_end[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 4.000 226.800 ;
    END
  END x_end[398]
  PIN x_end[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END x_end[399]
  PIN x_end[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 628.320 4.000 628.880 ;
    END
  END x_end[39]
  PIN x_end[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 668.640 4.000 669.200 ;
    END
  END x_end[3]
  PIN x_end[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END x_end[400]
  PIN x_end[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.880 4.000 223.440 ;
    END
  END x_end[401]
  PIN x_end[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END x_end[402]
  PIN x_end[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.640 4.000 221.200 ;
    END
  END x_end[403]
  PIN x_end[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.520 4.000 220.080 ;
    END
  END x_end[404]
  PIN x_end[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END x_end[405]
  PIN x_end[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.280 4.000 217.840 ;
    END
  END x_end[406]
  PIN x_end[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 4.000 216.720 ;
    END
  END x_end[407]
  PIN x_end[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 215.040 4.000 215.600 ;
    END
  END x_end[408]
  PIN x_end[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 4.000 214.480 ;
    END
  END x_end[409]
  PIN x_end[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 627.200 4.000 627.760 ;
    END
  END x_end[40]
  PIN x_end[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END x_end[410]
  PIN x_end[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END x_end[411]
  PIN x_end[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.560 4.000 211.120 ;
    END
  END x_end[412]
  PIN x_end[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 209.440 4.000 210.000 ;
    END
  END x_end[413]
  PIN x_end[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END x_end[414]
  PIN x_end[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END x_end[415]
  PIN x_end[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.080 4.000 206.640 ;
    END
  END x_end[416]
  PIN x_end[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END x_end[417]
  PIN x_end[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 203.840 4.000 204.400 ;
    END
  END x_end[418]
  PIN x_end[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.720 4.000 203.280 ;
    END
  END x_end[419]
  PIN x_end[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.080 4.000 626.640 ;
    END
  END x_end[41]
  PIN x_end[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END x_end[420]
  PIN x_end[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.480 4.000 201.040 ;
    END
  END x_end[421]
  PIN x_end[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END x_end[422]
  PIN x_end[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END x_end[423]
  PIN x_end[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.120 4.000 197.680 ;
    END
  END x_end[424]
  PIN x_end[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END x_end[425]
  PIN x_end[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END x_end[426]
  PIN x_end[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.760 4.000 194.320 ;
    END
  END x_end[427]
  PIN x_end[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 192.640 4.000 193.200 ;
    END
  END x_end[428]
  PIN x_end[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END x_end[429]
  PIN x_end[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END x_end[42]
  PIN x_end[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END x_end[430]
  PIN x_end[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END x_end[431]
  PIN x_end[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END x_end[432]
  PIN x_end[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 4.000 187.600 ;
    END
  END x_end[433]
  PIN x_end[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END x_end[434]
  PIN x_end[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END x_end[435]
  PIN x_end[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.680 4.000 184.240 ;
    END
  END x_end[436]
  PIN x_end[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 4.000 183.120 ;
    END
  END x_end[437]
  PIN x_end[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END x_end[438]
  PIN x_end[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END x_end[439]
  PIN x_end[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 623.840 4.000 624.400 ;
    END
  END x_end[43]
  PIN x_end[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END x_end[440]
  PIN x_end[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END x_end[441]
  PIN x_end[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END x_end[442]
  PIN x_end[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 175.840 4.000 176.400 ;
    END
  END x_end[443]
  PIN x_end[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END x_end[444]
  PIN x_end[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 4.000 174.160 ;
    END
  END x_end[445]
  PIN x_end[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.480 4.000 173.040 ;
    END
  END x_end[446]
  PIN x_end[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END x_end[447]
  PIN x_end[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.240 4.000 170.800 ;
    END
  END x_end[448]
  PIN x_end[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 4.000 169.680 ;
    END
  END x_end[449]
  PIN x_end[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 622.720 4.000 623.280 ;
    END
  END x_end[44]
  PIN x_end[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END x_end[450]
  PIN x_end[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END x_end[451]
  PIN x_end[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END x_end[452]
  PIN x_end[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END x_end[453]
  PIN x_end[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.520 4.000 164.080 ;
    END
  END x_end[454]
  PIN x_end[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 4.000 162.960 ;
    END
  END x_end[455]
  PIN x_end[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END x_end[456]
  PIN x_end[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 4.000 160.720 ;
    END
  END x_end[457]
  PIN x_end[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 4.000 159.600 ;
    END
  END x_end[458]
  PIN x_end[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END x_end[459]
  PIN x_end[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.600 4.000 622.160 ;
    END
  END x_end[45]
  PIN x_end[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END x_end[460]
  PIN x_end[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 4.000 156.240 ;
    END
  END x_end[461]
  PIN x_end[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END x_end[462]
  PIN x_end[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.440 4.000 154.000 ;
    END
  END x_end[463]
  PIN x_end[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END x_end[464]
  PIN x_end[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END x_end[465]
  PIN x_end[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.080 4.000 150.640 ;
    END
  END x_end[466]
  PIN x_end[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 4.000 149.520 ;
    END
  END x_end[467]
  PIN x_end[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END x_end[468]
  PIN x_end[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 4.000 147.280 ;
    END
  END x_end[469]
  PIN x_end[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 620.480 4.000 621.040 ;
    END
  END x_end[46]
  PIN x_end[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END x_end[470]
  PIN x_end[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END x_end[471]
  PIN x_end[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.360 4.000 143.920 ;
    END
  END x_end[472]
  PIN x_end[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 4.000 142.800 ;
    END
  END x_end[473]
  PIN x_end[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END x_end[474]
  PIN x_end[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END x_end[475]
  PIN x_end[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 138.880 4.000 139.440 ;
    END
  END x_end[476]
  PIN x_end[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END x_end[477]
  PIN x_end[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.640 4.000 137.200 ;
    END
  END x_end[478]
  PIN x_end[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 4.000 136.080 ;
    END
  END x_end[479]
  PIN x_end[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 619.360 4.000 619.920 ;
    END
  END x_end[47]
  PIN x_end[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END x_end[480]
  PIN x_end[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 4.000 133.840 ;
    END
  END x_end[481]
  PIN x_end[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END x_end[482]
  PIN x_end[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END x_end[483]
  PIN x_end[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END x_end[484]
  PIN x_end[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 4.000 129.360 ;
    END
  END x_end[485]
  PIN x_end[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END x_end[486]
  PIN x_end[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 4.000 127.120 ;
    END
  END x_end[487]
  PIN x_end[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 125.440 4.000 126.000 ;
    END
  END x_end[488]
  PIN x_end[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END x_end[489]
  PIN x_end[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 618.240 4.000 618.800 ;
    END
  END x_end[48]
  PIN x_end[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END x_end[490]
  PIN x_end[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 4.000 122.640 ;
    END
  END x_end[491]
  PIN x_end[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END x_end[492]
  PIN x_end[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.840 4.000 120.400 ;
    END
  END x_end[493]
  PIN x_end[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END x_end[494]
  PIN x_end[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END x_end[495]
  PIN x_end[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.480 4.000 117.040 ;
    END
  END x_end[496]
  PIN x_end[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END x_end[497]
  PIN x_end[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END x_end[498]
  PIN x_end[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 4.000 113.680 ;
    END
  END x_end[499]
  PIN x_end[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 617.120 4.000 617.680 ;
    END
  END x_end[49]
  PIN x_end[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 667.520 4.000 668.080 ;
    END
  END x_end[4]
  PIN x_end[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END x_end[500]
  PIN x_end[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END x_end[501]
  PIN x_end[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.760 4.000 110.320 ;
    END
  END x_end[502]
  PIN x_end[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 108.640 4.000 109.200 ;
    END
  END x_end[503]
  PIN x_end[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END x_end[504]
  PIN x_end[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END x_end[505]
  PIN x_end[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END x_end[506]
  PIN x_end[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END x_end[507]
  PIN x_end[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.040 4.000 103.600 ;
    END
  END x_end[508]
  PIN x_end[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 4.000 102.480 ;
    END
  END x_end[509]
  PIN x_end[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 616.000 4.000 616.560 ;
    END
  END x_end[50]
  PIN x_end[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END x_end[510]
  PIN x_end[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END x_end[511]
  PIN x_end[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END x_end[51]
  PIN x_end[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 613.760 4.000 614.320 ;
    END
  END x_end[52]
  PIN x_end[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 612.640 4.000 613.200 ;
    END
  END x_end[53]
  PIN x_end[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END x_end[54]
  PIN x_end[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 610.400 4.000 610.960 ;
    END
  END x_end[55]
  PIN x_end[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 609.280 4.000 609.840 ;
    END
  END x_end[56]
  PIN x_end[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END x_end[57]
  PIN x_end[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 607.040 4.000 607.600 ;
    END
  END x_end[58]
  PIN x_end[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 605.920 4.000 606.480 ;
    END
  END x_end[59]
  PIN x_end[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 666.400 4.000 666.960 ;
    END
  END x_end[5]
  PIN x_end[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END x_end[60]
  PIN x_end[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 603.680 4.000 604.240 ;
    END
  END x_end[61]
  PIN x_end[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.560 4.000 603.120 ;
    END
  END x_end[62]
  PIN x_end[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 601.440 4.000 602.000 ;
    END
  END x_end[63]
  PIN x_end[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 600.320 4.000 600.880 ;
    END
  END x_end[64]
  PIN x_end[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 599.200 4.000 599.760 ;
    END
  END x_end[65]
  PIN x_end[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 598.080 4.000 598.640 ;
    END
  END x_end[66]
  PIN x_end[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 596.960 4.000 597.520 ;
    END
  END x_end[67]
  PIN x_end[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END x_end[68]
  PIN x_end[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 4.000 595.280 ;
    END
  END x_end[69]
  PIN x_end[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END x_end[6]
  PIN x_end[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 593.600 4.000 594.160 ;
    END
  END x_end[70]
  PIN x_end[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 592.480 4.000 593.040 ;
    END
  END x_end[71]
  PIN x_end[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 591.360 4.000 591.920 ;
    END
  END x_end[72]
  PIN x_end[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 590.240 4.000 590.800 ;
    END
  END x_end[73]
  PIN x_end[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.120 4.000 589.680 ;
    END
  END x_end[74]
  PIN x_end[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 588.000 4.000 588.560 ;
    END
  END x_end[75]
  PIN x_end[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 586.880 4.000 587.440 ;
    END
  END x_end[76]
  PIN x_end[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 585.760 4.000 586.320 ;
    END
  END x_end[77]
  PIN x_end[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 584.640 4.000 585.200 ;
    END
  END x_end[78]
  PIN x_end[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 583.520 4.000 584.080 ;
    END
  END x_end[79]
  PIN x_end[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 664.160 4.000 664.720 ;
    END
  END x_end[7]
  PIN x_end[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 582.400 4.000 582.960 ;
    END
  END x_end[80]
  PIN x_end[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 4.000 581.840 ;
    END
  END x_end[81]
  PIN x_end[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 580.160 4.000 580.720 ;
    END
  END x_end[82]
  PIN x_end[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 579.040 4.000 579.600 ;
    END
  END x_end[83]
  PIN x_end[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END x_end[84]
  PIN x_end[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 576.800 4.000 577.360 ;
    END
  END x_end[85]
  PIN x_end[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 575.680 4.000 576.240 ;
    END
  END x_end[86]
  PIN x_end[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END x_end[87]
  PIN x_end[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 573.440 4.000 574.000 ;
    END
  END x_end[88]
  PIN x_end[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 572.320 4.000 572.880 ;
    END
  END x_end[89]
  PIN x_end[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.040 4.000 663.600 ;
    END
  END x_end[8]
  PIN x_end[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END x_end[90]
  PIN x_end[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 570.080 4.000 570.640 ;
    END
  END x_end[91]
  PIN x_end[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 568.960 4.000 569.520 ;
    END
  END x_end[92]
  PIN x_end[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 4.000 568.400 ;
    END
  END x_end[93]
  PIN x_end[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 566.720 4.000 567.280 ;
    END
  END x_end[94]
  PIN x_end[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.600 4.000 566.160 ;
    END
  END x_end[95]
  PIN x_end[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 564.480 4.000 565.040 ;
    END
  END x_end[96]
  PIN x_end[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 563.360 4.000 563.920 ;
    END
  END x_end[97]
  PIN x_end[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 562.240 4.000 562.800 ;
    END
  END x_end[98]
  PIN x_end[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END x_end[99]
  PIN x_end[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 661.920 4.000 662.480 ;
    END
  END x_end[9]
  PIN x_start[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 126.560 2800.000 127.120 ;
    END
  END x_start[0]
  PIN x_start[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 238.560 2800.000 239.120 ;
    END
  END x_start[100]
  PIN x_start[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 239.680 2800.000 240.240 ;
    END
  END x_start[101]
  PIN x_start[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 240.800 2800.000 241.360 ;
    END
  END x_start[102]
  PIN x_start[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 241.920 2800.000 242.480 ;
    END
  END x_start[103]
  PIN x_start[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 243.040 2800.000 243.600 ;
    END
  END x_start[104]
  PIN x_start[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 244.160 2800.000 244.720 ;
    END
  END x_start[105]
  PIN x_start[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 245.280 2800.000 245.840 ;
    END
  END x_start[106]
  PIN x_start[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 246.400 2800.000 246.960 ;
    END
  END x_start[107]
  PIN x_start[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 247.520 2800.000 248.080 ;
    END
  END x_start[108]
  PIN x_start[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 248.640 2800.000 249.200 ;
    END
  END x_start[109]
  PIN x_start[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 137.760 2800.000 138.320 ;
    END
  END x_start[10]
  PIN x_start[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 249.760 2800.000 250.320 ;
    END
  END x_start[110]
  PIN x_start[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 250.880 2800.000 251.440 ;
    END
  END x_start[111]
  PIN x_start[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 252.000 2800.000 252.560 ;
    END
  END x_start[112]
  PIN x_start[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 253.120 2800.000 253.680 ;
    END
  END x_start[113]
  PIN x_start[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 254.240 2800.000 254.800 ;
    END
  END x_start[114]
  PIN x_start[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 255.360 2800.000 255.920 ;
    END
  END x_start[115]
  PIN x_start[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 256.480 2800.000 257.040 ;
    END
  END x_start[116]
  PIN x_start[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 257.600 2800.000 258.160 ;
    END
  END x_start[117]
  PIN x_start[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 258.720 2800.000 259.280 ;
    END
  END x_start[118]
  PIN x_start[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 259.840 2800.000 260.400 ;
    END
  END x_start[119]
  PIN x_start[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 138.880 2800.000 139.440 ;
    END
  END x_start[11]
  PIN x_start[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 260.960 2800.000 261.520 ;
    END
  END x_start[120]
  PIN x_start[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 262.080 2800.000 262.640 ;
    END
  END x_start[121]
  PIN x_start[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 263.200 2800.000 263.760 ;
    END
  END x_start[122]
  PIN x_start[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 264.320 2800.000 264.880 ;
    END
  END x_start[123]
  PIN x_start[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 265.440 2800.000 266.000 ;
    END
  END x_start[124]
  PIN x_start[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 266.560 2800.000 267.120 ;
    END
  END x_start[125]
  PIN x_start[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 267.680 2800.000 268.240 ;
    END
  END x_start[126]
  PIN x_start[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 268.800 2800.000 269.360 ;
    END
  END x_start[127]
  PIN x_start[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 269.920 2800.000 270.480 ;
    END
  END x_start[128]
  PIN x_start[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 271.040 2800.000 271.600 ;
    END
  END x_start[129]
  PIN x_start[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 140.000 2800.000 140.560 ;
    END
  END x_start[12]
  PIN x_start[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 272.160 2800.000 272.720 ;
    END
  END x_start[130]
  PIN x_start[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 273.280 2800.000 273.840 ;
    END
  END x_start[131]
  PIN x_start[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 274.400 2800.000 274.960 ;
    END
  END x_start[132]
  PIN x_start[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 275.520 2800.000 276.080 ;
    END
  END x_start[133]
  PIN x_start[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 276.640 2800.000 277.200 ;
    END
  END x_start[134]
  PIN x_start[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 277.760 2800.000 278.320 ;
    END
  END x_start[135]
  PIN x_start[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 278.880 2800.000 279.440 ;
    END
  END x_start[136]
  PIN x_start[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 280.000 2800.000 280.560 ;
    END
  END x_start[137]
  PIN x_start[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 281.120 2800.000 281.680 ;
    END
  END x_start[138]
  PIN x_start[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 282.240 2800.000 282.800 ;
    END
  END x_start[139]
  PIN x_start[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 141.120 2800.000 141.680 ;
    END
  END x_start[13]
  PIN x_start[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 283.360 2800.000 283.920 ;
    END
  END x_start[140]
  PIN x_start[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 284.480 2800.000 285.040 ;
    END
  END x_start[141]
  PIN x_start[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 285.600 2800.000 286.160 ;
    END
  END x_start[142]
  PIN x_start[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 286.720 2800.000 287.280 ;
    END
  END x_start[143]
  PIN x_start[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 287.840 2800.000 288.400 ;
    END
  END x_start[144]
  PIN x_start[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 288.960 2800.000 289.520 ;
    END
  END x_start[145]
  PIN x_start[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 290.080 2800.000 290.640 ;
    END
  END x_start[146]
  PIN x_start[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 291.200 2800.000 291.760 ;
    END
  END x_start[147]
  PIN x_start[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 292.320 2800.000 292.880 ;
    END
  END x_start[148]
  PIN x_start[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 293.440 2800.000 294.000 ;
    END
  END x_start[149]
  PIN x_start[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 142.240 2800.000 142.800 ;
    END
  END x_start[14]
  PIN x_start[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 294.560 2800.000 295.120 ;
    END
  END x_start[150]
  PIN x_start[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 295.680 2800.000 296.240 ;
    END
  END x_start[151]
  PIN x_start[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 296.800 2800.000 297.360 ;
    END
  END x_start[152]
  PIN x_start[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 297.920 2800.000 298.480 ;
    END
  END x_start[153]
  PIN x_start[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 299.040 2800.000 299.600 ;
    END
  END x_start[154]
  PIN x_start[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 300.160 2800.000 300.720 ;
    END
  END x_start[155]
  PIN x_start[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 301.280 2800.000 301.840 ;
    END
  END x_start[156]
  PIN x_start[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 302.400 2800.000 302.960 ;
    END
  END x_start[157]
  PIN x_start[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 303.520 2800.000 304.080 ;
    END
  END x_start[158]
  PIN x_start[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 304.640 2800.000 305.200 ;
    END
  END x_start[159]
  PIN x_start[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 143.360 2800.000 143.920 ;
    END
  END x_start[15]
  PIN x_start[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 305.760 2800.000 306.320 ;
    END
  END x_start[160]
  PIN x_start[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 306.880 2800.000 307.440 ;
    END
  END x_start[161]
  PIN x_start[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 308.000 2800.000 308.560 ;
    END
  END x_start[162]
  PIN x_start[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 309.120 2800.000 309.680 ;
    END
  END x_start[163]
  PIN x_start[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 310.240 2800.000 310.800 ;
    END
  END x_start[164]
  PIN x_start[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 311.360 2800.000 311.920 ;
    END
  END x_start[165]
  PIN x_start[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 312.480 2800.000 313.040 ;
    END
  END x_start[166]
  PIN x_start[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 313.600 2800.000 314.160 ;
    END
  END x_start[167]
  PIN x_start[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 314.720 2800.000 315.280 ;
    END
  END x_start[168]
  PIN x_start[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 315.840 2800.000 316.400 ;
    END
  END x_start[169]
  PIN x_start[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 144.480 2800.000 145.040 ;
    END
  END x_start[16]
  PIN x_start[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 316.960 2800.000 317.520 ;
    END
  END x_start[170]
  PIN x_start[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 318.080 2800.000 318.640 ;
    END
  END x_start[171]
  PIN x_start[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 319.200 2800.000 319.760 ;
    END
  END x_start[172]
  PIN x_start[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 320.320 2800.000 320.880 ;
    END
  END x_start[173]
  PIN x_start[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 321.440 2800.000 322.000 ;
    END
  END x_start[174]
  PIN x_start[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 322.560 2800.000 323.120 ;
    END
  END x_start[175]
  PIN x_start[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 323.680 2800.000 324.240 ;
    END
  END x_start[176]
  PIN x_start[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 324.800 2800.000 325.360 ;
    END
  END x_start[177]
  PIN x_start[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 325.920 2800.000 326.480 ;
    END
  END x_start[178]
  PIN x_start[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 327.040 2800.000 327.600 ;
    END
  END x_start[179]
  PIN x_start[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 145.600 2800.000 146.160 ;
    END
  END x_start[17]
  PIN x_start[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 328.160 2800.000 328.720 ;
    END
  END x_start[180]
  PIN x_start[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 329.280 2800.000 329.840 ;
    END
  END x_start[181]
  PIN x_start[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 330.400 2800.000 330.960 ;
    END
  END x_start[182]
  PIN x_start[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 331.520 2800.000 332.080 ;
    END
  END x_start[183]
  PIN x_start[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 332.640 2800.000 333.200 ;
    END
  END x_start[184]
  PIN x_start[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 333.760 2800.000 334.320 ;
    END
  END x_start[185]
  PIN x_start[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 334.880 2800.000 335.440 ;
    END
  END x_start[186]
  PIN x_start[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 336.000 2800.000 336.560 ;
    END
  END x_start[187]
  PIN x_start[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 337.120 2800.000 337.680 ;
    END
  END x_start[188]
  PIN x_start[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 338.240 2800.000 338.800 ;
    END
  END x_start[189]
  PIN x_start[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 146.720 2800.000 147.280 ;
    END
  END x_start[18]
  PIN x_start[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 339.360 2800.000 339.920 ;
    END
  END x_start[190]
  PIN x_start[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 340.480 2800.000 341.040 ;
    END
  END x_start[191]
  PIN x_start[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 341.600 2800.000 342.160 ;
    END
  END x_start[192]
  PIN x_start[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 342.720 2800.000 343.280 ;
    END
  END x_start[193]
  PIN x_start[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 343.840 2800.000 344.400 ;
    END
  END x_start[194]
  PIN x_start[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 344.960 2800.000 345.520 ;
    END
  END x_start[195]
  PIN x_start[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 346.080 2800.000 346.640 ;
    END
  END x_start[196]
  PIN x_start[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 347.200 2800.000 347.760 ;
    END
  END x_start[197]
  PIN x_start[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 348.320 2800.000 348.880 ;
    END
  END x_start[198]
  PIN x_start[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 349.440 2800.000 350.000 ;
    END
  END x_start[199]
  PIN x_start[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 147.840 2800.000 148.400 ;
    END
  END x_start[19]
  PIN x_start[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 127.680 2800.000 128.240 ;
    END
  END x_start[1]
  PIN x_start[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 350.560 2800.000 351.120 ;
    END
  END x_start[200]
  PIN x_start[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 351.680 2800.000 352.240 ;
    END
  END x_start[201]
  PIN x_start[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 352.800 2800.000 353.360 ;
    END
  END x_start[202]
  PIN x_start[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 353.920 2800.000 354.480 ;
    END
  END x_start[203]
  PIN x_start[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 355.040 2800.000 355.600 ;
    END
  END x_start[204]
  PIN x_start[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 356.160 2800.000 356.720 ;
    END
  END x_start[205]
  PIN x_start[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 357.280 2800.000 357.840 ;
    END
  END x_start[206]
  PIN x_start[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 358.400 2800.000 358.960 ;
    END
  END x_start[207]
  PIN x_start[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 359.520 2800.000 360.080 ;
    END
  END x_start[208]
  PIN x_start[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 360.640 2800.000 361.200 ;
    END
  END x_start[209]
  PIN x_start[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 148.960 2800.000 149.520 ;
    END
  END x_start[20]
  PIN x_start[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 361.760 2800.000 362.320 ;
    END
  END x_start[210]
  PIN x_start[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 362.880 2800.000 363.440 ;
    END
  END x_start[211]
  PIN x_start[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 364.000 2800.000 364.560 ;
    END
  END x_start[212]
  PIN x_start[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 365.120 2800.000 365.680 ;
    END
  END x_start[213]
  PIN x_start[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 366.240 2800.000 366.800 ;
    END
  END x_start[214]
  PIN x_start[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 367.360 2800.000 367.920 ;
    END
  END x_start[215]
  PIN x_start[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 368.480 2800.000 369.040 ;
    END
  END x_start[216]
  PIN x_start[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 369.600 2800.000 370.160 ;
    END
  END x_start[217]
  PIN x_start[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 370.720 2800.000 371.280 ;
    END
  END x_start[218]
  PIN x_start[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 371.840 2800.000 372.400 ;
    END
  END x_start[219]
  PIN x_start[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 150.080 2800.000 150.640 ;
    END
  END x_start[21]
  PIN x_start[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 372.960 2800.000 373.520 ;
    END
  END x_start[220]
  PIN x_start[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 374.080 2800.000 374.640 ;
    END
  END x_start[221]
  PIN x_start[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 375.200 2800.000 375.760 ;
    END
  END x_start[222]
  PIN x_start[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 376.320 2800.000 376.880 ;
    END
  END x_start[223]
  PIN x_start[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 377.440 2800.000 378.000 ;
    END
  END x_start[224]
  PIN x_start[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 378.560 2800.000 379.120 ;
    END
  END x_start[225]
  PIN x_start[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 379.680 2800.000 380.240 ;
    END
  END x_start[226]
  PIN x_start[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 380.800 2800.000 381.360 ;
    END
  END x_start[227]
  PIN x_start[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 381.920 2800.000 382.480 ;
    END
  END x_start[228]
  PIN x_start[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 383.040 2800.000 383.600 ;
    END
  END x_start[229]
  PIN x_start[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 151.200 2800.000 151.760 ;
    END
  END x_start[22]
  PIN x_start[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 384.160 2800.000 384.720 ;
    END
  END x_start[230]
  PIN x_start[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 385.280 2800.000 385.840 ;
    END
  END x_start[231]
  PIN x_start[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 386.400 2800.000 386.960 ;
    END
  END x_start[232]
  PIN x_start[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 387.520 2800.000 388.080 ;
    END
  END x_start[233]
  PIN x_start[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 388.640 2800.000 389.200 ;
    END
  END x_start[234]
  PIN x_start[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 389.760 2800.000 390.320 ;
    END
  END x_start[235]
  PIN x_start[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 390.880 2800.000 391.440 ;
    END
  END x_start[236]
  PIN x_start[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 392.000 2800.000 392.560 ;
    END
  END x_start[237]
  PIN x_start[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 393.120 2800.000 393.680 ;
    END
  END x_start[238]
  PIN x_start[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 394.240 2800.000 394.800 ;
    END
  END x_start[239]
  PIN x_start[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 152.320 2800.000 152.880 ;
    END
  END x_start[23]
  PIN x_start[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 395.360 2800.000 395.920 ;
    END
  END x_start[240]
  PIN x_start[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 396.480 2800.000 397.040 ;
    END
  END x_start[241]
  PIN x_start[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 397.600 2800.000 398.160 ;
    END
  END x_start[242]
  PIN x_start[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 398.720 2800.000 399.280 ;
    END
  END x_start[243]
  PIN x_start[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 399.840 2800.000 400.400 ;
    END
  END x_start[244]
  PIN x_start[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 400.960 2800.000 401.520 ;
    END
  END x_start[245]
  PIN x_start[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 402.080 2800.000 402.640 ;
    END
  END x_start[246]
  PIN x_start[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 403.200 2800.000 403.760 ;
    END
  END x_start[247]
  PIN x_start[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 404.320 2800.000 404.880 ;
    END
  END x_start[248]
  PIN x_start[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 405.440 2800.000 406.000 ;
    END
  END x_start[249]
  PIN x_start[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 153.440 2800.000 154.000 ;
    END
  END x_start[24]
  PIN x_start[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 406.560 2800.000 407.120 ;
    END
  END x_start[250]
  PIN x_start[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 407.680 2800.000 408.240 ;
    END
  END x_start[251]
  PIN x_start[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 408.800 2800.000 409.360 ;
    END
  END x_start[252]
  PIN x_start[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 409.920 2800.000 410.480 ;
    END
  END x_start[253]
  PIN x_start[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 411.040 2800.000 411.600 ;
    END
  END x_start[254]
  PIN x_start[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 412.160 2800.000 412.720 ;
    END
  END x_start[255]
  PIN x_start[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 413.280 2800.000 413.840 ;
    END
  END x_start[256]
  PIN x_start[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 414.400 2800.000 414.960 ;
    END
  END x_start[257]
  PIN x_start[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 415.520 2800.000 416.080 ;
    END
  END x_start[258]
  PIN x_start[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 416.640 2800.000 417.200 ;
    END
  END x_start[259]
  PIN x_start[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 154.560 2800.000 155.120 ;
    END
  END x_start[25]
  PIN x_start[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 417.760 2800.000 418.320 ;
    END
  END x_start[260]
  PIN x_start[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 418.880 2800.000 419.440 ;
    END
  END x_start[261]
  PIN x_start[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 420.000 2800.000 420.560 ;
    END
  END x_start[262]
  PIN x_start[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 421.120 2800.000 421.680 ;
    END
  END x_start[263]
  PIN x_start[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 422.240 2800.000 422.800 ;
    END
  END x_start[264]
  PIN x_start[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 423.360 2800.000 423.920 ;
    END
  END x_start[265]
  PIN x_start[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 424.480 2800.000 425.040 ;
    END
  END x_start[266]
  PIN x_start[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 425.600 2800.000 426.160 ;
    END
  END x_start[267]
  PIN x_start[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 426.720 2800.000 427.280 ;
    END
  END x_start[268]
  PIN x_start[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 427.840 2800.000 428.400 ;
    END
  END x_start[269]
  PIN x_start[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 155.680 2800.000 156.240 ;
    END
  END x_start[26]
  PIN x_start[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 428.960 2800.000 429.520 ;
    END
  END x_start[270]
  PIN x_start[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 430.080 2800.000 430.640 ;
    END
  END x_start[271]
  PIN x_start[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 431.200 2800.000 431.760 ;
    END
  END x_start[272]
  PIN x_start[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 432.320 2800.000 432.880 ;
    END
  END x_start[273]
  PIN x_start[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 433.440 2800.000 434.000 ;
    END
  END x_start[274]
  PIN x_start[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 434.560 2800.000 435.120 ;
    END
  END x_start[275]
  PIN x_start[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 435.680 2800.000 436.240 ;
    END
  END x_start[276]
  PIN x_start[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 436.800 2800.000 437.360 ;
    END
  END x_start[277]
  PIN x_start[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 437.920 2800.000 438.480 ;
    END
  END x_start[278]
  PIN x_start[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 439.040 2800.000 439.600 ;
    END
  END x_start[279]
  PIN x_start[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 156.800 2800.000 157.360 ;
    END
  END x_start[27]
  PIN x_start[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 440.160 2800.000 440.720 ;
    END
  END x_start[280]
  PIN x_start[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 441.280 2800.000 441.840 ;
    END
  END x_start[281]
  PIN x_start[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 442.400 2800.000 442.960 ;
    END
  END x_start[282]
  PIN x_start[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 443.520 2800.000 444.080 ;
    END
  END x_start[283]
  PIN x_start[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 444.640 2800.000 445.200 ;
    END
  END x_start[284]
  PIN x_start[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 445.760 2800.000 446.320 ;
    END
  END x_start[285]
  PIN x_start[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 446.880 2800.000 447.440 ;
    END
  END x_start[286]
  PIN x_start[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 448.000 2800.000 448.560 ;
    END
  END x_start[287]
  PIN x_start[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 449.120 2800.000 449.680 ;
    END
  END x_start[288]
  PIN x_start[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 450.240 2800.000 450.800 ;
    END
  END x_start[289]
  PIN x_start[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 157.920 2800.000 158.480 ;
    END
  END x_start[28]
  PIN x_start[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 451.360 2800.000 451.920 ;
    END
  END x_start[290]
  PIN x_start[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 452.480 2800.000 453.040 ;
    END
  END x_start[291]
  PIN x_start[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 453.600 2800.000 454.160 ;
    END
  END x_start[292]
  PIN x_start[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 454.720 2800.000 455.280 ;
    END
  END x_start[293]
  PIN x_start[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 455.840 2800.000 456.400 ;
    END
  END x_start[294]
  PIN x_start[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 456.960 2800.000 457.520 ;
    END
  END x_start[295]
  PIN x_start[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 458.080 2800.000 458.640 ;
    END
  END x_start[296]
  PIN x_start[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 459.200 2800.000 459.760 ;
    END
  END x_start[297]
  PIN x_start[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 460.320 2800.000 460.880 ;
    END
  END x_start[298]
  PIN x_start[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 461.440 2800.000 462.000 ;
    END
  END x_start[299]
  PIN x_start[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 159.040 2800.000 159.600 ;
    END
  END x_start[29]
  PIN x_start[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 128.800 2800.000 129.360 ;
    END
  END x_start[2]
  PIN x_start[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 462.560 2800.000 463.120 ;
    END
  END x_start[300]
  PIN x_start[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 463.680 2800.000 464.240 ;
    END
  END x_start[301]
  PIN x_start[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 464.800 2800.000 465.360 ;
    END
  END x_start[302]
  PIN x_start[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 465.920 2800.000 466.480 ;
    END
  END x_start[303]
  PIN x_start[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 467.040 2800.000 467.600 ;
    END
  END x_start[304]
  PIN x_start[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 468.160 2800.000 468.720 ;
    END
  END x_start[305]
  PIN x_start[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 469.280 2800.000 469.840 ;
    END
  END x_start[306]
  PIN x_start[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 470.400 2800.000 470.960 ;
    END
  END x_start[307]
  PIN x_start[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 471.520 2800.000 472.080 ;
    END
  END x_start[308]
  PIN x_start[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 472.640 2800.000 473.200 ;
    END
  END x_start[309]
  PIN x_start[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 160.160 2800.000 160.720 ;
    END
  END x_start[30]
  PIN x_start[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 473.760 2800.000 474.320 ;
    END
  END x_start[310]
  PIN x_start[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 474.880 2800.000 475.440 ;
    END
  END x_start[311]
  PIN x_start[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 476.000 2800.000 476.560 ;
    END
  END x_start[312]
  PIN x_start[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 477.120 2800.000 477.680 ;
    END
  END x_start[313]
  PIN x_start[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 478.240 2800.000 478.800 ;
    END
  END x_start[314]
  PIN x_start[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 479.360 2800.000 479.920 ;
    END
  END x_start[315]
  PIN x_start[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 480.480 2800.000 481.040 ;
    END
  END x_start[316]
  PIN x_start[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 481.600 2800.000 482.160 ;
    END
  END x_start[317]
  PIN x_start[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 482.720 2800.000 483.280 ;
    END
  END x_start[318]
  PIN x_start[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 483.840 2800.000 484.400 ;
    END
  END x_start[319]
  PIN x_start[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 161.280 2800.000 161.840 ;
    END
  END x_start[31]
  PIN x_start[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 484.960 2800.000 485.520 ;
    END
  END x_start[320]
  PIN x_start[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 486.080 2800.000 486.640 ;
    END
  END x_start[321]
  PIN x_start[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 487.200 2800.000 487.760 ;
    END
  END x_start[322]
  PIN x_start[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 488.320 2800.000 488.880 ;
    END
  END x_start[323]
  PIN x_start[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 489.440 2800.000 490.000 ;
    END
  END x_start[324]
  PIN x_start[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 490.560 2800.000 491.120 ;
    END
  END x_start[325]
  PIN x_start[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 491.680 2800.000 492.240 ;
    END
  END x_start[326]
  PIN x_start[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 492.800 2800.000 493.360 ;
    END
  END x_start[327]
  PIN x_start[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 493.920 2800.000 494.480 ;
    END
  END x_start[328]
  PIN x_start[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 495.040 2800.000 495.600 ;
    END
  END x_start[329]
  PIN x_start[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 162.400 2800.000 162.960 ;
    END
  END x_start[32]
  PIN x_start[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 496.160 2800.000 496.720 ;
    END
  END x_start[330]
  PIN x_start[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 497.280 2800.000 497.840 ;
    END
  END x_start[331]
  PIN x_start[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 498.400 2800.000 498.960 ;
    END
  END x_start[332]
  PIN x_start[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 499.520 2800.000 500.080 ;
    END
  END x_start[333]
  PIN x_start[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 500.640 2800.000 501.200 ;
    END
  END x_start[334]
  PIN x_start[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 501.760 2800.000 502.320 ;
    END
  END x_start[335]
  PIN x_start[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 502.880 2800.000 503.440 ;
    END
  END x_start[336]
  PIN x_start[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 504.000 2800.000 504.560 ;
    END
  END x_start[337]
  PIN x_start[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 505.120 2800.000 505.680 ;
    END
  END x_start[338]
  PIN x_start[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 506.240 2800.000 506.800 ;
    END
  END x_start[339]
  PIN x_start[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 163.520 2800.000 164.080 ;
    END
  END x_start[33]
  PIN x_start[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 507.360 2800.000 507.920 ;
    END
  END x_start[340]
  PIN x_start[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 508.480 2800.000 509.040 ;
    END
  END x_start[341]
  PIN x_start[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 509.600 2800.000 510.160 ;
    END
  END x_start[342]
  PIN x_start[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 510.720 2800.000 511.280 ;
    END
  END x_start[343]
  PIN x_start[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 511.840 2800.000 512.400 ;
    END
  END x_start[344]
  PIN x_start[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 512.960 2800.000 513.520 ;
    END
  END x_start[345]
  PIN x_start[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 514.080 2800.000 514.640 ;
    END
  END x_start[346]
  PIN x_start[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 515.200 2800.000 515.760 ;
    END
  END x_start[347]
  PIN x_start[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 516.320 2800.000 516.880 ;
    END
  END x_start[348]
  PIN x_start[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 517.440 2800.000 518.000 ;
    END
  END x_start[349]
  PIN x_start[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 164.640 2800.000 165.200 ;
    END
  END x_start[34]
  PIN x_start[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 518.560 2800.000 519.120 ;
    END
  END x_start[350]
  PIN x_start[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 519.680 2800.000 520.240 ;
    END
  END x_start[351]
  PIN x_start[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 520.800 2800.000 521.360 ;
    END
  END x_start[352]
  PIN x_start[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 521.920 2800.000 522.480 ;
    END
  END x_start[353]
  PIN x_start[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 523.040 2800.000 523.600 ;
    END
  END x_start[354]
  PIN x_start[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 524.160 2800.000 524.720 ;
    END
  END x_start[355]
  PIN x_start[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 525.280 2800.000 525.840 ;
    END
  END x_start[356]
  PIN x_start[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 526.400 2800.000 526.960 ;
    END
  END x_start[357]
  PIN x_start[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 527.520 2800.000 528.080 ;
    END
  END x_start[358]
  PIN x_start[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 528.640 2800.000 529.200 ;
    END
  END x_start[359]
  PIN x_start[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 165.760 2800.000 166.320 ;
    END
  END x_start[35]
  PIN x_start[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 529.760 2800.000 530.320 ;
    END
  END x_start[360]
  PIN x_start[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 530.880 2800.000 531.440 ;
    END
  END x_start[361]
  PIN x_start[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 532.000 2800.000 532.560 ;
    END
  END x_start[362]
  PIN x_start[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 533.120 2800.000 533.680 ;
    END
  END x_start[363]
  PIN x_start[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 534.240 2800.000 534.800 ;
    END
  END x_start[364]
  PIN x_start[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 535.360 2800.000 535.920 ;
    END
  END x_start[365]
  PIN x_start[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 536.480 2800.000 537.040 ;
    END
  END x_start[366]
  PIN x_start[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 537.600 2800.000 538.160 ;
    END
  END x_start[367]
  PIN x_start[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 538.720 2800.000 539.280 ;
    END
  END x_start[368]
  PIN x_start[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 539.840 2800.000 540.400 ;
    END
  END x_start[369]
  PIN x_start[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 166.880 2800.000 167.440 ;
    END
  END x_start[36]
  PIN x_start[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 540.960 2800.000 541.520 ;
    END
  END x_start[370]
  PIN x_start[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 542.080 2800.000 542.640 ;
    END
  END x_start[371]
  PIN x_start[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 543.200 2800.000 543.760 ;
    END
  END x_start[372]
  PIN x_start[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 544.320 2800.000 544.880 ;
    END
  END x_start[373]
  PIN x_start[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 545.440 2800.000 546.000 ;
    END
  END x_start[374]
  PIN x_start[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 546.560 2800.000 547.120 ;
    END
  END x_start[375]
  PIN x_start[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 547.680 2800.000 548.240 ;
    END
  END x_start[376]
  PIN x_start[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 548.800 2800.000 549.360 ;
    END
  END x_start[377]
  PIN x_start[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 549.920 2800.000 550.480 ;
    END
  END x_start[378]
  PIN x_start[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 551.040 2800.000 551.600 ;
    END
  END x_start[379]
  PIN x_start[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 168.000 2800.000 168.560 ;
    END
  END x_start[37]
  PIN x_start[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 552.160 2800.000 552.720 ;
    END
  END x_start[380]
  PIN x_start[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 553.280 2800.000 553.840 ;
    END
  END x_start[381]
  PIN x_start[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 554.400 2800.000 554.960 ;
    END
  END x_start[382]
  PIN x_start[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 555.520 2800.000 556.080 ;
    END
  END x_start[383]
  PIN x_start[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 556.640 2800.000 557.200 ;
    END
  END x_start[384]
  PIN x_start[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 557.760 2800.000 558.320 ;
    END
  END x_start[385]
  PIN x_start[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 558.880 2800.000 559.440 ;
    END
  END x_start[386]
  PIN x_start[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 560.000 2800.000 560.560 ;
    END
  END x_start[387]
  PIN x_start[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 561.120 2800.000 561.680 ;
    END
  END x_start[388]
  PIN x_start[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 562.240 2800.000 562.800 ;
    END
  END x_start[389]
  PIN x_start[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 169.120 2800.000 169.680 ;
    END
  END x_start[38]
  PIN x_start[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 563.360 2800.000 563.920 ;
    END
  END x_start[390]
  PIN x_start[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 564.480 2800.000 565.040 ;
    END
  END x_start[391]
  PIN x_start[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 565.600 2800.000 566.160 ;
    END
  END x_start[392]
  PIN x_start[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 566.720 2800.000 567.280 ;
    END
  END x_start[393]
  PIN x_start[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 567.840 2800.000 568.400 ;
    END
  END x_start[394]
  PIN x_start[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 568.960 2800.000 569.520 ;
    END
  END x_start[395]
  PIN x_start[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 570.080 2800.000 570.640 ;
    END
  END x_start[396]
  PIN x_start[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 571.200 2800.000 571.760 ;
    END
  END x_start[397]
  PIN x_start[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 572.320 2800.000 572.880 ;
    END
  END x_start[398]
  PIN x_start[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 573.440 2800.000 574.000 ;
    END
  END x_start[399]
  PIN x_start[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 170.240 2800.000 170.800 ;
    END
  END x_start[39]
  PIN x_start[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 129.920 2800.000 130.480 ;
    END
  END x_start[3]
  PIN x_start[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 574.560 2800.000 575.120 ;
    END
  END x_start[400]
  PIN x_start[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 575.680 2800.000 576.240 ;
    END
  END x_start[401]
  PIN x_start[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 576.800 2800.000 577.360 ;
    END
  END x_start[402]
  PIN x_start[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 577.920 2800.000 578.480 ;
    END
  END x_start[403]
  PIN x_start[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 579.040 2800.000 579.600 ;
    END
  END x_start[404]
  PIN x_start[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 580.160 2800.000 580.720 ;
    END
  END x_start[405]
  PIN x_start[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 581.280 2800.000 581.840 ;
    END
  END x_start[406]
  PIN x_start[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 582.400 2800.000 582.960 ;
    END
  END x_start[407]
  PIN x_start[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 583.520 2800.000 584.080 ;
    END
  END x_start[408]
  PIN x_start[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 584.640 2800.000 585.200 ;
    END
  END x_start[409]
  PIN x_start[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 171.360 2800.000 171.920 ;
    END
  END x_start[40]
  PIN x_start[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 585.760 2800.000 586.320 ;
    END
  END x_start[410]
  PIN x_start[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 586.880 2800.000 587.440 ;
    END
  END x_start[411]
  PIN x_start[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 588.000 2800.000 588.560 ;
    END
  END x_start[412]
  PIN x_start[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 589.120 2800.000 589.680 ;
    END
  END x_start[413]
  PIN x_start[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 590.240 2800.000 590.800 ;
    END
  END x_start[414]
  PIN x_start[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 591.360 2800.000 591.920 ;
    END
  END x_start[415]
  PIN x_start[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 592.480 2800.000 593.040 ;
    END
  END x_start[416]
  PIN x_start[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 593.600 2800.000 594.160 ;
    END
  END x_start[417]
  PIN x_start[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 594.720 2800.000 595.280 ;
    END
  END x_start[418]
  PIN x_start[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 595.840 2800.000 596.400 ;
    END
  END x_start[419]
  PIN x_start[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 172.480 2800.000 173.040 ;
    END
  END x_start[41]
  PIN x_start[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 596.960 2800.000 597.520 ;
    END
  END x_start[420]
  PIN x_start[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 598.080 2800.000 598.640 ;
    END
  END x_start[421]
  PIN x_start[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 599.200 2800.000 599.760 ;
    END
  END x_start[422]
  PIN x_start[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 600.320 2800.000 600.880 ;
    END
  END x_start[423]
  PIN x_start[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 601.440 2800.000 602.000 ;
    END
  END x_start[424]
  PIN x_start[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 602.560 2800.000 603.120 ;
    END
  END x_start[425]
  PIN x_start[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 603.680 2800.000 604.240 ;
    END
  END x_start[426]
  PIN x_start[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 604.800 2800.000 605.360 ;
    END
  END x_start[427]
  PIN x_start[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 605.920 2800.000 606.480 ;
    END
  END x_start[428]
  PIN x_start[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 607.040 2800.000 607.600 ;
    END
  END x_start[429]
  PIN x_start[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 173.600 2800.000 174.160 ;
    END
  END x_start[42]
  PIN x_start[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 608.160 2800.000 608.720 ;
    END
  END x_start[430]
  PIN x_start[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 609.280 2800.000 609.840 ;
    END
  END x_start[431]
  PIN x_start[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 610.400 2800.000 610.960 ;
    END
  END x_start[432]
  PIN x_start[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 611.520 2800.000 612.080 ;
    END
  END x_start[433]
  PIN x_start[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 612.640 2800.000 613.200 ;
    END
  END x_start[434]
  PIN x_start[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 613.760 2800.000 614.320 ;
    END
  END x_start[435]
  PIN x_start[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 614.880 2800.000 615.440 ;
    END
  END x_start[436]
  PIN x_start[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 616.000 2800.000 616.560 ;
    END
  END x_start[437]
  PIN x_start[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 617.120 2800.000 617.680 ;
    END
  END x_start[438]
  PIN x_start[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 618.240 2800.000 618.800 ;
    END
  END x_start[439]
  PIN x_start[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 174.720 2800.000 175.280 ;
    END
  END x_start[43]
  PIN x_start[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 619.360 2800.000 619.920 ;
    END
  END x_start[440]
  PIN x_start[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 620.480 2800.000 621.040 ;
    END
  END x_start[441]
  PIN x_start[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 621.600 2800.000 622.160 ;
    END
  END x_start[442]
  PIN x_start[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 622.720 2800.000 623.280 ;
    END
  END x_start[443]
  PIN x_start[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 623.840 2800.000 624.400 ;
    END
  END x_start[444]
  PIN x_start[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 624.960 2800.000 625.520 ;
    END
  END x_start[445]
  PIN x_start[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 626.080 2800.000 626.640 ;
    END
  END x_start[446]
  PIN x_start[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 627.200 2800.000 627.760 ;
    END
  END x_start[447]
  PIN x_start[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 628.320 2800.000 628.880 ;
    END
  END x_start[448]
  PIN x_start[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 629.440 2800.000 630.000 ;
    END
  END x_start[449]
  PIN x_start[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 175.840 2800.000 176.400 ;
    END
  END x_start[44]
  PIN x_start[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 630.560 2800.000 631.120 ;
    END
  END x_start[450]
  PIN x_start[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 631.680 2800.000 632.240 ;
    END
  END x_start[451]
  PIN x_start[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 632.800 2800.000 633.360 ;
    END
  END x_start[452]
  PIN x_start[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 633.920 2800.000 634.480 ;
    END
  END x_start[453]
  PIN x_start[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 635.040 2800.000 635.600 ;
    END
  END x_start[454]
  PIN x_start[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 636.160 2800.000 636.720 ;
    END
  END x_start[455]
  PIN x_start[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 637.280 2800.000 637.840 ;
    END
  END x_start[456]
  PIN x_start[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 638.400 2800.000 638.960 ;
    END
  END x_start[457]
  PIN x_start[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 639.520 2800.000 640.080 ;
    END
  END x_start[458]
  PIN x_start[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 640.640 2800.000 641.200 ;
    END
  END x_start[459]
  PIN x_start[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 176.960 2800.000 177.520 ;
    END
  END x_start[45]
  PIN x_start[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 641.760 2800.000 642.320 ;
    END
  END x_start[460]
  PIN x_start[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 642.880 2800.000 643.440 ;
    END
  END x_start[461]
  PIN x_start[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 644.000 2800.000 644.560 ;
    END
  END x_start[462]
  PIN x_start[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 645.120 2800.000 645.680 ;
    END
  END x_start[463]
  PIN x_start[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 646.240 2800.000 646.800 ;
    END
  END x_start[464]
  PIN x_start[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 647.360 2800.000 647.920 ;
    END
  END x_start[465]
  PIN x_start[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 648.480 2800.000 649.040 ;
    END
  END x_start[466]
  PIN x_start[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 649.600 2800.000 650.160 ;
    END
  END x_start[467]
  PIN x_start[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 650.720 2800.000 651.280 ;
    END
  END x_start[468]
  PIN x_start[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 651.840 2800.000 652.400 ;
    END
  END x_start[469]
  PIN x_start[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 178.080 2800.000 178.640 ;
    END
  END x_start[46]
  PIN x_start[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 652.960 2800.000 653.520 ;
    END
  END x_start[470]
  PIN x_start[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 654.080 2800.000 654.640 ;
    END
  END x_start[471]
  PIN x_start[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 655.200 2800.000 655.760 ;
    END
  END x_start[472]
  PIN x_start[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 656.320 2800.000 656.880 ;
    END
  END x_start[473]
  PIN x_start[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 657.440 2800.000 658.000 ;
    END
  END x_start[474]
  PIN x_start[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 658.560 2800.000 659.120 ;
    END
  END x_start[475]
  PIN x_start[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 659.680 2800.000 660.240 ;
    END
  END x_start[476]
  PIN x_start[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 660.800 2800.000 661.360 ;
    END
  END x_start[477]
  PIN x_start[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 661.920 2800.000 662.480 ;
    END
  END x_start[478]
  PIN x_start[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 663.040 2800.000 663.600 ;
    END
  END x_start[479]
  PIN x_start[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 179.200 2800.000 179.760 ;
    END
  END x_start[47]
  PIN x_start[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 664.160 2800.000 664.720 ;
    END
  END x_start[480]
  PIN x_start[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 665.280 2800.000 665.840 ;
    END
  END x_start[481]
  PIN x_start[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 666.400 2800.000 666.960 ;
    END
  END x_start[482]
  PIN x_start[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 667.520 2800.000 668.080 ;
    END
  END x_start[483]
  PIN x_start[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 668.640 2800.000 669.200 ;
    END
  END x_start[484]
  PIN x_start[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 669.760 2800.000 670.320 ;
    END
  END x_start[485]
  PIN x_start[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 670.880 2800.000 671.440 ;
    END
  END x_start[486]
  PIN x_start[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 672.000 2800.000 672.560 ;
    END
  END x_start[487]
  PIN x_start[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 673.120 2800.000 673.680 ;
    END
  END x_start[488]
  PIN x_start[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 674.240 2800.000 674.800 ;
    END
  END x_start[489]
  PIN x_start[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 180.320 2800.000 180.880 ;
    END
  END x_start[48]
  PIN x_start[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 675.360 2800.000 675.920 ;
    END
  END x_start[490]
  PIN x_start[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 676.480 2800.000 677.040 ;
    END
  END x_start[491]
  PIN x_start[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 677.600 2800.000 678.160 ;
    END
  END x_start[492]
  PIN x_start[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 678.720 2800.000 679.280 ;
    END
  END x_start[493]
  PIN x_start[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 679.840 2800.000 680.400 ;
    END
  END x_start[494]
  PIN x_start[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 680.960 2800.000 681.520 ;
    END
  END x_start[495]
  PIN x_start[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 682.080 2800.000 682.640 ;
    END
  END x_start[496]
  PIN x_start[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 683.200 2800.000 683.760 ;
    END
  END x_start[497]
  PIN x_start[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 684.320 2800.000 684.880 ;
    END
  END x_start[498]
  PIN x_start[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 685.440 2800.000 686.000 ;
    END
  END x_start[499]
  PIN x_start[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 181.440 2800.000 182.000 ;
    END
  END x_start[49]
  PIN x_start[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 131.040 2800.000 131.600 ;
    END
  END x_start[4]
  PIN x_start[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 686.560 2800.000 687.120 ;
    END
  END x_start[500]
  PIN x_start[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 687.680 2800.000 688.240 ;
    END
  END x_start[501]
  PIN x_start[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 688.800 2800.000 689.360 ;
    END
  END x_start[502]
  PIN x_start[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 689.920 2800.000 690.480 ;
    END
  END x_start[503]
  PIN x_start[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 691.040 2800.000 691.600 ;
    END
  END x_start[504]
  PIN x_start[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 692.160 2800.000 692.720 ;
    END
  END x_start[505]
  PIN x_start[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 693.280 2800.000 693.840 ;
    END
  END x_start[506]
  PIN x_start[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 694.400 2800.000 694.960 ;
    END
  END x_start[507]
  PIN x_start[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 695.520 2800.000 696.080 ;
    END
  END x_start[508]
  PIN x_start[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 696.640 2800.000 697.200 ;
    END
  END x_start[509]
  PIN x_start[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 182.560 2800.000 183.120 ;
    END
  END x_start[50]
  PIN x_start[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 697.760 2800.000 698.320 ;
    END
  END x_start[510]
  PIN x_start[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 698.880 2800.000 699.440 ;
    END
  END x_start[511]
  PIN x_start[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 183.680 2800.000 184.240 ;
    END
  END x_start[51]
  PIN x_start[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 184.800 2800.000 185.360 ;
    END
  END x_start[52]
  PIN x_start[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 185.920 2800.000 186.480 ;
    END
  END x_start[53]
  PIN x_start[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 187.040 2800.000 187.600 ;
    END
  END x_start[54]
  PIN x_start[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 188.160 2800.000 188.720 ;
    END
  END x_start[55]
  PIN x_start[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 189.280 2800.000 189.840 ;
    END
  END x_start[56]
  PIN x_start[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 190.400 2800.000 190.960 ;
    END
  END x_start[57]
  PIN x_start[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 191.520 2800.000 192.080 ;
    END
  END x_start[58]
  PIN x_start[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 192.640 2800.000 193.200 ;
    END
  END x_start[59]
  PIN x_start[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 132.160 2800.000 132.720 ;
    END
  END x_start[5]
  PIN x_start[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 193.760 2800.000 194.320 ;
    END
  END x_start[60]
  PIN x_start[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 194.880 2800.000 195.440 ;
    END
  END x_start[61]
  PIN x_start[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 196.000 2800.000 196.560 ;
    END
  END x_start[62]
  PIN x_start[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 197.120 2800.000 197.680 ;
    END
  END x_start[63]
  PIN x_start[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 198.240 2800.000 198.800 ;
    END
  END x_start[64]
  PIN x_start[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 199.360 2800.000 199.920 ;
    END
  END x_start[65]
  PIN x_start[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 200.480 2800.000 201.040 ;
    END
  END x_start[66]
  PIN x_start[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 201.600 2800.000 202.160 ;
    END
  END x_start[67]
  PIN x_start[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 202.720 2800.000 203.280 ;
    END
  END x_start[68]
  PIN x_start[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 203.840 2800.000 204.400 ;
    END
  END x_start[69]
  PIN x_start[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 133.280 2800.000 133.840 ;
    END
  END x_start[6]
  PIN x_start[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 204.960 2800.000 205.520 ;
    END
  END x_start[70]
  PIN x_start[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 206.080 2800.000 206.640 ;
    END
  END x_start[71]
  PIN x_start[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 207.200 2800.000 207.760 ;
    END
  END x_start[72]
  PIN x_start[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 208.320 2800.000 208.880 ;
    END
  END x_start[73]
  PIN x_start[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 209.440 2800.000 210.000 ;
    END
  END x_start[74]
  PIN x_start[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 210.560 2800.000 211.120 ;
    END
  END x_start[75]
  PIN x_start[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 211.680 2800.000 212.240 ;
    END
  END x_start[76]
  PIN x_start[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 212.800 2800.000 213.360 ;
    END
  END x_start[77]
  PIN x_start[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 213.920 2800.000 214.480 ;
    END
  END x_start[78]
  PIN x_start[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 215.040 2800.000 215.600 ;
    END
  END x_start[79]
  PIN x_start[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 134.400 2800.000 134.960 ;
    END
  END x_start[7]
  PIN x_start[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 216.160 2800.000 216.720 ;
    END
  END x_start[80]
  PIN x_start[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 217.280 2800.000 217.840 ;
    END
  END x_start[81]
  PIN x_start[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 218.400 2800.000 218.960 ;
    END
  END x_start[82]
  PIN x_start[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 219.520 2800.000 220.080 ;
    END
  END x_start[83]
  PIN x_start[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 220.640 2800.000 221.200 ;
    END
  END x_start[84]
  PIN x_start[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 221.760 2800.000 222.320 ;
    END
  END x_start[85]
  PIN x_start[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 222.880 2800.000 223.440 ;
    END
  END x_start[86]
  PIN x_start[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 224.000 2800.000 224.560 ;
    END
  END x_start[87]
  PIN x_start[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 225.120 2800.000 225.680 ;
    END
  END x_start[88]
  PIN x_start[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 226.240 2800.000 226.800 ;
    END
  END x_start[89]
  PIN x_start[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 135.520 2800.000 136.080 ;
    END
  END x_start[8]
  PIN x_start[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 227.360 2800.000 227.920 ;
    END
  END x_start[90]
  PIN x_start[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 228.480 2800.000 229.040 ;
    END
  END x_start[91]
  PIN x_start[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 229.600 2800.000 230.160 ;
    END
  END x_start[92]
  PIN x_start[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 230.720 2800.000 231.280 ;
    END
  END x_start[93]
  PIN x_start[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 231.840 2800.000 232.400 ;
    END
  END x_start[94]
  PIN x_start[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 232.960 2800.000 233.520 ;
    END
  END x_start[95]
  PIN x_start[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 234.080 2800.000 234.640 ;
    END
  END x_start[96]
  PIN x_start[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 235.200 2800.000 235.760 ;
    END
  END x_start[97]
  PIN x_start[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 236.320 2800.000 236.880 ;
    END
  END x_start[98]
  PIN x_start[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 237.440 2800.000 238.000 ;
    END
  END x_start[99]
  PIN x_start[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 136.640 2800.000 137.200 ;
    END
  END x_start[9]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1046.080 0.000 1046.640 4.000 ;
    END
  END y[0]
  PIN y[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1382.080 0.000 1382.640 4.000 ;
    END
  END y[100]
  PIN y[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1385.440 0.000 1386.000 4.000 ;
    END
  END y[101]
  PIN y[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1388.800 0.000 1389.360 4.000 ;
    END
  END y[102]
  PIN y[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1392.160 0.000 1392.720 4.000 ;
    END
  END y[103]
  PIN y[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1395.520 0.000 1396.080 4.000 ;
    END
  END y[104]
  PIN y[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1398.880 0.000 1399.440 4.000 ;
    END
  END y[105]
  PIN y[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1402.240 0.000 1402.800 4.000 ;
    END
  END y[106]
  PIN y[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1405.600 0.000 1406.160 4.000 ;
    END
  END y[107]
  PIN y[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1408.960 0.000 1409.520 4.000 ;
    END
  END y[108]
  PIN y[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1412.320 0.000 1412.880 4.000 ;
    END
  END y[109]
  PIN y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1079.680 0.000 1080.240 4.000 ;
    END
  END y[10]
  PIN y[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1415.680 0.000 1416.240 4.000 ;
    END
  END y[110]
  PIN y[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1419.040 0.000 1419.600 4.000 ;
    END
  END y[111]
  PIN y[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1422.400 0.000 1422.960 4.000 ;
    END
  END y[112]
  PIN y[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1425.760 0.000 1426.320 4.000 ;
    END
  END y[113]
  PIN y[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1429.120 0.000 1429.680 4.000 ;
    END
  END y[114]
  PIN y[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1432.480 0.000 1433.040 4.000 ;
    END
  END y[115]
  PIN y[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1435.840 0.000 1436.400 4.000 ;
    END
  END y[116]
  PIN y[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1439.200 0.000 1439.760 4.000 ;
    END
  END y[117]
  PIN y[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1442.560 0.000 1443.120 4.000 ;
    END
  END y[118]
  PIN y[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1445.920 0.000 1446.480 4.000 ;
    END
  END y[119]
  PIN y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1083.040 0.000 1083.600 4.000 ;
    END
  END y[11]
  PIN y[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1449.280 0.000 1449.840 4.000 ;
    END
  END y[120]
  PIN y[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1452.640 0.000 1453.200 4.000 ;
    END
  END y[121]
  PIN y[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1456.000 0.000 1456.560 4.000 ;
    END
  END y[122]
  PIN y[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1459.360 0.000 1459.920 4.000 ;
    END
  END y[123]
  PIN y[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1462.720 0.000 1463.280 4.000 ;
    END
  END y[124]
  PIN y[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1466.080 0.000 1466.640 4.000 ;
    END
  END y[125]
  PIN y[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1469.440 0.000 1470.000 4.000 ;
    END
  END y[126]
  PIN y[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1472.800 0.000 1473.360 4.000 ;
    END
  END y[127]
  PIN y[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1476.160 0.000 1476.720 4.000 ;
    END
  END y[128]
  PIN y[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1479.520 0.000 1480.080 4.000 ;
    END
  END y[129]
  PIN y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1086.400 0.000 1086.960 4.000 ;
    END
  END y[12]
  PIN y[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1482.880 0.000 1483.440 4.000 ;
    END
  END y[130]
  PIN y[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1486.240 0.000 1486.800 4.000 ;
    END
  END y[131]
  PIN y[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1489.600 0.000 1490.160 4.000 ;
    END
  END y[132]
  PIN y[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1492.960 0.000 1493.520 4.000 ;
    END
  END y[133]
  PIN y[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1496.320 0.000 1496.880 4.000 ;
    END
  END y[134]
  PIN y[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1499.680 0.000 1500.240 4.000 ;
    END
  END y[135]
  PIN y[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1503.040 0.000 1503.600 4.000 ;
    END
  END y[136]
  PIN y[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1506.400 0.000 1506.960 4.000 ;
    END
  END y[137]
  PIN y[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1509.760 0.000 1510.320 4.000 ;
    END
  END y[138]
  PIN y[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1513.120 0.000 1513.680 4.000 ;
    END
  END y[139]
  PIN y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1089.760 0.000 1090.320 4.000 ;
    END
  END y[13]
  PIN y[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1516.480 0.000 1517.040 4.000 ;
    END
  END y[140]
  PIN y[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1519.840 0.000 1520.400 4.000 ;
    END
  END y[141]
  PIN y[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1523.200 0.000 1523.760 4.000 ;
    END
  END y[142]
  PIN y[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1526.560 0.000 1527.120 4.000 ;
    END
  END y[143]
  PIN y[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1529.920 0.000 1530.480 4.000 ;
    END
  END y[144]
  PIN y[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1533.280 0.000 1533.840 4.000 ;
    END
  END y[145]
  PIN y[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1536.640 0.000 1537.200 4.000 ;
    END
  END y[146]
  PIN y[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1540.000 0.000 1540.560 4.000 ;
    END
  END y[147]
  PIN y[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1543.360 0.000 1543.920 4.000 ;
    END
  END y[148]
  PIN y[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1546.720 0.000 1547.280 4.000 ;
    END
  END y[149]
  PIN y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1093.120 0.000 1093.680 4.000 ;
    END
  END y[14]
  PIN y[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1550.080 0.000 1550.640 4.000 ;
    END
  END y[150]
  PIN y[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1553.440 0.000 1554.000 4.000 ;
    END
  END y[151]
  PIN y[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1556.800 0.000 1557.360 4.000 ;
    END
  END y[152]
  PIN y[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1560.160 0.000 1560.720 4.000 ;
    END
  END y[153]
  PIN y[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1563.520 0.000 1564.080 4.000 ;
    END
  END y[154]
  PIN y[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1566.880 0.000 1567.440 4.000 ;
    END
  END y[155]
  PIN y[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1570.240 0.000 1570.800 4.000 ;
    END
  END y[156]
  PIN y[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1573.600 0.000 1574.160 4.000 ;
    END
  END y[157]
  PIN y[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1576.960 0.000 1577.520 4.000 ;
    END
  END y[158]
  PIN y[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1580.320 0.000 1580.880 4.000 ;
    END
  END y[159]
  PIN y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 0.000 1097.040 4.000 ;
    END
  END y[15]
  PIN y[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1583.680 0.000 1584.240 4.000 ;
    END
  END y[160]
  PIN y[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1587.040 0.000 1587.600 4.000 ;
    END
  END y[161]
  PIN y[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1590.400 0.000 1590.960 4.000 ;
    END
  END y[162]
  PIN y[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1593.760 0.000 1594.320 4.000 ;
    END
  END y[163]
  PIN y[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1597.120 0.000 1597.680 4.000 ;
    END
  END y[164]
  PIN y[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1600.480 0.000 1601.040 4.000 ;
    END
  END y[165]
  PIN y[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1603.840 0.000 1604.400 4.000 ;
    END
  END y[166]
  PIN y[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1607.200 0.000 1607.760 4.000 ;
    END
  END y[167]
  PIN y[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1610.560 0.000 1611.120 4.000 ;
    END
  END y[168]
  PIN y[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1613.920 0.000 1614.480 4.000 ;
    END
  END y[169]
  PIN y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1099.840 0.000 1100.400 4.000 ;
    END
  END y[16]
  PIN y[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1617.280 0.000 1617.840 4.000 ;
    END
  END y[170]
  PIN y[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1620.640 0.000 1621.200 4.000 ;
    END
  END y[171]
  PIN y[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1624.000 0.000 1624.560 4.000 ;
    END
  END y[172]
  PIN y[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1627.360 0.000 1627.920 4.000 ;
    END
  END y[173]
  PIN y[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1630.720 0.000 1631.280 4.000 ;
    END
  END y[174]
  PIN y[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1634.080 0.000 1634.640 4.000 ;
    END
  END y[175]
  PIN y[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1637.440 0.000 1638.000 4.000 ;
    END
  END y[176]
  PIN y[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1640.800 0.000 1641.360 4.000 ;
    END
  END y[177]
  PIN y[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1644.160 0.000 1644.720 4.000 ;
    END
  END y[178]
  PIN y[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1647.520 0.000 1648.080 4.000 ;
    END
  END y[179]
  PIN y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1103.200 0.000 1103.760 4.000 ;
    END
  END y[17]
  PIN y[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1650.880 0.000 1651.440 4.000 ;
    END
  END y[180]
  PIN y[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1654.240 0.000 1654.800 4.000 ;
    END
  END y[181]
  PIN y[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1657.600 0.000 1658.160 4.000 ;
    END
  END y[182]
  PIN y[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1660.960 0.000 1661.520 4.000 ;
    END
  END y[183]
  PIN y[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1664.320 0.000 1664.880 4.000 ;
    END
  END y[184]
  PIN y[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1667.680 0.000 1668.240 4.000 ;
    END
  END y[185]
  PIN y[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1671.040 0.000 1671.600 4.000 ;
    END
  END y[186]
  PIN y[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1674.400 0.000 1674.960 4.000 ;
    END
  END y[187]
  PIN y[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1677.760 0.000 1678.320 4.000 ;
    END
  END y[188]
  PIN y[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1681.120 0.000 1681.680 4.000 ;
    END
  END y[189]
  PIN y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1106.560 0.000 1107.120 4.000 ;
    END
  END y[18]
  PIN y[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1684.480 0.000 1685.040 4.000 ;
    END
  END y[190]
  PIN y[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1687.840 0.000 1688.400 4.000 ;
    END
  END y[191]
  PIN y[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1691.200 0.000 1691.760 4.000 ;
    END
  END y[192]
  PIN y[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1694.560 0.000 1695.120 4.000 ;
    END
  END y[193]
  PIN y[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1697.920 0.000 1698.480 4.000 ;
    END
  END y[194]
  PIN y[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1701.280 0.000 1701.840 4.000 ;
    END
  END y[195]
  PIN y[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1704.640 0.000 1705.200 4.000 ;
    END
  END y[196]
  PIN y[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1708.000 0.000 1708.560 4.000 ;
    END
  END y[197]
  PIN y[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1711.360 0.000 1711.920 4.000 ;
    END
  END y[198]
  PIN y[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1714.720 0.000 1715.280 4.000 ;
    END
  END y[199]
  PIN y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1109.920 0.000 1110.480 4.000 ;
    END
  END y[19]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1049.440 0.000 1050.000 4.000 ;
    END
  END y[1]
  PIN y[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1718.080 0.000 1718.640 4.000 ;
    END
  END y[200]
  PIN y[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1721.440 0.000 1722.000 4.000 ;
    END
  END y[201]
  PIN y[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1724.800 0.000 1725.360 4.000 ;
    END
  END y[202]
  PIN y[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1728.160 0.000 1728.720 4.000 ;
    END
  END y[203]
  PIN y[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1731.520 0.000 1732.080 4.000 ;
    END
  END y[204]
  PIN y[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1734.880 0.000 1735.440 4.000 ;
    END
  END y[205]
  PIN y[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1738.240 0.000 1738.800 4.000 ;
    END
  END y[206]
  PIN y[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1741.600 0.000 1742.160 4.000 ;
    END
  END y[207]
  PIN y[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1744.960 0.000 1745.520 4.000 ;
    END
  END y[208]
  PIN y[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1748.320 0.000 1748.880 4.000 ;
    END
  END y[209]
  PIN y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1113.280 0.000 1113.840 4.000 ;
    END
  END y[20]
  PIN y[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1751.680 0.000 1752.240 4.000 ;
    END
  END y[210]
  PIN y[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1755.040 0.000 1755.600 4.000 ;
    END
  END y[211]
  PIN y[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1758.400 0.000 1758.960 4.000 ;
    END
  END y[212]
  PIN y[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1761.760 0.000 1762.320 4.000 ;
    END
  END y[213]
  PIN y[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1765.120 0.000 1765.680 4.000 ;
    END
  END y[214]
  PIN y[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1768.480 0.000 1769.040 4.000 ;
    END
  END y[215]
  PIN y[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1771.840 0.000 1772.400 4.000 ;
    END
  END y[216]
  PIN y[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1775.200 0.000 1775.760 4.000 ;
    END
  END y[217]
  PIN y[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1778.560 0.000 1779.120 4.000 ;
    END
  END y[218]
  PIN y[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1781.920 0.000 1782.480 4.000 ;
    END
  END y[219]
  PIN y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1116.640 0.000 1117.200 4.000 ;
    END
  END y[21]
  PIN y[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1785.280 0.000 1785.840 4.000 ;
    END
  END y[220]
  PIN y[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1788.640 0.000 1789.200 4.000 ;
    END
  END y[221]
  PIN y[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1792.000 0.000 1792.560 4.000 ;
    END
  END y[222]
  PIN y[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1795.360 0.000 1795.920 4.000 ;
    END
  END y[223]
  PIN y[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1798.720 0.000 1799.280 4.000 ;
    END
  END y[224]
  PIN y[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1802.080 0.000 1802.640 4.000 ;
    END
  END y[225]
  PIN y[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1805.440 0.000 1806.000 4.000 ;
    END
  END y[226]
  PIN y[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1808.800 0.000 1809.360 4.000 ;
    END
  END y[227]
  PIN y[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1812.160 0.000 1812.720 4.000 ;
    END
  END y[228]
  PIN y[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1815.520 0.000 1816.080 4.000 ;
    END
  END y[229]
  PIN y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1120.000 0.000 1120.560 4.000 ;
    END
  END y[22]
  PIN y[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1818.880 0.000 1819.440 4.000 ;
    END
  END y[230]
  PIN y[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1822.240 0.000 1822.800 4.000 ;
    END
  END y[231]
  PIN y[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1825.600 0.000 1826.160 4.000 ;
    END
  END y[232]
  PIN y[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1828.960 0.000 1829.520 4.000 ;
    END
  END y[233]
  PIN y[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1832.320 0.000 1832.880 4.000 ;
    END
  END y[234]
  PIN y[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1835.680 0.000 1836.240 4.000 ;
    END
  END y[235]
  PIN y[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1839.040 0.000 1839.600 4.000 ;
    END
  END y[236]
  PIN y[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1842.400 0.000 1842.960 4.000 ;
    END
  END y[237]
  PIN y[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1845.760 0.000 1846.320 4.000 ;
    END
  END y[238]
  PIN y[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1849.120 0.000 1849.680 4.000 ;
    END
  END y[239]
  PIN y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1123.360 0.000 1123.920 4.000 ;
    END
  END y[23]
  PIN y[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1852.480 0.000 1853.040 4.000 ;
    END
  END y[240]
  PIN y[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1855.840 0.000 1856.400 4.000 ;
    END
  END y[241]
  PIN y[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1859.200 0.000 1859.760 4.000 ;
    END
  END y[242]
  PIN y[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1862.560 0.000 1863.120 4.000 ;
    END
  END y[243]
  PIN y[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1865.920 0.000 1866.480 4.000 ;
    END
  END y[244]
  PIN y[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1869.280 0.000 1869.840 4.000 ;
    END
  END y[245]
  PIN y[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1872.640 0.000 1873.200 4.000 ;
    END
  END y[246]
  PIN y[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1876.000 0.000 1876.560 4.000 ;
    END
  END y[247]
  PIN y[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1879.360 0.000 1879.920 4.000 ;
    END
  END y[248]
  PIN y[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1882.720 0.000 1883.280 4.000 ;
    END
  END y[249]
  PIN y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1126.720 0.000 1127.280 4.000 ;
    END
  END y[24]
  PIN y[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1886.080 0.000 1886.640 4.000 ;
    END
  END y[250]
  PIN y[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1889.440 0.000 1890.000 4.000 ;
    END
  END y[251]
  PIN y[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1892.800 0.000 1893.360 4.000 ;
    END
  END y[252]
  PIN y[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1896.160 0.000 1896.720 4.000 ;
    END
  END y[253]
  PIN y[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1899.520 0.000 1900.080 4.000 ;
    END
  END y[254]
  PIN y[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1902.880 0.000 1903.440 4.000 ;
    END
  END y[255]
  PIN y[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1906.240 0.000 1906.800 4.000 ;
    END
  END y[256]
  PIN y[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1909.600 0.000 1910.160 4.000 ;
    END
  END y[257]
  PIN y[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1912.960 0.000 1913.520 4.000 ;
    END
  END y[258]
  PIN y[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1916.320 0.000 1916.880 4.000 ;
    END
  END y[259]
  PIN y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1130.080 0.000 1130.640 4.000 ;
    END
  END y[25]
  PIN y[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1919.680 0.000 1920.240 4.000 ;
    END
  END y[260]
  PIN y[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1923.040 0.000 1923.600 4.000 ;
    END
  END y[261]
  PIN y[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1926.400 0.000 1926.960 4.000 ;
    END
  END y[262]
  PIN y[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1929.760 0.000 1930.320 4.000 ;
    END
  END y[263]
  PIN y[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1933.120 0.000 1933.680 4.000 ;
    END
  END y[264]
  PIN y[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1936.480 0.000 1937.040 4.000 ;
    END
  END y[265]
  PIN y[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1939.840 0.000 1940.400 4.000 ;
    END
  END y[266]
  PIN y[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1943.200 0.000 1943.760 4.000 ;
    END
  END y[267]
  PIN y[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1946.560 0.000 1947.120 4.000 ;
    END
  END y[268]
  PIN y[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1949.920 0.000 1950.480 4.000 ;
    END
  END y[269]
  PIN y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1133.440 0.000 1134.000 4.000 ;
    END
  END y[26]
  PIN y[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1953.280 0.000 1953.840 4.000 ;
    END
  END y[270]
  PIN y[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1956.640 0.000 1957.200 4.000 ;
    END
  END y[271]
  PIN y[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1960.000 0.000 1960.560 4.000 ;
    END
  END y[272]
  PIN y[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1963.360 0.000 1963.920 4.000 ;
    END
  END y[273]
  PIN y[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1966.720 0.000 1967.280 4.000 ;
    END
  END y[274]
  PIN y[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1970.080 0.000 1970.640 4.000 ;
    END
  END y[275]
  PIN y[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1973.440 0.000 1974.000 4.000 ;
    END
  END y[276]
  PIN y[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1976.800 0.000 1977.360 4.000 ;
    END
  END y[277]
  PIN y[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1980.160 0.000 1980.720 4.000 ;
    END
  END y[278]
  PIN y[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1983.520 0.000 1984.080 4.000 ;
    END
  END y[279]
  PIN y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1136.800 0.000 1137.360 4.000 ;
    END
  END y[27]
  PIN y[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1986.880 0.000 1987.440 4.000 ;
    END
  END y[280]
  PIN y[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1990.240 0.000 1990.800 4.000 ;
    END
  END y[281]
  PIN y[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1993.600 0.000 1994.160 4.000 ;
    END
  END y[282]
  PIN y[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1996.960 0.000 1997.520 4.000 ;
    END
  END y[283]
  PIN y[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2000.320 0.000 2000.880 4.000 ;
    END
  END y[284]
  PIN y[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2003.680 0.000 2004.240 4.000 ;
    END
  END y[285]
  PIN y[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2007.040 0.000 2007.600 4.000 ;
    END
  END y[286]
  PIN y[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2010.400 0.000 2010.960 4.000 ;
    END
  END y[287]
  PIN y[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2013.760 0.000 2014.320 4.000 ;
    END
  END y[288]
  PIN y[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2017.120 0.000 2017.680 4.000 ;
    END
  END y[289]
  PIN y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1140.160 0.000 1140.720 4.000 ;
    END
  END y[28]
  PIN y[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2020.480 0.000 2021.040 4.000 ;
    END
  END y[290]
  PIN y[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2023.840 0.000 2024.400 4.000 ;
    END
  END y[291]
  PIN y[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2027.200 0.000 2027.760 4.000 ;
    END
  END y[292]
  PIN y[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2030.560 0.000 2031.120 4.000 ;
    END
  END y[293]
  PIN y[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2033.920 0.000 2034.480 4.000 ;
    END
  END y[294]
  PIN y[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2037.280 0.000 2037.840 4.000 ;
    END
  END y[295]
  PIN y[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2040.640 0.000 2041.200 4.000 ;
    END
  END y[296]
  PIN y[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2044.000 0.000 2044.560 4.000 ;
    END
  END y[297]
  PIN y[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2047.360 0.000 2047.920 4.000 ;
    END
  END y[298]
  PIN y[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2050.720 0.000 2051.280 4.000 ;
    END
  END y[299]
  PIN y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1143.520 0.000 1144.080 4.000 ;
    END
  END y[29]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1052.800 0.000 1053.360 4.000 ;
    END
  END y[2]
  PIN y[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2054.080 0.000 2054.640 4.000 ;
    END
  END y[300]
  PIN y[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2057.440 0.000 2058.000 4.000 ;
    END
  END y[301]
  PIN y[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2060.800 0.000 2061.360 4.000 ;
    END
  END y[302]
  PIN y[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2064.160 0.000 2064.720 4.000 ;
    END
  END y[303]
  PIN y[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2067.520 0.000 2068.080 4.000 ;
    END
  END y[304]
  PIN y[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2070.880 0.000 2071.440 4.000 ;
    END
  END y[305]
  PIN y[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2074.240 0.000 2074.800 4.000 ;
    END
  END y[306]
  PIN y[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2077.600 0.000 2078.160 4.000 ;
    END
  END y[307]
  PIN y[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2080.960 0.000 2081.520 4.000 ;
    END
  END y[308]
  PIN y[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2084.320 0.000 2084.880 4.000 ;
    END
  END y[309]
  PIN y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1146.880 0.000 1147.440 4.000 ;
    END
  END y[30]
  PIN y[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2087.680 0.000 2088.240 4.000 ;
    END
  END y[310]
  PIN y[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2091.040 0.000 2091.600 4.000 ;
    END
  END y[311]
  PIN y[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2094.400 0.000 2094.960 4.000 ;
    END
  END y[312]
  PIN y[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2097.760 0.000 2098.320 4.000 ;
    END
  END y[313]
  PIN y[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2101.120 0.000 2101.680 4.000 ;
    END
  END y[314]
  PIN y[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2104.480 0.000 2105.040 4.000 ;
    END
  END y[315]
  PIN y[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2107.840 0.000 2108.400 4.000 ;
    END
  END y[316]
  PIN y[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2111.200 0.000 2111.760 4.000 ;
    END
  END y[317]
  PIN y[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2114.560 0.000 2115.120 4.000 ;
    END
  END y[318]
  PIN y[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2117.920 0.000 2118.480 4.000 ;
    END
  END y[319]
  PIN y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1150.240 0.000 1150.800 4.000 ;
    END
  END y[31]
  PIN y[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2121.280 0.000 2121.840 4.000 ;
    END
  END y[320]
  PIN y[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2124.640 0.000 2125.200 4.000 ;
    END
  END y[321]
  PIN y[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2128.000 0.000 2128.560 4.000 ;
    END
  END y[322]
  PIN y[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2131.360 0.000 2131.920 4.000 ;
    END
  END y[323]
  PIN y[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2134.720 0.000 2135.280 4.000 ;
    END
  END y[324]
  PIN y[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2138.080 0.000 2138.640 4.000 ;
    END
  END y[325]
  PIN y[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2141.440 0.000 2142.000 4.000 ;
    END
  END y[326]
  PIN y[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2144.800 0.000 2145.360 4.000 ;
    END
  END y[327]
  PIN y[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2148.160 0.000 2148.720 4.000 ;
    END
  END y[328]
  PIN y[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2151.520 0.000 2152.080 4.000 ;
    END
  END y[329]
  PIN y[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1153.600 0.000 1154.160 4.000 ;
    END
  END y[32]
  PIN y[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2154.880 0.000 2155.440 4.000 ;
    END
  END y[330]
  PIN y[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2158.240 0.000 2158.800 4.000 ;
    END
  END y[331]
  PIN y[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2161.600 0.000 2162.160 4.000 ;
    END
  END y[332]
  PIN y[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2164.960 0.000 2165.520 4.000 ;
    END
  END y[333]
  PIN y[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2168.320 0.000 2168.880 4.000 ;
    END
  END y[334]
  PIN y[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2171.680 0.000 2172.240 4.000 ;
    END
  END y[335]
  PIN y[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2175.040 0.000 2175.600 4.000 ;
    END
  END y[336]
  PIN y[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2178.400 0.000 2178.960 4.000 ;
    END
  END y[337]
  PIN y[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2181.760 0.000 2182.320 4.000 ;
    END
  END y[338]
  PIN y[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2185.120 0.000 2185.680 4.000 ;
    END
  END y[339]
  PIN y[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1156.960 0.000 1157.520 4.000 ;
    END
  END y[33]
  PIN y[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2188.480 0.000 2189.040 4.000 ;
    END
  END y[340]
  PIN y[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2191.840 0.000 2192.400 4.000 ;
    END
  END y[341]
  PIN y[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2195.200 0.000 2195.760 4.000 ;
    END
  END y[342]
  PIN y[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2198.560 0.000 2199.120 4.000 ;
    END
  END y[343]
  PIN y[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2201.920 0.000 2202.480 4.000 ;
    END
  END y[344]
  PIN y[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2205.280 0.000 2205.840 4.000 ;
    END
  END y[345]
  PIN y[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2208.640 0.000 2209.200 4.000 ;
    END
  END y[346]
  PIN y[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2212.000 0.000 2212.560 4.000 ;
    END
  END y[347]
  PIN y[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2215.360 0.000 2215.920 4.000 ;
    END
  END y[348]
  PIN y[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2218.720 0.000 2219.280 4.000 ;
    END
  END y[349]
  PIN y[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1160.320 0.000 1160.880 4.000 ;
    END
  END y[34]
  PIN y[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2222.080 0.000 2222.640 4.000 ;
    END
  END y[350]
  PIN y[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2225.440 0.000 2226.000 4.000 ;
    END
  END y[351]
  PIN y[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2228.800 0.000 2229.360 4.000 ;
    END
  END y[352]
  PIN y[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2232.160 0.000 2232.720 4.000 ;
    END
  END y[353]
  PIN y[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2235.520 0.000 2236.080 4.000 ;
    END
  END y[354]
  PIN y[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2238.880 0.000 2239.440 4.000 ;
    END
  END y[355]
  PIN y[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2242.240 0.000 2242.800 4.000 ;
    END
  END y[356]
  PIN y[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2245.600 0.000 2246.160 4.000 ;
    END
  END y[357]
  PIN y[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2248.960 0.000 2249.520 4.000 ;
    END
  END y[358]
  PIN y[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2252.320 0.000 2252.880 4.000 ;
    END
  END y[359]
  PIN y[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1163.680 0.000 1164.240 4.000 ;
    END
  END y[35]
  PIN y[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2255.680 0.000 2256.240 4.000 ;
    END
  END y[360]
  PIN y[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2259.040 0.000 2259.600 4.000 ;
    END
  END y[361]
  PIN y[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2262.400 0.000 2262.960 4.000 ;
    END
  END y[362]
  PIN y[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2265.760 0.000 2266.320 4.000 ;
    END
  END y[363]
  PIN y[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2269.120 0.000 2269.680 4.000 ;
    END
  END y[364]
  PIN y[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2272.480 0.000 2273.040 4.000 ;
    END
  END y[365]
  PIN y[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2275.840 0.000 2276.400 4.000 ;
    END
  END y[366]
  PIN y[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2279.200 0.000 2279.760 4.000 ;
    END
  END y[367]
  PIN y[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2282.560 0.000 2283.120 4.000 ;
    END
  END y[368]
  PIN y[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2285.920 0.000 2286.480 4.000 ;
    END
  END y[369]
  PIN y[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1167.040 0.000 1167.600 4.000 ;
    END
  END y[36]
  PIN y[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2289.280 0.000 2289.840 4.000 ;
    END
  END y[370]
  PIN y[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2292.640 0.000 2293.200 4.000 ;
    END
  END y[371]
  PIN y[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2296.000 0.000 2296.560 4.000 ;
    END
  END y[372]
  PIN y[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2299.360 0.000 2299.920 4.000 ;
    END
  END y[373]
  PIN y[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2302.720 0.000 2303.280 4.000 ;
    END
  END y[374]
  PIN y[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2306.080 0.000 2306.640 4.000 ;
    END
  END y[375]
  PIN y[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2309.440 0.000 2310.000 4.000 ;
    END
  END y[376]
  PIN y[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2312.800 0.000 2313.360 4.000 ;
    END
  END y[377]
  PIN y[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2316.160 0.000 2316.720 4.000 ;
    END
  END y[378]
  PIN y[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2319.520 0.000 2320.080 4.000 ;
    END
  END y[379]
  PIN y[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1170.400 0.000 1170.960 4.000 ;
    END
  END y[37]
  PIN y[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2322.880 0.000 2323.440 4.000 ;
    END
  END y[380]
  PIN y[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2326.240 0.000 2326.800 4.000 ;
    END
  END y[381]
  PIN y[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2329.600 0.000 2330.160 4.000 ;
    END
  END y[382]
  PIN y[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2332.960 0.000 2333.520 4.000 ;
    END
  END y[383]
  PIN y[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2336.320 0.000 2336.880 4.000 ;
    END
  END y[384]
  PIN y[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2339.680 0.000 2340.240 4.000 ;
    END
  END y[385]
  PIN y[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2343.040 0.000 2343.600 4.000 ;
    END
  END y[386]
  PIN y[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2346.400 0.000 2346.960 4.000 ;
    END
  END y[387]
  PIN y[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2349.760 0.000 2350.320 4.000 ;
    END
  END y[388]
  PIN y[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2353.120 0.000 2353.680 4.000 ;
    END
  END y[389]
  PIN y[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1173.760 0.000 1174.320 4.000 ;
    END
  END y[38]
  PIN y[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2356.480 0.000 2357.040 4.000 ;
    END
  END y[390]
  PIN y[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2359.840 0.000 2360.400 4.000 ;
    END
  END y[391]
  PIN y[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2363.200 0.000 2363.760 4.000 ;
    END
  END y[392]
  PIN y[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2366.560 0.000 2367.120 4.000 ;
    END
  END y[393]
  PIN y[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2369.920 0.000 2370.480 4.000 ;
    END
  END y[394]
  PIN y[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2373.280 0.000 2373.840 4.000 ;
    END
  END y[395]
  PIN y[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2376.640 0.000 2377.200 4.000 ;
    END
  END y[396]
  PIN y[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2380.000 0.000 2380.560 4.000 ;
    END
  END y[397]
  PIN y[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2383.360 0.000 2383.920 4.000 ;
    END
  END y[398]
  PIN y[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2386.720 0.000 2387.280 4.000 ;
    END
  END y[399]
  PIN y[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1177.120 0.000 1177.680 4.000 ;
    END
  END y[39]
  PIN y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.160 0.000 1056.720 4.000 ;
    END
  END y[3]
  PIN y[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2390.080 0.000 2390.640 4.000 ;
    END
  END y[400]
  PIN y[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2393.440 0.000 2394.000 4.000 ;
    END
  END y[401]
  PIN y[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2396.800 0.000 2397.360 4.000 ;
    END
  END y[402]
  PIN y[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2400.160 0.000 2400.720 4.000 ;
    END
  END y[403]
  PIN y[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2403.520 0.000 2404.080 4.000 ;
    END
  END y[404]
  PIN y[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2406.880 0.000 2407.440 4.000 ;
    END
  END y[405]
  PIN y[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2410.240 0.000 2410.800 4.000 ;
    END
  END y[406]
  PIN y[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2413.600 0.000 2414.160 4.000 ;
    END
  END y[407]
  PIN y[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2416.960 0.000 2417.520 4.000 ;
    END
  END y[408]
  PIN y[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2420.320 0.000 2420.880 4.000 ;
    END
  END y[409]
  PIN y[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1180.480 0.000 1181.040 4.000 ;
    END
  END y[40]
  PIN y[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2423.680 0.000 2424.240 4.000 ;
    END
  END y[410]
  PIN y[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2427.040 0.000 2427.600 4.000 ;
    END
  END y[411]
  PIN y[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2430.400 0.000 2430.960 4.000 ;
    END
  END y[412]
  PIN y[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2433.760 0.000 2434.320 4.000 ;
    END
  END y[413]
  PIN y[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2437.120 0.000 2437.680 4.000 ;
    END
  END y[414]
  PIN y[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2440.480 0.000 2441.040 4.000 ;
    END
  END y[415]
  PIN y[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2443.840 0.000 2444.400 4.000 ;
    END
  END y[416]
  PIN y[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2447.200 0.000 2447.760 4.000 ;
    END
  END y[417]
  PIN y[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2450.560 0.000 2451.120 4.000 ;
    END
  END y[418]
  PIN y[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2453.920 0.000 2454.480 4.000 ;
    END
  END y[419]
  PIN y[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1183.840 0.000 1184.400 4.000 ;
    END
  END y[41]
  PIN y[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2457.280 0.000 2457.840 4.000 ;
    END
  END y[420]
  PIN y[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2460.640 0.000 2461.200 4.000 ;
    END
  END y[421]
  PIN y[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2464.000 0.000 2464.560 4.000 ;
    END
  END y[422]
  PIN y[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2467.360 0.000 2467.920 4.000 ;
    END
  END y[423]
  PIN y[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2470.720 0.000 2471.280 4.000 ;
    END
  END y[424]
  PIN y[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2474.080 0.000 2474.640 4.000 ;
    END
  END y[425]
  PIN y[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2477.440 0.000 2478.000 4.000 ;
    END
  END y[426]
  PIN y[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2480.800 0.000 2481.360 4.000 ;
    END
  END y[427]
  PIN y[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2484.160 0.000 2484.720 4.000 ;
    END
  END y[428]
  PIN y[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2487.520 0.000 2488.080 4.000 ;
    END
  END y[429]
  PIN y[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1187.200 0.000 1187.760 4.000 ;
    END
  END y[42]
  PIN y[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2490.880 0.000 2491.440 4.000 ;
    END
  END y[430]
  PIN y[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2494.240 0.000 2494.800 4.000 ;
    END
  END y[431]
  PIN y[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2497.600 0.000 2498.160 4.000 ;
    END
  END y[432]
  PIN y[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2500.960 0.000 2501.520 4.000 ;
    END
  END y[433]
  PIN y[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2504.320 0.000 2504.880 4.000 ;
    END
  END y[434]
  PIN y[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2507.680 0.000 2508.240 4.000 ;
    END
  END y[435]
  PIN y[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2511.040 0.000 2511.600 4.000 ;
    END
  END y[436]
  PIN y[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2514.400 0.000 2514.960 4.000 ;
    END
  END y[437]
  PIN y[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2517.760 0.000 2518.320 4.000 ;
    END
  END y[438]
  PIN y[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2521.120 0.000 2521.680 4.000 ;
    END
  END y[439]
  PIN y[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1190.560 0.000 1191.120 4.000 ;
    END
  END y[43]
  PIN y[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2524.480 0.000 2525.040 4.000 ;
    END
  END y[440]
  PIN y[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2527.840 0.000 2528.400 4.000 ;
    END
  END y[441]
  PIN y[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2531.200 0.000 2531.760 4.000 ;
    END
  END y[442]
  PIN y[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2534.560 0.000 2535.120 4.000 ;
    END
  END y[443]
  PIN y[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2537.920 0.000 2538.480 4.000 ;
    END
  END y[444]
  PIN y[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2541.280 0.000 2541.840 4.000 ;
    END
  END y[445]
  PIN y[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2544.640 0.000 2545.200 4.000 ;
    END
  END y[446]
  PIN y[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2548.000 0.000 2548.560 4.000 ;
    END
  END y[447]
  PIN y[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2551.360 0.000 2551.920 4.000 ;
    END
  END y[448]
  PIN y[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2554.720 0.000 2555.280 4.000 ;
    END
  END y[449]
  PIN y[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1193.920 0.000 1194.480 4.000 ;
    END
  END y[44]
  PIN y[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2558.080 0.000 2558.640 4.000 ;
    END
  END y[450]
  PIN y[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2561.440 0.000 2562.000 4.000 ;
    END
  END y[451]
  PIN y[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2564.800 0.000 2565.360 4.000 ;
    END
  END y[452]
  PIN y[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2568.160 0.000 2568.720 4.000 ;
    END
  END y[453]
  PIN y[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2571.520 0.000 2572.080 4.000 ;
    END
  END y[454]
  PIN y[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2574.880 0.000 2575.440 4.000 ;
    END
  END y[455]
  PIN y[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2578.240 0.000 2578.800 4.000 ;
    END
  END y[456]
  PIN y[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2581.600 0.000 2582.160 4.000 ;
    END
  END y[457]
  PIN y[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2584.960 0.000 2585.520 4.000 ;
    END
  END y[458]
  PIN y[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2588.320 0.000 2588.880 4.000 ;
    END
  END y[459]
  PIN y[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1197.280 0.000 1197.840 4.000 ;
    END
  END y[45]
  PIN y[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2591.680 0.000 2592.240 4.000 ;
    END
  END y[460]
  PIN y[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2595.040 0.000 2595.600 4.000 ;
    END
  END y[461]
  PIN y[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2598.400 0.000 2598.960 4.000 ;
    END
  END y[462]
  PIN y[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2601.760 0.000 2602.320 4.000 ;
    END
  END y[463]
  PIN y[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2605.120 0.000 2605.680 4.000 ;
    END
  END y[464]
  PIN y[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2608.480 0.000 2609.040 4.000 ;
    END
  END y[465]
  PIN y[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2611.840 0.000 2612.400 4.000 ;
    END
  END y[466]
  PIN y[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2615.200 0.000 2615.760 4.000 ;
    END
  END y[467]
  PIN y[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2618.560 0.000 2619.120 4.000 ;
    END
  END y[468]
  PIN y[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2621.920 0.000 2622.480 4.000 ;
    END
  END y[469]
  PIN y[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1200.640 0.000 1201.200 4.000 ;
    END
  END y[46]
  PIN y[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2625.280 0.000 2625.840 4.000 ;
    END
  END y[470]
  PIN y[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2628.640 0.000 2629.200 4.000 ;
    END
  END y[471]
  PIN y[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2632.000 0.000 2632.560 4.000 ;
    END
  END y[472]
  PIN y[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2635.360 0.000 2635.920 4.000 ;
    END
  END y[473]
  PIN y[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2638.720 0.000 2639.280 4.000 ;
    END
  END y[474]
  PIN y[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2642.080 0.000 2642.640 4.000 ;
    END
  END y[475]
  PIN y[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2645.440 0.000 2646.000 4.000 ;
    END
  END y[476]
  PIN y[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2648.800 0.000 2649.360 4.000 ;
    END
  END y[477]
  PIN y[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2652.160 0.000 2652.720 4.000 ;
    END
  END y[478]
  PIN y[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2655.520 0.000 2656.080 4.000 ;
    END
  END y[479]
  PIN y[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1204.000 0.000 1204.560 4.000 ;
    END
  END y[47]
  PIN y[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2658.880 0.000 2659.440 4.000 ;
    END
  END y[480]
  PIN y[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2662.240 0.000 2662.800 4.000 ;
    END
  END y[481]
  PIN y[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2665.600 0.000 2666.160 4.000 ;
    END
  END y[482]
  PIN y[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2668.960 0.000 2669.520 4.000 ;
    END
  END y[483]
  PIN y[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2672.320 0.000 2672.880 4.000 ;
    END
  END y[484]
  PIN y[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2675.680 0.000 2676.240 4.000 ;
    END
  END y[485]
  PIN y[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2679.040 0.000 2679.600 4.000 ;
    END
  END y[486]
  PIN y[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2682.400 0.000 2682.960 4.000 ;
    END
  END y[487]
  PIN y[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2685.760 0.000 2686.320 4.000 ;
    END
  END y[488]
  PIN y[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2689.120 0.000 2689.680 4.000 ;
    END
  END y[489]
  PIN y[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1207.360 0.000 1207.920 4.000 ;
    END
  END y[48]
  PIN y[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2692.480 0.000 2693.040 4.000 ;
    END
  END y[490]
  PIN y[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2695.840 0.000 2696.400 4.000 ;
    END
  END y[491]
  PIN y[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2699.200 0.000 2699.760 4.000 ;
    END
  END y[492]
  PIN y[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2702.560 0.000 2703.120 4.000 ;
    END
  END y[493]
  PIN y[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2705.920 0.000 2706.480 4.000 ;
    END
  END y[494]
  PIN y[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2709.280 0.000 2709.840 4.000 ;
    END
  END y[495]
  PIN y[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2712.640 0.000 2713.200 4.000 ;
    END
  END y[496]
  PIN y[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2716.000 0.000 2716.560 4.000 ;
    END
  END y[497]
  PIN y[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2719.360 0.000 2719.920 4.000 ;
    END
  END y[498]
  PIN y[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2722.720 0.000 2723.280 4.000 ;
    END
  END y[499]
  PIN y[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1210.720 0.000 1211.280 4.000 ;
    END
  END y[49]
  PIN y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1059.520 0.000 1060.080 4.000 ;
    END
  END y[4]
  PIN y[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2726.080 0.000 2726.640 4.000 ;
    END
  END y[500]
  PIN y[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2729.440 0.000 2730.000 4.000 ;
    END
  END y[501]
  PIN y[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2732.800 0.000 2733.360 4.000 ;
    END
  END y[502]
  PIN y[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2736.160 0.000 2736.720 4.000 ;
    END
  END y[503]
  PIN y[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2739.520 0.000 2740.080 4.000 ;
    END
  END y[504]
  PIN y[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2742.880 0.000 2743.440 4.000 ;
    END
  END y[505]
  PIN y[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2746.240 0.000 2746.800 4.000 ;
    END
  END y[506]
  PIN y[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2749.600 0.000 2750.160 4.000 ;
    END
  END y[507]
  PIN y[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2752.960 0.000 2753.520 4.000 ;
    END
  END y[508]
  PIN y[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2756.320 0.000 2756.880 4.000 ;
    END
  END y[509]
  PIN y[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1214.080 0.000 1214.640 4.000 ;
    END
  END y[50]
  PIN y[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2759.680 0.000 2760.240 4.000 ;
    END
  END y[510]
  PIN y[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2763.040 0.000 2763.600 4.000 ;
    END
  END y[511]
  PIN y[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1217.440 0.000 1218.000 4.000 ;
    END
  END y[51]
  PIN y[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1220.800 0.000 1221.360 4.000 ;
    END
  END y[52]
  PIN y[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1224.160 0.000 1224.720 4.000 ;
    END
  END y[53]
  PIN y[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1227.520 0.000 1228.080 4.000 ;
    END
  END y[54]
  PIN y[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1230.880 0.000 1231.440 4.000 ;
    END
  END y[55]
  PIN y[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1234.240 0.000 1234.800 4.000 ;
    END
  END y[56]
  PIN y[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1237.600 0.000 1238.160 4.000 ;
    END
  END y[57]
  PIN y[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1240.960 0.000 1241.520 4.000 ;
    END
  END y[58]
  PIN y[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1244.320 0.000 1244.880 4.000 ;
    END
  END y[59]
  PIN y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1062.880 0.000 1063.440 4.000 ;
    END
  END y[5]
  PIN y[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1247.680 0.000 1248.240 4.000 ;
    END
  END y[60]
  PIN y[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1251.040 0.000 1251.600 4.000 ;
    END
  END y[61]
  PIN y[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1254.400 0.000 1254.960 4.000 ;
    END
  END y[62]
  PIN y[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1257.760 0.000 1258.320 4.000 ;
    END
  END y[63]
  PIN y[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1261.120 0.000 1261.680 4.000 ;
    END
  END y[64]
  PIN y[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1264.480 0.000 1265.040 4.000 ;
    END
  END y[65]
  PIN y[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1267.840 0.000 1268.400 4.000 ;
    END
  END y[66]
  PIN y[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1271.200 0.000 1271.760 4.000 ;
    END
  END y[67]
  PIN y[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1274.560 0.000 1275.120 4.000 ;
    END
  END y[68]
  PIN y[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1277.920 0.000 1278.480 4.000 ;
    END
  END y[69]
  PIN y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1066.240 0.000 1066.800 4.000 ;
    END
  END y[6]
  PIN y[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1281.280 0.000 1281.840 4.000 ;
    END
  END y[70]
  PIN y[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1284.640 0.000 1285.200 4.000 ;
    END
  END y[71]
  PIN y[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1288.000 0.000 1288.560 4.000 ;
    END
  END y[72]
  PIN y[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1291.360 0.000 1291.920 4.000 ;
    END
  END y[73]
  PIN y[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1294.720 0.000 1295.280 4.000 ;
    END
  END y[74]
  PIN y[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1298.080 0.000 1298.640 4.000 ;
    END
  END y[75]
  PIN y[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1301.440 0.000 1302.000 4.000 ;
    END
  END y[76]
  PIN y[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1304.800 0.000 1305.360 4.000 ;
    END
  END y[77]
  PIN y[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1308.160 0.000 1308.720 4.000 ;
    END
  END y[78]
  PIN y[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1311.520 0.000 1312.080 4.000 ;
    END
  END y[79]
  PIN y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1069.600 0.000 1070.160 4.000 ;
    END
  END y[7]
  PIN y[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1314.880 0.000 1315.440 4.000 ;
    END
  END y[80]
  PIN y[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1318.240 0.000 1318.800 4.000 ;
    END
  END y[81]
  PIN y[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1321.600 0.000 1322.160 4.000 ;
    END
  END y[82]
  PIN y[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1324.960 0.000 1325.520 4.000 ;
    END
  END y[83]
  PIN y[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1328.320 0.000 1328.880 4.000 ;
    END
  END y[84]
  PIN y[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1331.680 0.000 1332.240 4.000 ;
    END
  END y[85]
  PIN y[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1335.040 0.000 1335.600 4.000 ;
    END
  END y[86]
  PIN y[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1338.400 0.000 1338.960 4.000 ;
    END
  END y[87]
  PIN y[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1341.760 0.000 1342.320 4.000 ;
    END
  END y[88]
  PIN y[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1345.120 0.000 1345.680 4.000 ;
    END
  END y[89]
  PIN y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1072.960 0.000 1073.520 4.000 ;
    END
  END y[8]
  PIN y[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1348.480 0.000 1349.040 4.000 ;
    END
  END y[90]
  PIN y[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1351.840 0.000 1352.400 4.000 ;
    END
  END y[91]
  PIN y[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1355.200 0.000 1355.760 4.000 ;
    END
  END y[92]
  PIN y[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1358.560 0.000 1359.120 4.000 ;
    END
  END y[93]
  PIN y[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1361.920 0.000 1362.480 4.000 ;
    END
  END y[94]
  PIN y[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1365.280 0.000 1365.840 4.000 ;
    END
  END y[95]
  PIN y[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1368.640 0.000 1369.200 4.000 ;
    END
  END y[96]
  PIN y[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1372.000 0.000 1372.560 4.000 ;
    END
  END y[97]
  PIN y[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1375.360 0.000 1375.920 4.000 ;
    END
  END y[98]
  PIN y[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1378.720 0.000 1379.280 4.000 ;
    END
  END y[99]
  PIN y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1076.320 0.000 1076.880 4.000 ;
    END
  END y[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 2793.280 788.890 ;
      LAYER Metal2 ;
        RECT 7.980 795.700 36.660 796.000 ;
        RECT 37.820 795.700 57.940 796.000 ;
        RECT 59.100 795.700 79.220 796.000 ;
        RECT 80.380 795.700 100.500 796.000 ;
        RECT 101.660 795.700 121.780 796.000 ;
        RECT 122.940 795.700 143.060 796.000 ;
        RECT 144.220 795.700 164.340 796.000 ;
        RECT 165.500 795.700 185.620 796.000 ;
        RECT 186.780 795.700 206.900 796.000 ;
        RECT 208.060 795.700 228.180 796.000 ;
        RECT 229.340 795.700 249.460 796.000 ;
        RECT 250.620 795.700 270.740 796.000 ;
        RECT 271.900 795.700 292.020 796.000 ;
        RECT 293.180 795.700 313.300 796.000 ;
        RECT 314.460 795.700 334.580 796.000 ;
        RECT 335.740 795.700 355.860 796.000 ;
        RECT 357.020 795.700 377.140 796.000 ;
        RECT 378.300 795.700 398.420 796.000 ;
        RECT 399.580 795.700 419.700 796.000 ;
        RECT 420.860 795.700 440.980 796.000 ;
        RECT 442.140 795.700 462.260 796.000 ;
        RECT 463.420 795.700 483.540 796.000 ;
        RECT 484.700 795.700 504.820 796.000 ;
        RECT 505.980 795.700 526.100 796.000 ;
        RECT 527.260 795.700 547.380 796.000 ;
        RECT 548.540 795.700 568.660 796.000 ;
        RECT 569.820 795.700 589.940 796.000 ;
        RECT 591.100 795.700 611.220 796.000 ;
        RECT 612.380 795.700 632.500 796.000 ;
        RECT 633.660 795.700 653.780 796.000 ;
        RECT 654.940 795.700 675.060 796.000 ;
        RECT 676.220 795.700 696.340 796.000 ;
        RECT 697.500 795.700 717.620 796.000 ;
        RECT 718.780 795.700 738.900 796.000 ;
        RECT 740.060 795.700 760.180 796.000 ;
        RECT 761.340 795.700 781.460 796.000 ;
        RECT 782.620 795.700 802.740 796.000 ;
        RECT 803.900 795.700 824.020 796.000 ;
        RECT 825.180 795.700 845.300 796.000 ;
        RECT 846.460 795.700 866.580 796.000 ;
        RECT 867.740 795.700 887.860 796.000 ;
        RECT 889.020 795.700 909.140 796.000 ;
        RECT 910.300 795.700 930.420 796.000 ;
        RECT 931.580 795.700 951.700 796.000 ;
        RECT 952.860 795.700 972.980 796.000 ;
        RECT 974.140 795.700 994.260 796.000 ;
        RECT 995.420 795.700 1015.540 796.000 ;
        RECT 1016.700 795.700 1036.820 796.000 ;
        RECT 1037.980 795.700 1058.100 796.000 ;
        RECT 1059.260 795.700 1079.380 796.000 ;
        RECT 1080.540 795.700 1100.660 796.000 ;
        RECT 1101.820 795.700 1121.940 796.000 ;
        RECT 1123.100 795.700 1143.220 796.000 ;
        RECT 1144.380 795.700 1164.500 796.000 ;
        RECT 1165.660 795.700 1185.780 796.000 ;
        RECT 1186.940 795.700 1207.060 796.000 ;
        RECT 1208.220 795.700 1228.340 796.000 ;
        RECT 1229.500 795.700 1249.620 796.000 ;
        RECT 1250.780 795.700 1270.900 796.000 ;
        RECT 1272.060 795.700 1292.180 796.000 ;
        RECT 1293.340 795.700 1313.460 796.000 ;
        RECT 1314.620 795.700 1334.740 796.000 ;
        RECT 1335.900 795.700 1356.020 796.000 ;
        RECT 1357.180 795.700 1377.300 796.000 ;
        RECT 1378.460 795.700 1398.580 796.000 ;
        RECT 1399.740 795.700 1419.860 796.000 ;
        RECT 1421.020 795.700 1441.140 796.000 ;
        RECT 1442.300 795.700 1462.420 796.000 ;
        RECT 1463.580 795.700 1483.700 796.000 ;
        RECT 1484.860 795.700 1504.980 796.000 ;
        RECT 1506.140 795.700 1526.260 796.000 ;
        RECT 1527.420 795.700 1547.540 796.000 ;
        RECT 1548.700 795.700 1568.820 796.000 ;
        RECT 1569.980 795.700 1590.100 796.000 ;
        RECT 1591.260 795.700 1611.380 796.000 ;
        RECT 1612.540 795.700 1632.660 796.000 ;
        RECT 1633.820 795.700 1653.940 796.000 ;
        RECT 1655.100 795.700 1675.220 796.000 ;
        RECT 1676.380 795.700 1696.500 796.000 ;
        RECT 1697.660 795.700 1717.780 796.000 ;
        RECT 1718.940 795.700 1739.060 796.000 ;
        RECT 1740.220 795.700 1760.340 796.000 ;
        RECT 1761.500 795.700 1781.620 796.000 ;
        RECT 1782.780 795.700 1802.900 796.000 ;
        RECT 1804.060 795.700 1824.180 796.000 ;
        RECT 1825.340 795.700 1845.460 796.000 ;
        RECT 1846.620 795.700 1866.740 796.000 ;
        RECT 1867.900 795.700 1888.020 796.000 ;
        RECT 1889.180 795.700 1909.300 796.000 ;
        RECT 1910.460 795.700 1930.580 796.000 ;
        RECT 1931.740 795.700 1951.860 796.000 ;
        RECT 1953.020 795.700 1973.140 796.000 ;
        RECT 1974.300 795.700 1994.420 796.000 ;
        RECT 1995.580 795.700 2015.700 796.000 ;
        RECT 2016.860 795.700 2036.980 796.000 ;
        RECT 2038.140 795.700 2058.260 796.000 ;
        RECT 2059.420 795.700 2079.540 796.000 ;
        RECT 2080.700 795.700 2100.820 796.000 ;
        RECT 2101.980 795.700 2122.100 796.000 ;
        RECT 2123.260 795.700 2143.380 796.000 ;
        RECT 2144.540 795.700 2164.660 796.000 ;
        RECT 2165.820 795.700 2185.940 796.000 ;
        RECT 2187.100 795.700 2207.220 796.000 ;
        RECT 2208.380 795.700 2228.500 796.000 ;
        RECT 2229.660 795.700 2249.780 796.000 ;
        RECT 2250.940 795.700 2271.060 796.000 ;
        RECT 2272.220 795.700 2292.340 796.000 ;
        RECT 2293.500 795.700 2313.620 796.000 ;
        RECT 2314.780 795.700 2334.900 796.000 ;
        RECT 2336.060 795.700 2356.180 796.000 ;
        RECT 2357.340 795.700 2377.460 796.000 ;
        RECT 2378.620 795.700 2398.740 796.000 ;
        RECT 2399.900 795.700 2420.020 796.000 ;
        RECT 2421.180 795.700 2441.300 796.000 ;
        RECT 2442.460 795.700 2462.580 796.000 ;
        RECT 2463.740 795.700 2483.860 796.000 ;
        RECT 2485.020 795.700 2505.140 796.000 ;
        RECT 2506.300 795.700 2526.420 796.000 ;
        RECT 2527.580 795.700 2547.700 796.000 ;
        RECT 2548.860 795.700 2568.980 796.000 ;
        RECT 2570.140 795.700 2590.260 796.000 ;
        RECT 2591.420 795.700 2611.540 796.000 ;
        RECT 2612.700 795.700 2632.820 796.000 ;
        RECT 2633.980 795.700 2654.100 796.000 ;
        RECT 2655.260 795.700 2675.380 796.000 ;
        RECT 2676.540 795.700 2696.660 796.000 ;
        RECT 2697.820 795.700 2717.940 796.000 ;
        RECT 2719.100 795.700 2739.220 796.000 ;
        RECT 2740.380 795.700 2760.500 796.000 ;
        RECT 2761.660 795.700 2791.460 796.000 ;
        RECT 7.980 4.300 2791.460 795.700 ;
        RECT 7.980 4.000 34.420 4.300 ;
        RECT 35.580 4.000 37.780 4.300 ;
        RECT 38.940 4.000 41.140 4.300 ;
        RECT 42.300 4.000 44.500 4.300 ;
        RECT 45.660 4.000 47.860 4.300 ;
        RECT 49.020 4.000 51.220 4.300 ;
        RECT 52.380 4.000 54.580 4.300 ;
        RECT 55.740 4.000 57.940 4.300 ;
        RECT 59.100 4.000 61.300 4.300 ;
        RECT 62.460 4.000 64.660 4.300 ;
        RECT 65.820 4.000 68.020 4.300 ;
        RECT 69.180 4.000 71.380 4.300 ;
        RECT 72.540 4.000 74.740 4.300 ;
        RECT 75.900 4.000 78.100 4.300 ;
        RECT 79.260 4.000 81.460 4.300 ;
        RECT 82.620 4.000 84.820 4.300 ;
        RECT 85.980 4.000 88.180 4.300 ;
        RECT 89.340 4.000 91.540 4.300 ;
        RECT 92.700 4.000 94.900 4.300 ;
        RECT 96.060 4.000 98.260 4.300 ;
        RECT 99.420 4.000 101.620 4.300 ;
        RECT 102.780 4.000 104.980 4.300 ;
        RECT 106.140 4.000 108.340 4.300 ;
        RECT 109.500 4.000 111.700 4.300 ;
        RECT 112.860 4.000 115.060 4.300 ;
        RECT 116.220 4.000 118.420 4.300 ;
        RECT 119.580 4.000 121.780 4.300 ;
        RECT 122.940 4.000 125.140 4.300 ;
        RECT 126.300 4.000 128.500 4.300 ;
        RECT 129.660 4.000 131.860 4.300 ;
        RECT 133.020 4.000 135.220 4.300 ;
        RECT 136.380 4.000 138.580 4.300 ;
        RECT 139.740 4.000 141.940 4.300 ;
        RECT 143.100 4.000 145.300 4.300 ;
        RECT 146.460 4.000 148.660 4.300 ;
        RECT 149.820 4.000 152.020 4.300 ;
        RECT 153.180 4.000 155.380 4.300 ;
        RECT 156.540 4.000 158.740 4.300 ;
        RECT 159.900 4.000 162.100 4.300 ;
        RECT 163.260 4.000 165.460 4.300 ;
        RECT 166.620 4.000 168.820 4.300 ;
        RECT 169.980 4.000 172.180 4.300 ;
        RECT 173.340 4.000 175.540 4.300 ;
        RECT 176.700 4.000 178.900 4.300 ;
        RECT 180.060 4.000 182.260 4.300 ;
        RECT 183.420 4.000 185.620 4.300 ;
        RECT 186.780 4.000 188.980 4.300 ;
        RECT 190.140 4.000 192.340 4.300 ;
        RECT 193.500 4.000 195.700 4.300 ;
        RECT 196.860 4.000 199.060 4.300 ;
        RECT 200.220 4.000 202.420 4.300 ;
        RECT 203.580 4.000 205.780 4.300 ;
        RECT 206.940 4.000 209.140 4.300 ;
        RECT 210.300 4.000 212.500 4.300 ;
        RECT 213.660 4.000 215.860 4.300 ;
        RECT 217.020 4.000 219.220 4.300 ;
        RECT 220.380 4.000 222.580 4.300 ;
        RECT 223.740 4.000 225.940 4.300 ;
        RECT 227.100 4.000 229.300 4.300 ;
        RECT 230.460 4.000 232.660 4.300 ;
        RECT 233.820 4.000 236.020 4.300 ;
        RECT 237.180 4.000 239.380 4.300 ;
        RECT 240.540 4.000 242.740 4.300 ;
        RECT 243.900 4.000 246.100 4.300 ;
        RECT 247.260 4.000 249.460 4.300 ;
        RECT 250.620 4.000 252.820 4.300 ;
        RECT 253.980 4.000 256.180 4.300 ;
        RECT 257.340 4.000 259.540 4.300 ;
        RECT 260.700 4.000 262.900 4.300 ;
        RECT 264.060 4.000 266.260 4.300 ;
        RECT 267.420 4.000 269.620 4.300 ;
        RECT 270.780 4.000 272.980 4.300 ;
        RECT 274.140 4.000 276.340 4.300 ;
        RECT 277.500 4.000 279.700 4.300 ;
        RECT 280.860 4.000 283.060 4.300 ;
        RECT 284.220 4.000 286.420 4.300 ;
        RECT 287.580 4.000 289.780 4.300 ;
        RECT 290.940 4.000 293.140 4.300 ;
        RECT 294.300 4.000 296.500 4.300 ;
        RECT 297.660 4.000 299.860 4.300 ;
        RECT 301.020 4.000 303.220 4.300 ;
        RECT 304.380 4.000 306.580 4.300 ;
        RECT 307.740 4.000 309.940 4.300 ;
        RECT 311.100 4.000 313.300 4.300 ;
        RECT 314.460 4.000 316.660 4.300 ;
        RECT 317.820 4.000 320.020 4.300 ;
        RECT 321.180 4.000 323.380 4.300 ;
        RECT 324.540 4.000 326.740 4.300 ;
        RECT 327.900 4.000 330.100 4.300 ;
        RECT 331.260 4.000 333.460 4.300 ;
        RECT 334.620 4.000 336.820 4.300 ;
        RECT 337.980 4.000 340.180 4.300 ;
        RECT 341.340 4.000 343.540 4.300 ;
        RECT 344.700 4.000 346.900 4.300 ;
        RECT 348.060 4.000 350.260 4.300 ;
        RECT 351.420 4.000 353.620 4.300 ;
        RECT 354.780 4.000 356.980 4.300 ;
        RECT 358.140 4.000 360.340 4.300 ;
        RECT 361.500 4.000 363.700 4.300 ;
        RECT 364.860 4.000 367.060 4.300 ;
        RECT 368.220 4.000 370.420 4.300 ;
        RECT 371.580 4.000 373.780 4.300 ;
        RECT 374.940 4.000 377.140 4.300 ;
        RECT 378.300 4.000 380.500 4.300 ;
        RECT 381.660 4.000 383.860 4.300 ;
        RECT 385.020 4.000 387.220 4.300 ;
        RECT 388.380 4.000 390.580 4.300 ;
        RECT 391.740 4.000 393.940 4.300 ;
        RECT 395.100 4.000 397.300 4.300 ;
        RECT 398.460 4.000 400.660 4.300 ;
        RECT 401.820 4.000 404.020 4.300 ;
        RECT 405.180 4.000 407.380 4.300 ;
        RECT 408.540 4.000 410.740 4.300 ;
        RECT 411.900 4.000 414.100 4.300 ;
        RECT 415.260 4.000 417.460 4.300 ;
        RECT 418.620 4.000 420.820 4.300 ;
        RECT 421.980 4.000 424.180 4.300 ;
        RECT 425.340 4.000 427.540 4.300 ;
        RECT 428.700 4.000 430.900 4.300 ;
        RECT 432.060 4.000 434.260 4.300 ;
        RECT 435.420 4.000 437.620 4.300 ;
        RECT 438.780 4.000 440.980 4.300 ;
        RECT 442.140 4.000 444.340 4.300 ;
        RECT 445.500 4.000 447.700 4.300 ;
        RECT 448.860 4.000 451.060 4.300 ;
        RECT 452.220 4.000 454.420 4.300 ;
        RECT 455.580 4.000 457.780 4.300 ;
        RECT 458.940 4.000 461.140 4.300 ;
        RECT 462.300 4.000 464.500 4.300 ;
        RECT 465.660 4.000 467.860 4.300 ;
        RECT 469.020 4.000 471.220 4.300 ;
        RECT 472.380 4.000 474.580 4.300 ;
        RECT 475.740 4.000 477.940 4.300 ;
        RECT 479.100 4.000 481.300 4.300 ;
        RECT 482.460 4.000 484.660 4.300 ;
        RECT 485.820 4.000 488.020 4.300 ;
        RECT 489.180 4.000 491.380 4.300 ;
        RECT 492.540 4.000 494.740 4.300 ;
        RECT 495.900 4.000 498.100 4.300 ;
        RECT 499.260 4.000 501.460 4.300 ;
        RECT 502.620 4.000 504.820 4.300 ;
        RECT 505.980 4.000 508.180 4.300 ;
        RECT 509.340 4.000 511.540 4.300 ;
        RECT 512.700 4.000 514.900 4.300 ;
        RECT 516.060 4.000 518.260 4.300 ;
        RECT 519.420 4.000 521.620 4.300 ;
        RECT 522.780 4.000 524.980 4.300 ;
        RECT 526.140 4.000 528.340 4.300 ;
        RECT 529.500 4.000 531.700 4.300 ;
        RECT 532.860 4.000 535.060 4.300 ;
        RECT 536.220 4.000 538.420 4.300 ;
        RECT 539.580 4.000 541.780 4.300 ;
        RECT 542.940 4.000 545.140 4.300 ;
        RECT 546.300 4.000 548.500 4.300 ;
        RECT 549.660 4.000 551.860 4.300 ;
        RECT 553.020 4.000 555.220 4.300 ;
        RECT 556.380 4.000 558.580 4.300 ;
        RECT 559.740 4.000 561.940 4.300 ;
        RECT 563.100 4.000 565.300 4.300 ;
        RECT 566.460 4.000 568.660 4.300 ;
        RECT 569.820 4.000 572.020 4.300 ;
        RECT 573.180 4.000 575.380 4.300 ;
        RECT 576.540 4.000 578.740 4.300 ;
        RECT 579.900 4.000 582.100 4.300 ;
        RECT 583.260 4.000 585.460 4.300 ;
        RECT 586.620 4.000 588.820 4.300 ;
        RECT 589.980 4.000 592.180 4.300 ;
        RECT 593.340 4.000 595.540 4.300 ;
        RECT 596.700 4.000 598.900 4.300 ;
        RECT 600.060 4.000 602.260 4.300 ;
        RECT 603.420 4.000 605.620 4.300 ;
        RECT 606.780 4.000 608.980 4.300 ;
        RECT 610.140 4.000 612.340 4.300 ;
        RECT 613.500 4.000 615.700 4.300 ;
        RECT 616.860 4.000 619.060 4.300 ;
        RECT 620.220 4.000 622.420 4.300 ;
        RECT 623.580 4.000 625.780 4.300 ;
        RECT 626.940 4.000 629.140 4.300 ;
        RECT 630.300 4.000 632.500 4.300 ;
        RECT 633.660 4.000 635.860 4.300 ;
        RECT 637.020 4.000 639.220 4.300 ;
        RECT 640.380 4.000 642.580 4.300 ;
        RECT 643.740 4.000 645.940 4.300 ;
        RECT 647.100 4.000 649.300 4.300 ;
        RECT 650.460 4.000 652.660 4.300 ;
        RECT 653.820 4.000 656.020 4.300 ;
        RECT 657.180 4.000 659.380 4.300 ;
        RECT 660.540 4.000 662.740 4.300 ;
        RECT 663.900 4.000 666.100 4.300 ;
        RECT 667.260 4.000 669.460 4.300 ;
        RECT 670.620 4.000 672.820 4.300 ;
        RECT 673.980 4.000 676.180 4.300 ;
        RECT 677.340 4.000 679.540 4.300 ;
        RECT 680.700 4.000 682.900 4.300 ;
        RECT 684.060 4.000 686.260 4.300 ;
        RECT 687.420 4.000 689.620 4.300 ;
        RECT 690.780 4.000 692.980 4.300 ;
        RECT 694.140 4.000 696.340 4.300 ;
        RECT 697.500 4.000 699.700 4.300 ;
        RECT 700.860 4.000 703.060 4.300 ;
        RECT 704.220 4.000 706.420 4.300 ;
        RECT 707.580 4.000 709.780 4.300 ;
        RECT 710.940 4.000 713.140 4.300 ;
        RECT 714.300 4.000 716.500 4.300 ;
        RECT 717.660 4.000 719.860 4.300 ;
        RECT 721.020 4.000 723.220 4.300 ;
        RECT 724.380 4.000 726.580 4.300 ;
        RECT 727.740 4.000 729.940 4.300 ;
        RECT 731.100 4.000 733.300 4.300 ;
        RECT 734.460 4.000 736.660 4.300 ;
        RECT 737.820 4.000 740.020 4.300 ;
        RECT 741.180 4.000 743.380 4.300 ;
        RECT 744.540 4.000 746.740 4.300 ;
        RECT 747.900 4.000 750.100 4.300 ;
        RECT 751.260 4.000 753.460 4.300 ;
        RECT 754.620 4.000 756.820 4.300 ;
        RECT 757.980 4.000 760.180 4.300 ;
        RECT 761.340 4.000 763.540 4.300 ;
        RECT 764.700 4.000 766.900 4.300 ;
        RECT 768.060 4.000 770.260 4.300 ;
        RECT 771.420 4.000 773.620 4.300 ;
        RECT 774.780 4.000 776.980 4.300 ;
        RECT 778.140 4.000 780.340 4.300 ;
        RECT 781.500 4.000 783.700 4.300 ;
        RECT 784.860 4.000 787.060 4.300 ;
        RECT 788.220 4.000 790.420 4.300 ;
        RECT 791.580 4.000 793.780 4.300 ;
        RECT 794.940 4.000 797.140 4.300 ;
        RECT 798.300 4.000 800.500 4.300 ;
        RECT 801.660 4.000 803.860 4.300 ;
        RECT 805.020 4.000 807.220 4.300 ;
        RECT 808.380 4.000 810.580 4.300 ;
        RECT 811.740 4.000 813.940 4.300 ;
        RECT 815.100 4.000 817.300 4.300 ;
        RECT 818.460 4.000 820.660 4.300 ;
        RECT 821.820 4.000 824.020 4.300 ;
        RECT 825.180 4.000 827.380 4.300 ;
        RECT 828.540 4.000 830.740 4.300 ;
        RECT 831.900 4.000 834.100 4.300 ;
        RECT 835.260 4.000 837.460 4.300 ;
        RECT 838.620 4.000 840.820 4.300 ;
        RECT 841.980 4.000 844.180 4.300 ;
        RECT 845.340 4.000 847.540 4.300 ;
        RECT 848.700 4.000 850.900 4.300 ;
        RECT 852.060 4.000 854.260 4.300 ;
        RECT 855.420 4.000 857.620 4.300 ;
        RECT 858.780 4.000 860.980 4.300 ;
        RECT 862.140 4.000 864.340 4.300 ;
        RECT 865.500 4.000 867.700 4.300 ;
        RECT 868.860 4.000 871.060 4.300 ;
        RECT 872.220 4.000 874.420 4.300 ;
        RECT 875.580 4.000 877.780 4.300 ;
        RECT 878.940 4.000 881.140 4.300 ;
        RECT 882.300 4.000 884.500 4.300 ;
        RECT 885.660 4.000 887.860 4.300 ;
        RECT 889.020 4.000 891.220 4.300 ;
        RECT 892.380 4.000 894.580 4.300 ;
        RECT 895.740 4.000 897.940 4.300 ;
        RECT 899.100 4.000 901.300 4.300 ;
        RECT 902.460 4.000 904.660 4.300 ;
        RECT 905.820 4.000 908.020 4.300 ;
        RECT 909.180 4.000 911.380 4.300 ;
        RECT 912.540 4.000 914.740 4.300 ;
        RECT 915.900 4.000 918.100 4.300 ;
        RECT 919.260 4.000 921.460 4.300 ;
        RECT 922.620 4.000 924.820 4.300 ;
        RECT 925.980 4.000 928.180 4.300 ;
        RECT 929.340 4.000 931.540 4.300 ;
        RECT 932.700 4.000 934.900 4.300 ;
        RECT 936.060 4.000 938.260 4.300 ;
        RECT 939.420 4.000 941.620 4.300 ;
        RECT 942.780 4.000 944.980 4.300 ;
        RECT 946.140 4.000 948.340 4.300 ;
        RECT 949.500 4.000 951.700 4.300 ;
        RECT 952.860 4.000 955.060 4.300 ;
        RECT 956.220 4.000 958.420 4.300 ;
        RECT 959.580 4.000 961.780 4.300 ;
        RECT 962.940 4.000 965.140 4.300 ;
        RECT 966.300 4.000 968.500 4.300 ;
        RECT 969.660 4.000 971.860 4.300 ;
        RECT 973.020 4.000 975.220 4.300 ;
        RECT 976.380 4.000 978.580 4.300 ;
        RECT 979.740 4.000 981.940 4.300 ;
        RECT 983.100 4.000 985.300 4.300 ;
        RECT 986.460 4.000 988.660 4.300 ;
        RECT 989.820 4.000 992.020 4.300 ;
        RECT 993.180 4.000 995.380 4.300 ;
        RECT 996.540 4.000 998.740 4.300 ;
        RECT 999.900 4.000 1002.100 4.300 ;
        RECT 1003.260 4.000 1005.460 4.300 ;
        RECT 1006.620 4.000 1008.820 4.300 ;
        RECT 1009.980 4.000 1012.180 4.300 ;
        RECT 1013.340 4.000 1015.540 4.300 ;
        RECT 1016.700 4.000 1018.900 4.300 ;
        RECT 1020.060 4.000 1022.260 4.300 ;
        RECT 1023.420 4.000 1025.620 4.300 ;
        RECT 1026.780 4.000 1028.980 4.300 ;
        RECT 1030.140 4.000 1032.340 4.300 ;
        RECT 1033.500 4.000 1035.700 4.300 ;
        RECT 1036.860 4.000 1039.060 4.300 ;
        RECT 1040.220 4.000 1042.420 4.300 ;
        RECT 1043.580 4.000 1045.780 4.300 ;
        RECT 1046.940 4.000 1049.140 4.300 ;
        RECT 1050.300 4.000 1052.500 4.300 ;
        RECT 1053.660 4.000 1055.860 4.300 ;
        RECT 1057.020 4.000 1059.220 4.300 ;
        RECT 1060.380 4.000 1062.580 4.300 ;
        RECT 1063.740 4.000 1065.940 4.300 ;
        RECT 1067.100 4.000 1069.300 4.300 ;
        RECT 1070.460 4.000 1072.660 4.300 ;
        RECT 1073.820 4.000 1076.020 4.300 ;
        RECT 1077.180 4.000 1079.380 4.300 ;
        RECT 1080.540 4.000 1082.740 4.300 ;
        RECT 1083.900 4.000 1086.100 4.300 ;
        RECT 1087.260 4.000 1089.460 4.300 ;
        RECT 1090.620 4.000 1092.820 4.300 ;
        RECT 1093.980 4.000 1096.180 4.300 ;
        RECT 1097.340 4.000 1099.540 4.300 ;
        RECT 1100.700 4.000 1102.900 4.300 ;
        RECT 1104.060 4.000 1106.260 4.300 ;
        RECT 1107.420 4.000 1109.620 4.300 ;
        RECT 1110.780 4.000 1112.980 4.300 ;
        RECT 1114.140 4.000 1116.340 4.300 ;
        RECT 1117.500 4.000 1119.700 4.300 ;
        RECT 1120.860 4.000 1123.060 4.300 ;
        RECT 1124.220 4.000 1126.420 4.300 ;
        RECT 1127.580 4.000 1129.780 4.300 ;
        RECT 1130.940 4.000 1133.140 4.300 ;
        RECT 1134.300 4.000 1136.500 4.300 ;
        RECT 1137.660 4.000 1139.860 4.300 ;
        RECT 1141.020 4.000 1143.220 4.300 ;
        RECT 1144.380 4.000 1146.580 4.300 ;
        RECT 1147.740 4.000 1149.940 4.300 ;
        RECT 1151.100 4.000 1153.300 4.300 ;
        RECT 1154.460 4.000 1156.660 4.300 ;
        RECT 1157.820 4.000 1160.020 4.300 ;
        RECT 1161.180 4.000 1163.380 4.300 ;
        RECT 1164.540 4.000 1166.740 4.300 ;
        RECT 1167.900 4.000 1170.100 4.300 ;
        RECT 1171.260 4.000 1173.460 4.300 ;
        RECT 1174.620 4.000 1176.820 4.300 ;
        RECT 1177.980 4.000 1180.180 4.300 ;
        RECT 1181.340 4.000 1183.540 4.300 ;
        RECT 1184.700 4.000 1186.900 4.300 ;
        RECT 1188.060 4.000 1190.260 4.300 ;
        RECT 1191.420 4.000 1193.620 4.300 ;
        RECT 1194.780 4.000 1196.980 4.300 ;
        RECT 1198.140 4.000 1200.340 4.300 ;
        RECT 1201.500 4.000 1203.700 4.300 ;
        RECT 1204.860 4.000 1207.060 4.300 ;
        RECT 1208.220 4.000 1210.420 4.300 ;
        RECT 1211.580 4.000 1213.780 4.300 ;
        RECT 1214.940 4.000 1217.140 4.300 ;
        RECT 1218.300 4.000 1220.500 4.300 ;
        RECT 1221.660 4.000 1223.860 4.300 ;
        RECT 1225.020 4.000 1227.220 4.300 ;
        RECT 1228.380 4.000 1230.580 4.300 ;
        RECT 1231.740 4.000 1233.940 4.300 ;
        RECT 1235.100 4.000 1237.300 4.300 ;
        RECT 1238.460 4.000 1240.660 4.300 ;
        RECT 1241.820 4.000 1244.020 4.300 ;
        RECT 1245.180 4.000 1247.380 4.300 ;
        RECT 1248.540 4.000 1250.740 4.300 ;
        RECT 1251.900 4.000 1254.100 4.300 ;
        RECT 1255.260 4.000 1257.460 4.300 ;
        RECT 1258.620 4.000 1260.820 4.300 ;
        RECT 1261.980 4.000 1264.180 4.300 ;
        RECT 1265.340 4.000 1267.540 4.300 ;
        RECT 1268.700 4.000 1270.900 4.300 ;
        RECT 1272.060 4.000 1274.260 4.300 ;
        RECT 1275.420 4.000 1277.620 4.300 ;
        RECT 1278.780 4.000 1280.980 4.300 ;
        RECT 1282.140 4.000 1284.340 4.300 ;
        RECT 1285.500 4.000 1287.700 4.300 ;
        RECT 1288.860 4.000 1291.060 4.300 ;
        RECT 1292.220 4.000 1294.420 4.300 ;
        RECT 1295.580 4.000 1297.780 4.300 ;
        RECT 1298.940 4.000 1301.140 4.300 ;
        RECT 1302.300 4.000 1304.500 4.300 ;
        RECT 1305.660 4.000 1307.860 4.300 ;
        RECT 1309.020 4.000 1311.220 4.300 ;
        RECT 1312.380 4.000 1314.580 4.300 ;
        RECT 1315.740 4.000 1317.940 4.300 ;
        RECT 1319.100 4.000 1321.300 4.300 ;
        RECT 1322.460 4.000 1324.660 4.300 ;
        RECT 1325.820 4.000 1328.020 4.300 ;
        RECT 1329.180 4.000 1331.380 4.300 ;
        RECT 1332.540 4.000 1334.740 4.300 ;
        RECT 1335.900 4.000 1338.100 4.300 ;
        RECT 1339.260 4.000 1341.460 4.300 ;
        RECT 1342.620 4.000 1344.820 4.300 ;
        RECT 1345.980 4.000 1348.180 4.300 ;
        RECT 1349.340 4.000 1351.540 4.300 ;
        RECT 1352.700 4.000 1354.900 4.300 ;
        RECT 1356.060 4.000 1358.260 4.300 ;
        RECT 1359.420 4.000 1361.620 4.300 ;
        RECT 1362.780 4.000 1364.980 4.300 ;
        RECT 1366.140 4.000 1368.340 4.300 ;
        RECT 1369.500 4.000 1371.700 4.300 ;
        RECT 1372.860 4.000 1375.060 4.300 ;
        RECT 1376.220 4.000 1378.420 4.300 ;
        RECT 1379.580 4.000 1381.780 4.300 ;
        RECT 1382.940 4.000 1385.140 4.300 ;
        RECT 1386.300 4.000 1388.500 4.300 ;
        RECT 1389.660 4.000 1391.860 4.300 ;
        RECT 1393.020 4.000 1395.220 4.300 ;
        RECT 1396.380 4.000 1398.580 4.300 ;
        RECT 1399.740 4.000 1401.940 4.300 ;
        RECT 1403.100 4.000 1405.300 4.300 ;
        RECT 1406.460 4.000 1408.660 4.300 ;
        RECT 1409.820 4.000 1412.020 4.300 ;
        RECT 1413.180 4.000 1415.380 4.300 ;
        RECT 1416.540 4.000 1418.740 4.300 ;
        RECT 1419.900 4.000 1422.100 4.300 ;
        RECT 1423.260 4.000 1425.460 4.300 ;
        RECT 1426.620 4.000 1428.820 4.300 ;
        RECT 1429.980 4.000 1432.180 4.300 ;
        RECT 1433.340 4.000 1435.540 4.300 ;
        RECT 1436.700 4.000 1438.900 4.300 ;
        RECT 1440.060 4.000 1442.260 4.300 ;
        RECT 1443.420 4.000 1445.620 4.300 ;
        RECT 1446.780 4.000 1448.980 4.300 ;
        RECT 1450.140 4.000 1452.340 4.300 ;
        RECT 1453.500 4.000 1455.700 4.300 ;
        RECT 1456.860 4.000 1459.060 4.300 ;
        RECT 1460.220 4.000 1462.420 4.300 ;
        RECT 1463.580 4.000 1465.780 4.300 ;
        RECT 1466.940 4.000 1469.140 4.300 ;
        RECT 1470.300 4.000 1472.500 4.300 ;
        RECT 1473.660 4.000 1475.860 4.300 ;
        RECT 1477.020 4.000 1479.220 4.300 ;
        RECT 1480.380 4.000 1482.580 4.300 ;
        RECT 1483.740 4.000 1485.940 4.300 ;
        RECT 1487.100 4.000 1489.300 4.300 ;
        RECT 1490.460 4.000 1492.660 4.300 ;
        RECT 1493.820 4.000 1496.020 4.300 ;
        RECT 1497.180 4.000 1499.380 4.300 ;
        RECT 1500.540 4.000 1502.740 4.300 ;
        RECT 1503.900 4.000 1506.100 4.300 ;
        RECT 1507.260 4.000 1509.460 4.300 ;
        RECT 1510.620 4.000 1512.820 4.300 ;
        RECT 1513.980 4.000 1516.180 4.300 ;
        RECT 1517.340 4.000 1519.540 4.300 ;
        RECT 1520.700 4.000 1522.900 4.300 ;
        RECT 1524.060 4.000 1526.260 4.300 ;
        RECT 1527.420 4.000 1529.620 4.300 ;
        RECT 1530.780 4.000 1532.980 4.300 ;
        RECT 1534.140 4.000 1536.340 4.300 ;
        RECT 1537.500 4.000 1539.700 4.300 ;
        RECT 1540.860 4.000 1543.060 4.300 ;
        RECT 1544.220 4.000 1546.420 4.300 ;
        RECT 1547.580 4.000 1549.780 4.300 ;
        RECT 1550.940 4.000 1553.140 4.300 ;
        RECT 1554.300 4.000 1556.500 4.300 ;
        RECT 1557.660 4.000 1559.860 4.300 ;
        RECT 1561.020 4.000 1563.220 4.300 ;
        RECT 1564.380 4.000 1566.580 4.300 ;
        RECT 1567.740 4.000 1569.940 4.300 ;
        RECT 1571.100 4.000 1573.300 4.300 ;
        RECT 1574.460 4.000 1576.660 4.300 ;
        RECT 1577.820 4.000 1580.020 4.300 ;
        RECT 1581.180 4.000 1583.380 4.300 ;
        RECT 1584.540 4.000 1586.740 4.300 ;
        RECT 1587.900 4.000 1590.100 4.300 ;
        RECT 1591.260 4.000 1593.460 4.300 ;
        RECT 1594.620 4.000 1596.820 4.300 ;
        RECT 1597.980 4.000 1600.180 4.300 ;
        RECT 1601.340 4.000 1603.540 4.300 ;
        RECT 1604.700 4.000 1606.900 4.300 ;
        RECT 1608.060 4.000 1610.260 4.300 ;
        RECT 1611.420 4.000 1613.620 4.300 ;
        RECT 1614.780 4.000 1616.980 4.300 ;
        RECT 1618.140 4.000 1620.340 4.300 ;
        RECT 1621.500 4.000 1623.700 4.300 ;
        RECT 1624.860 4.000 1627.060 4.300 ;
        RECT 1628.220 4.000 1630.420 4.300 ;
        RECT 1631.580 4.000 1633.780 4.300 ;
        RECT 1634.940 4.000 1637.140 4.300 ;
        RECT 1638.300 4.000 1640.500 4.300 ;
        RECT 1641.660 4.000 1643.860 4.300 ;
        RECT 1645.020 4.000 1647.220 4.300 ;
        RECT 1648.380 4.000 1650.580 4.300 ;
        RECT 1651.740 4.000 1653.940 4.300 ;
        RECT 1655.100 4.000 1657.300 4.300 ;
        RECT 1658.460 4.000 1660.660 4.300 ;
        RECT 1661.820 4.000 1664.020 4.300 ;
        RECT 1665.180 4.000 1667.380 4.300 ;
        RECT 1668.540 4.000 1670.740 4.300 ;
        RECT 1671.900 4.000 1674.100 4.300 ;
        RECT 1675.260 4.000 1677.460 4.300 ;
        RECT 1678.620 4.000 1680.820 4.300 ;
        RECT 1681.980 4.000 1684.180 4.300 ;
        RECT 1685.340 4.000 1687.540 4.300 ;
        RECT 1688.700 4.000 1690.900 4.300 ;
        RECT 1692.060 4.000 1694.260 4.300 ;
        RECT 1695.420 4.000 1697.620 4.300 ;
        RECT 1698.780 4.000 1700.980 4.300 ;
        RECT 1702.140 4.000 1704.340 4.300 ;
        RECT 1705.500 4.000 1707.700 4.300 ;
        RECT 1708.860 4.000 1711.060 4.300 ;
        RECT 1712.220 4.000 1714.420 4.300 ;
        RECT 1715.580 4.000 1717.780 4.300 ;
        RECT 1718.940 4.000 1721.140 4.300 ;
        RECT 1722.300 4.000 1724.500 4.300 ;
        RECT 1725.660 4.000 1727.860 4.300 ;
        RECT 1729.020 4.000 1731.220 4.300 ;
        RECT 1732.380 4.000 1734.580 4.300 ;
        RECT 1735.740 4.000 1737.940 4.300 ;
        RECT 1739.100 4.000 1741.300 4.300 ;
        RECT 1742.460 4.000 1744.660 4.300 ;
        RECT 1745.820 4.000 1748.020 4.300 ;
        RECT 1749.180 4.000 1751.380 4.300 ;
        RECT 1752.540 4.000 1754.740 4.300 ;
        RECT 1755.900 4.000 1758.100 4.300 ;
        RECT 1759.260 4.000 1761.460 4.300 ;
        RECT 1762.620 4.000 1764.820 4.300 ;
        RECT 1765.980 4.000 1768.180 4.300 ;
        RECT 1769.340 4.000 1771.540 4.300 ;
        RECT 1772.700 4.000 1774.900 4.300 ;
        RECT 1776.060 4.000 1778.260 4.300 ;
        RECT 1779.420 4.000 1781.620 4.300 ;
        RECT 1782.780 4.000 1784.980 4.300 ;
        RECT 1786.140 4.000 1788.340 4.300 ;
        RECT 1789.500 4.000 1791.700 4.300 ;
        RECT 1792.860 4.000 1795.060 4.300 ;
        RECT 1796.220 4.000 1798.420 4.300 ;
        RECT 1799.580 4.000 1801.780 4.300 ;
        RECT 1802.940 4.000 1805.140 4.300 ;
        RECT 1806.300 4.000 1808.500 4.300 ;
        RECT 1809.660 4.000 1811.860 4.300 ;
        RECT 1813.020 4.000 1815.220 4.300 ;
        RECT 1816.380 4.000 1818.580 4.300 ;
        RECT 1819.740 4.000 1821.940 4.300 ;
        RECT 1823.100 4.000 1825.300 4.300 ;
        RECT 1826.460 4.000 1828.660 4.300 ;
        RECT 1829.820 4.000 1832.020 4.300 ;
        RECT 1833.180 4.000 1835.380 4.300 ;
        RECT 1836.540 4.000 1838.740 4.300 ;
        RECT 1839.900 4.000 1842.100 4.300 ;
        RECT 1843.260 4.000 1845.460 4.300 ;
        RECT 1846.620 4.000 1848.820 4.300 ;
        RECT 1849.980 4.000 1852.180 4.300 ;
        RECT 1853.340 4.000 1855.540 4.300 ;
        RECT 1856.700 4.000 1858.900 4.300 ;
        RECT 1860.060 4.000 1862.260 4.300 ;
        RECT 1863.420 4.000 1865.620 4.300 ;
        RECT 1866.780 4.000 1868.980 4.300 ;
        RECT 1870.140 4.000 1872.340 4.300 ;
        RECT 1873.500 4.000 1875.700 4.300 ;
        RECT 1876.860 4.000 1879.060 4.300 ;
        RECT 1880.220 4.000 1882.420 4.300 ;
        RECT 1883.580 4.000 1885.780 4.300 ;
        RECT 1886.940 4.000 1889.140 4.300 ;
        RECT 1890.300 4.000 1892.500 4.300 ;
        RECT 1893.660 4.000 1895.860 4.300 ;
        RECT 1897.020 4.000 1899.220 4.300 ;
        RECT 1900.380 4.000 1902.580 4.300 ;
        RECT 1903.740 4.000 1905.940 4.300 ;
        RECT 1907.100 4.000 1909.300 4.300 ;
        RECT 1910.460 4.000 1912.660 4.300 ;
        RECT 1913.820 4.000 1916.020 4.300 ;
        RECT 1917.180 4.000 1919.380 4.300 ;
        RECT 1920.540 4.000 1922.740 4.300 ;
        RECT 1923.900 4.000 1926.100 4.300 ;
        RECT 1927.260 4.000 1929.460 4.300 ;
        RECT 1930.620 4.000 1932.820 4.300 ;
        RECT 1933.980 4.000 1936.180 4.300 ;
        RECT 1937.340 4.000 1939.540 4.300 ;
        RECT 1940.700 4.000 1942.900 4.300 ;
        RECT 1944.060 4.000 1946.260 4.300 ;
        RECT 1947.420 4.000 1949.620 4.300 ;
        RECT 1950.780 4.000 1952.980 4.300 ;
        RECT 1954.140 4.000 1956.340 4.300 ;
        RECT 1957.500 4.000 1959.700 4.300 ;
        RECT 1960.860 4.000 1963.060 4.300 ;
        RECT 1964.220 4.000 1966.420 4.300 ;
        RECT 1967.580 4.000 1969.780 4.300 ;
        RECT 1970.940 4.000 1973.140 4.300 ;
        RECT 1974.300 4.000 1976.500 4.300 ;
        RECT 1977.660 4.000 1979.860 4.300 ;
        RECT 1981.020 4.000 1983.220 4.300 ;
        RECT 1984.380 4.000 1986.580 4.300 ;
        RECT 1987.740 4.000 1989.940 4.300 ;
        RECT 1991.100 4.000 1993.300 4.300 ;
        RECT 1994.460 4.000 1996.660 4.300 ;
        RECT 1997.820 4.000 2000.020 4.300 ;
        RECT 2001.180 4.000 2003.380 4.300 ;
        RECT 2004.540 4.000 2006.740 4.300 ;
        RECT 2007.900 4.000 2010.100 4.300 ;
        RECT 2011.260 4.000 2013.460 4.300 ;
        RECT 2014.620 4.000 2016.820 4.300 ;
        RECT 2017.980 4.000 2020.180 4.300 ;
        RECT 2021.340 4.000 2023.540 4.300 ;
        RECT 2024.700 4.000 2026.900 4.300 ;
        RECT 2028.060 4.000 2030.260 4.300 ;
        RECT 2031.420 4.000 2033.620 4.300 ;
        RECT 2034.780 4.000 2036.980 4.300 ;
        RECT 2038.140 4.000 2040.340 4.300 ;
        RECT 2041.500 4.000 2043.700 4.300 ;
        RECT 2044.860 4.000 2047.060 4.300 ;
        RECT 2048.220 4.000 2050.420 4.300 ;
        RECT 2051.580 4.000 2053.780 4.300 ;
        RECT 2054.940 4.000 2057.140 4.300 ;
        RECT 2058.300 4.000 2060.500 4.300 ;
        RECT 2061.660 4.000 2063.860 4.300 ;
        RECT 2065.020 4.000 2067.220 4.300 ;
        RECT 2068.380 4.000 2070.580 4.300 ;
        RECT 2071.740 4.000 2073.940 4.300 ;
        RECT 2075.100 4.000 2077.300 4.300 ;
        RECT 2078.460 4.000 2080.660 4.300 ;
        RECT 2081.820 4.000 2084.020 4.300 ;
        RECT 2085.180 4.000 2087.380 4.300 ;
        RECT 2088.540 4.000 2090.740 4.300 ;
        RECT 2091.900 4.000 2094.100 4.300 ;
        RECT 2095.260 4.000 2097.460 4.300 ;
        RECT 2098.620 4.000 2100.820 4.300 ;
        RECT 2101.980 4.000 2104.180 4.300 ;
        RECT 2105.340 4.000 2107.540 4.300 ;
        RECT 2108.700 4.000 2110.900 4.300 ;
        RECT 2112.060 4.000 2114.260 4.300 ;
        RECT 2115.420 4.000 2117.620 4.300 ;
        RECT 2118.780 4.000 2120.980 4.300 ;
        RECT 2122.140 4.000 2124.340 4.300 ;
        RECT 2125.500 4.000 2127.700 4.300 ;
        RECT 2128.860 4.000 2131.060 4.300 ;
        RECT 2132.220 4.000 2134.420 4.300 ;
        RECT 2135.580 4.000 2137.780 4.300 ;
        RECT 2138.940 4.000 2141.140 4.300 ;
        RECT 2142.300 4.000 2144.500 4.300 ;
        RECT 2145.660 4.000 2147.860 4.300 ;
        RECT 2149.020 4.000 2151.220 4.300 ;
        RECT 2152.380 4.000 2154.580 4.300 ;
        RECT 2155.740 4.000 2157.940 4.300 ;
        RECT 2159.100 4.000 2161.300 4.300 ;
        RECT 2162.460 4.000 2164.660 4.300 ;
        RECT 2165.820 4.000 2168.020 4.300 ;
        RECT 2169.180 4.000 2171.380 4.300 ;
        RECT 2172.540 4.000 2174.740 4.300 ;
        RECT 2175.900 4.000 2178.100 4.300 ;
        RECT 2179.260 4.000 2181.460 4.300 ;
        RECT 2182.620 4.000 2184.820 4.300 ;
        RECT 2185.980 4.000 2188.180 4.300 ;
        RECT 2189.340 4.000 2191.540 4.300 ;
        RECT 2192.700 4.000 2194.900 4.300 ;
        RECT 2196.060 4.000 2198.260 4.300 ;
        RECT 2199.420 4.000 2201.620 4.300 ;
        RECT 2202.780 4.000 2204.980 4.300 ;
        RECT 2206.140 4.000 2208.340 4.300 ;
        RECT 2209.500 4.000 2211.700 4.300 ;
        RECT 2212.860 4.000 2215.060 4.300 ;
        RECT 2216.220 4.000 2218.420 4.300 ;
        RECT 2219.580 4.000 2221.780 4.300 ;
        RECT 2222.940 4.000 2225.140 4.300 ;
        RECT 2226.300 4.000 2228.500 4.300 ;
        RECT 2229.660 4.000 2231.860 4.300 ;
        RECT 2233.020 4.000 2235.220 4.300 ;
        RECT 2236.380 4.000 2238.580 4.300 ;
        RECT 2239.740 4.000 2241.940 4.300 ;
        RECT 2243.100 4.000 2245.300 4.300 ;
        RECT 2246.460 4.000 2248.660 4.300 ;
        RECT 2249.820 4.000 2252.020 4.300 ;
        RECT 2253.180 4.000 2255.380 4.300 ;
        RECT 2256.540 4.000 2258.740 4.300 ;
        RECT 2259.900 4.000 2262.100 4.300 ;
        RECT 2263.260 4.000 2265.460 4.300 ;
        RECT 2266.620 4.000 2268.820 4.300 ;
        RECT 2269.980 4.000 2272.180 4.300 ;
        RECT 2273.340 4.000 2275.540 4.300 ;
        RECT 2276.700 4.000 2278.900 4.300 ;
        RECT 2280.060 4.000 2282.260 4.300 ;
        RECT 2283.420 4.000 2285.620 4.300 ;
        RECT 2286.780 4.000 2288.980 4.300 ;
        RECT 2290.140 4.000 2292.340 4.300 ;
        RECT 2293.500 4.000 2295.700 4.300 ;
        RECT 2296.860 4.000 2299.060 4.300 ;
        RECT 2300.220 4.000 2302.420 4.300 ;
        RECT 2303.580 4.000 2305.780 4.300 ;
        RECT 2306.940 4.000 2309.140 4.300 ;
        RECT 2310.300 4.000 2312.500 4.300 ;
        RECT 2313.660 4.000 2315.860 4.300 ;
        RECT 2317.020 4.000 2319.220 4.300 ;
        RECT 2320.380 4.000 2322.580 4.300 ;
        RECT 2323.740 4.000 2325.940 4.300 ;
        RECT 2327.100 4.000 2329.300 4.300 ;
        RECT 2330.460 4.000 2332.660 4.300 ;
        RECT 2333.820 4.000 2336.020 4.300 ;
        RECT 2337.180 4.000 2339.380 4.300 ;
        RECT 2340.540 4.000 2342.740 4.300 ;
        RECT 2343.900 4.000 2346.100 4.300 ;
        RECT 2347.260 4.000 2349.460 4.300 ;
        RECT 2350.620 4.000 2352.820 4.300 ;
        RECT 2353.980 4.000 2356.180 4.300 ;
        RECT 2357.340 4.000 2359.540 4.300 ;
        RECT 2360.700 4.000 2362.900 4.300 ;
        RECT 2364.060 4.000 2366.260 4.300 ;
        RECT 2367.420 4.000 2369.620 4.300 ;
        RECT 2370.780 4.000 2372.980 4.300 ;
        RECT 2374.140 4.000 2376.340 4.300 ;
        RECT 2377.500 4.000 2379.700 4.300 ;
        RECT 2380.860 4.000 2383.060 4.300 ;
        RECT 2384.220 4.000 2386.420 4.300 ;
        RECT 2387.580 4.000 2389.780 4.300 ;
        RECT 2390.940 4.000 2393.140 4.300 ;
        RECT 2394.300 4.000 2396.500 4.300 ;
        RECT 2397.660 4.000 2399.860 4.300 ;
        RECT 2401.020 4.000 2403.220 4.300 ;
        RECT 2404.380 4.000 2406.580 4.300 ;
        RECT 2407.740 4.000 2409.940 4.300 ;
        RECT 2411.100 4.000 2413.300 4.300 ;
        RECT 2414.460 4.000 2416.660 4.300 ;
        RECT 2417.820 4.000 2420.020 4.300 ;
        RECT 2421.180 4.000 2423.380 4.300 ;
        RECT 2424.540 4.000 2426.740 4.300 ;
        RECT 2427.900 4.000 2430.100 4.300 ;
        RECT 2431.260 4.000 2433.460 4.300 ;
        RECT 2434.620 4.000 2436.820 4.300 ;
        RECT 2437.980 4.000 2440.180 4.300 ;
        RECT 2441.340 4.000 2443.540 4.300 ;
        RECT 2444.700 4.000 2446.900 4.300 ;
        RECT 2448.060 4.000 2450.260 4.300 ;
        RECT 2451.420 4.000 2453.620 4.300 ;
        RECT 2454.780 4.000 2456.980 4.300 ;
        RECT 2458.140 4.000 2460.340 4.300 ;
        RECT 2461.500 4.000 2463.700 4.300 ;
        RECT 2464.860 4.000 2467.060 4.300 ;
        RECT 2468.220 4.000 2470.420 4.300 ;
        RECT 2471.580 4.000 2473.780 4.300 ;
        RECT 2474.940 4.000 2477.140 4.300 ;
        RECT 2478.300 4.000 2480.500 4.300 ;
        RECT 2481.660 4.000 2483.860 4.300 ;
        RECT 2485.020 4.000 2487.220 4.300 ;
        RECT 2488.380 4.000 2490.580 4.300 ;
        RECT 2491.740 4.000 2493.940 4.300 ;
        RECT 2495.100 4.000 2497.300 4.300 ;
        RECT 2498.460 4.000 2500.660 4.300 ;
        RECT 2501.820 4.000 2504.020 4.300 ;
        RECT 2505.180 4.000 2507.380 4.300 ;
        RECT 2508.540 4.000 2510.740 4.300 ;
        RECT 2511.900 4.000 2514.100 4.300 ;
        RECT 2515.260 4.000 2517.460 4.300 ;
        RECT 2518.620 4.000 2520.820 4.300 ;
        RECT 2521.980 4.000 2524.180 4.300 ;
        RECT 2525.340 4.000 2527.540 4.300 ;
        RECT 2528.700 4.000 2530.900 4.300 ;
        RECT 2532.060 4.000 2534.260 4.300 ;
        RECT 2535.420 4.000 2537.620 4.300 ;
        RECT 2538.780 4.000 2540.980 4.300 ;
        RECT 2542.140 4.000 2544.340 4.300 ;
        RECT 2545.500 4.000 2547.700 4.300 ;
        RECT 2548.860 4.000 2551.060 4.300 ;
        RECT 2552.220 4.000 2554.420 4.300 ;
        RECT 2555.580 4.000 2557.780 4.300 ;
        RECT 2558.940 4.000 2561.140 4.300 ;
        RECT 2562.300 4.000 2564.500 4.300 ;
        RECT 2565.660 4.000 2567.860 4.300 ;
        RECT 2569.020 4.000 2571.220 4.300 ;
        RECT 2572.380 4.000 2574.580 4.300 ;
        RECT 2575.740 4.000 2577.940 4.300 ;
        RECT 2579.100 4.000 2581.300 4.300 ;
        RECT 2582.460 4.000 2584.660 4.300 ;
        RECT 2585.820 4.000 2588.020 4.300 ;
        RECT 2589.180 4.000 2591.380 4.300 ;
        RECT 2592.540 4.000 2594.740 4.300 ;
        RECT 2595.900 4.000 2598.100 4.300 ;
        RECT 2599.260 4.000 2601.460 4.300 ;
        RECT 2602.620 4.000 2604.820 4.300 ;
        RECT 2605.980 4.000 2608.180 4.300 ;
        RECT 2609.340 4.000 2611.540 4.300 ;
        RECT 2612.700 4.000 2614.900 4.300 ;
        RECT 2616.060 4.000 2618.260 4.300 ;
        RECT 2619.420 4.000 2621.620 4.300 ;
        RECT 2622.780 4.000 2624.980 4.300 ;
        RECT 2626.140 4.000 2628.340 4.300 ;
        RECT 2629.500 4.000 2631.700 4.300 ;
        RECT 2632.860 4.000 2635.060 4.300 ;
        RECT 2636.220 4.000 2638.420 4.300 ;
        RECT 2639.580 4.000 2641.780 4.300 ;
        RECT 2642.940 4.000 2645.140 4.300 ;
        RECT 2646.300 4.000 2648.500 4.300 ;
        RECT 2649.660 4.000 2651.860 4.300 ;
        RECT 2653.020 4.000 2655.220 4.300 ;
        RECT 2656.380 4.000 2658.580 4.300 ;
        RECT 2659.740 4.000 2661.940 4.300 ;
        RECT 2663.100 4.000 2665.300 4.300 ;
        RECT 2666.460 4.000 2668.660 4.300 ;
        RECT 2669.820 4.000 2672.020 4.300 ;
        RECT 2673.180 4.000 2675.380 4.300 ;
        RECT 2676.540 4.000 2678.740 4.300 ;
        RECT 2679.900 4.000 2682.100 4.300 ;
        RECT 2683.260 4.000 2685.460 4.300 ;
        RECT 2686.620 4.000 2688.820 4.300 ;
        RECT 2689.980 4.000 2692.180 4.300 ;
        RECT 2693.340 4.000 2695.540 4.300 ;
        RECT 2696.700 4.000 2698.900 4.300 ;
        RECT 2700.060 4.000 2702.260 4.300 ;
        RECT 2703.420 4.000 2705.620 4.300 ;
        RECT 2706.780 4.000 2708.980 4.300 ;
        RECT 2710.140 4.000 2712.340 4.300 ;
        RECT 2713.500 4.000 2715.700 4.300 ;
        RECT 2716.860 4.000 2719.060 4.300 ;
        RECT 2720.220 4.000 2722.420 4.300 ;
        RECT 2723.580 4.000 2725.780 4.300 ;
        RECT 2726.940 4.000 2729.140 4.300 ;
        RECT 2730.300 4.000 2732.500 4.300 ;
        RECT 2733.660 4.000 2735.860 4.300 ;
        RECT 2737.020 4.000 2739.220 4.300 ;
        RECT 2740.380 4.000 2742.580 4.300 ;
        RECT 2743.740 4.000 2745.940 4.300 ;
        RECT 2747.100 4.000 2749.300 4.300 ;
        RECT 2750.460 4.000 2752.660 4.300 ;
        RECT 2753.820 4.000 2756.020 4.300 ;
        RECT 2757.180 4.000 2759.380 4.300 ;
        RECT 2760.540 4.000 2762.740 4.300 ;
        RECT 2763.900 4.000 2791.460 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 699.740 2796.000 793.380 ;
        RECT 4.300 99.380 2795.700 699.740 ;
        RECT 4.000 15.540 2796.000 99.380 ;
      LAYER Metal4 ;
        RECT 777.420 763.930 789.940 774.390 ;
        RECT 792.140 763.930 866.740 774.390 ;
        RECT 868.940 763.930 943.540 774.390 ;
        RECT 945.740 763.930 1020.340 774.390 ;
        RECT 1022.540 763.930 1097.140 774.390 ;
        RECT 1099.340 763.930 1173.940 774.390 ;
        RECT 1176.140 763.930 1250.740 774.390 ;
        RECT 1252.940 763.930 1327.540 774.390 ;
        RECT 1329.740 763.930 1404.340 774.390 ;
        RECT 1406.540 763.930 1481.140 774.390 ;
        RECT 1483.340 763.930 1557.940 774.390 ;
        RECT 1560.140 763.930 1634.740 774.390 ;
        RECT 1636.940 763.930 1711.540 774.390 ;
        RECT 1713.740 763.930 1747.620 774.390 ;
  END
END tjrpu
END LIBRARY

