magic
tech gf180mcuD
magscale 1 10
timestamp 1701035930
<< nwell >>
rect 1258 196377 198662 196870
rect 1258 196352 78396 196377
rect 1258 195623 58989 195648
rect 1258 194809 198662 195623
rect 1258 194784 69629 194809
rect 1258 194055 46109 194080
rect 1258 193241 198662 194055
rect 1258 193216 34349 193241
rect 1258 192487 67725 192512
rect 1258 191673 198662 192487
rect 1258 191648 39389 191673
rect 1258 190919 45437 190944
rect 1258 190105 198662 190919
rect 1258 190080 56301 190105
rect 1258 189351 31144 189376
rect 1258 188537 198662 189351
rect 1258 188512 33341 188537
rect 1258 187783 30429 187808
rect 1258 186969 198662 187783
rect 1258 186944 39613 186969
rect 1258 186215 44317 186240
rect 1258 185401 198662 186215
rect 1258 185376 71869 185401
rect 1258 184647 27517 184672
rect 1258 183833 198662 184647
rect 1258 183808 65709 183833
rect 1258 183079 27181 183104
rect 1258 182265 198662 183079
rect 1258 182240 54845 182265
rect 1258 181511 43757 181536
rect 1258 180697 198662 181511
rect 1258 180672 23821 180697
rect 1258 179943 38269 179968
rect 1258 179129 198662 179943
rect 1258 179104 24605 179129
rect 1258 178375 49693 178400
rect 1258 177561 198662 178375
rect 1258 177536 87144 177561
rect 1258 176807 43757 176832
rect 1258 175993 198662 176807
rect 1258 175968 65597 175993
rect 1258 175239 22589 175264
rect 1258 174425 198662 175239
rect 1258 174400 22141 174425
rect 1258 173671 90125 173696
rect 1258 172857 198662 173671
rect 1258 172832 96509 172857
rect 1258 172103 37149 172128
rect 1258 171289 198662 172103
rect 1258 171264 42120 171289
rect 1258 170535 18221 170560
rect 1258 169721 198662 170535
rect 1258 169696 22477 169721
rect 1258 168967 28861 168992
rect 1258 168153 198662 168967
rect 1258 168128 16765 168153
rect 1258 167399 12173 167424
rect 1258 166585 198662 167399
rect 1258 166560 10829 166585
rect 1258 165831 74893 165856
rect 1258 165017 198662 165831
rect 1258 164992 15869 165017
rect 1258 164263 22141 164288
rect 1258 163449 198662 164263
rect 1258 163424 22141 163449
rect 1258 162695 10381 162720
rect 1258 161881 198662 162695
rect 1258 161856 9149 161881
rect 1258 161127 4557 161152
rect 1258 160313 198662 161127
rect 1258 160288 27861 160313
rect 1258 159559 4893 159584
rect 1258 158745 198662 159559
rect 1258 158720 2989 158745
rect 1258 157991 20909 158016
rect 1258 157177 198662 157991
rect 1258 157152 26983 157177
rect 1258 156423 20168 156448
rect 1258 155609 198662 156423
rect 1258 155584 26983 155609
rect 1258 154855 3661 154880
rect 1258 154041 198662 154855
rect 1258 154016 2989 154041
rect 1258 153287 68061 153312
rect 1258 152473 198662 153287
rect 1258 152448 34125 152473
rect 1258 151719 21917 151744
rect 1258 150905 198662 151719
rect 1258 150880 17549 150905
rect 1258 150151 3213 150176
rect 1258 149337 198662 150151
rect 1258 149312 9485 149337
rect 1258 148583 3213 148608
rect 1258 147769 198662 148583
rect 1258 147744 37821 147769
rect 1258 147015 20797 147040
rect 1258 146201 198662 147015
rect 1258 146176 143727 146201
rect 1258 145447 59793 145472
rect 1258 144633 198662 145447
rect 1258 144608 2989 144633
rect 1258 143879 3437 143904
rect 1258 143065 198662 143879
rect 1258 143040 23597 143065
rect 1258 142311 61135 142336
rect 1258 141497 198662 142311
rect 1258 141472 62481 141497
rect 1258 140743 21357 140768
rect 1258 139929 198662 140743
rect 1258 139904 10829 139929
rect 1258 139175 3773 139200
rect 1258 138361 198662 139175
rect 1258 138336 2989 138361
rect 1258 137607 45370 137632
rect 1258 136793 198662 137607
rect 1258 136768 16808 136793
rect 1258 136039 3213 136064
rect 1258 135225 198662 136039
rect 1258 135200 39432 135225
rect 1258 134471 10381 134496
rect 1258 133657 198662 134471
rect 1258 133632 9261 133657
rect 1258 132903 3885 132928
rect 1258 132089 198662 132903
rect 1258 132064 40509 132089
rect 1258 131335 4333 131360
rect 1258 130521 198662 131335
rect 1258 130496 2989 130521
rect 1258 129767 109566 129792
rect 1258 128953 198662 129767
rect 1258 128928 37821 128953
rect 1258 128199 21581 128224
rect 1258 127385 198662 128199
rect 1258 127360 9821 127385
rect 1258 126631 4893 126656
rect 1258 125817 198662 126631
rect 1258 125792 2989 125817
rect 1258 125063 37597 125088
rect 1258 124249 198662 125063
rect 1258 124224 34237 124249
rect 1258 123495 19453 123520
rect 1258 122681 198662 123495
rect 1258 122656 8701 122681
rect 1258 121927 3325 121952
rect 1258 121113 198662 121927
rect 1258 121088 2989 121113
rect 1258 120359 3997 120384
rect 1258 119545 198662 120359
rect 1258 119520 22737 119545
rect 1258 118791 12285 118816
rect 1258 117977 198662 118791
rect 1258 117952 37821 117977
rect 1258 117223 30429 117248
rect 1258 116409 198662 117223
rect 1258 116384 18221 116409
rect 1258 115655 10381 115680
rect 1258 114841 198662 115655
rect 1258 114816 2877 114841
rect 1258 114087 2989 114112
rect 1258 113273 198662 114087
rect 1258 113248 7805 113273
rect 1258 112519 30429 112544
rect 1258 111705 198662 112519
rect 1258 111680 10829 111705
rect 1258 110951 12509 110976
rect 1258 110137 198662 110951
rect 1258 110112 47229 110137
rect 1258 109383 3325 109408
rect 1258 108569 198662 109383
rect 1258 108544 2989 108569
rect 1258 107815 36632 107840
rect 1258 107001 198662 107815
rect 1258 106976 39389 107001
rect 1258 106247 10381 106272
rect 1258 105433 198662 106247
rect 1258 105408 14525 105433
rect 1258 104679 3661 104704
rect 1258 103865 198662 104679
rect 1258 103840 6573 103865
rect 1258 103111 2989 103136
rect 1258 102297 198662 103111
rect 1258 102272 123622 102297
rect 1258 101543 20685 101568
rect 1258 100729 198662 101543
rect 1258 100704 48013 100729
rect 1258 99975 10717 100000
rect 1258 99161 198662 99975
rect 1258 99136 10381 99161
rect 1258 98407 5341 98432
rect 1258 97593 198662 98407
rect 1258 97568 2877 97593
rect 1258 96839 4669 96864
rect 1258 96025 198662 96839
rect 1258 96000 46109 96025
rect 1258 95271 10829 95296
rect 1258 94457 198662 95271
rect 1258 94432 10269 94457
rect 1258 93703 42413 93728
rect 1258 92889 198662 93703
rect 1258 92864 6461 92889
rect 1258 92135 13517 92160
rect 1258 91321 198662 92135
rect 1258 91296 25165 91321
rect 1258 90567 22141 90592
rect 1258 89753 198662 90567
rect 1258 89728 10493 89753
rect 1258 88999 36520 89024
rect 1258 88185 198662 88999
rect 1258 88160 8925 88185
rect 1258 87431 33901 87456
rect 1258 86617 198662 87431
rect 1258 86592 18152 86617
rect 1258 85863 10717 85888
rect 1258 85049 198662 85863
rect 1258 85024 22253 85049
rect 1258 84295 28301 84320
rect 1258 83481 198662 84295
rect 1258 83456 26509 83481
rect 1258 82727 14077 82752
rect 1258 81913 198662 82727
rect 1258 81888 16429 81913
rect 1258 81159 20237 81184
rect 1258 80345 198662 81159
rect 1258 80320 15757 80345
rect 1258 79591 34952 79616
rect 1258 78777 198662 79591
rect 1258 78752 18669 78777
rect 1258 78023 28301 78048
rect 1258 77209 198662 78023
rect 1258 77184 18669 77209
rect 1258 76455 28077 76480
rect 1258 75641 198662 76455
rect 1258 75616 39725 75641
rect 1258 74887 33901 74912
rect 1258 74073 198662 74887
rect 1258 74048 32893 74073
rect 1258 73319 21245 73344
rect 1258 72505 198662 73319
rect 1258 72480 15981 72505
rect 1258 71751 21021 71776
rect 1258 70937 198662 71751
rect 1258 70912 16205 70937
rect 1258 70183 30429 70208
rect 1258 69369 198662 70183
rect 1258 69344 33160 69369
rect 1258 68615 52941 68640
rect 1258 67801 198662 68615
rect 1258 67776 18669 67801
rect 1258 67047 18221 67072
rect 1258 66233 198662 67047
rect 1258 66208 43457 66233
rect 1258 65479 14749 65504
rect 1258 64665 198662 65479
rect 1258 64640 23597 64665
rect 1258 63911 15800 63936
rect 1258 63097 198662 63911
rect 1258 63072 31437 63097
rect 1258 62343 63057 62368
rect 1258 61529 198662 62343
rect 1258 61504 24269 61529
rect 1258 60775 21245 60800
rect 1258 59961 198662 60775
rect 1258 59936 17325 59961
rect 1258 59207 43787 59232
rect 1258 58393 198662 59207
rect 1258 58368 156942 58393
rect 1258 57639 14749 57664
rect 1258 56825 198662 57639
rect 1258 56800 30129 56825
rect 1258 56071 14749 56096
rect 1258 55257 198662 56071
rect 1258 55232 40433 55257
rect 1258 54503 14413 54528
rect 1258 53689 198662 54503
rect 1258 53664 40545 53689
rect 1258 52935 68061 52960
rect 1258 52121 198662 52935
rect 1258 52096 38872 52121
rect 1258 51367 13069 51392
rect 1258 50553 198662 51367
rect 1258 50528 40097 50553
rect 1258 49799 43533 49824
rect 1258 48985 198662 49799
rect 1258 48960 26285 48985
rect 1258 48231 11725 48256
rect 1258 47417 198662 48231
rect 1258 47392 10829 47417
rect 1258 46663 26397 46688
rect 1258 45849 198662 46663
rect 1258 45824 37821 45849
rect 1258 45095 20237 45120
rect 1258 44281 198662 45095
rect 1258 44256 14301 44281
rect 1258 43527 19789 43552
rect 1258 42713 198662 43527
rect 1258 42688 14301 42713
rect 1258 41959 20013 41984
rect 1258 41145 198662 41959
rect 1258 41120 55965 41145
rect 1258 40391 84568 40416
rect 1258 39577 198662 40391
rect 1258 39552 39165 39577
rect 1258 38823 38269 38848
rect 1258 38009 198662 38823
rect 1258 37984 15421 38009
rect 1258 37255 28232 37280
rect 1258 36441 198662 37255
rect 1258 36416 50029 36441
rect 1258 35687 13517 35712
rect 1258 34873 198662 35687
rect 1258 34848 34833 34873
rect 1258 34119 12621 34144
rect 1258 33305 198662 34119
rect 1258 33280 39389 33305
rect 1258 32551 12845 32576
rect 1258 31737 198662 32551
rect 1258 31712 32593 31737
rect 1258 30983 18221 31008
rect 1258 30169 198662 30983
rect 1258 30144 16653 30169
rect 1258 29415 27560 29440
rect 1258 28601 198662 29415
rect 1258 28576 65640 28601
rect 1258 27847 14189 27872
rect 1258 27033 198662 27847
rect 1258 27008 32145 27033
rect 1258 26279 14637 26304
rect 1258 25465 198662 26279
rect 1258 25440 22141 25465
rect 1258 24711 53949 24736
rect 1258 23897 198662 24711
rect 1258 23872 26509 23897
rect 1258 23143 43197 23168
rect 1258 22329 198662 23143
rect 1258 22304 15645 22329
rect 1258 21575 41741 21600
rect 1258 20761 198662 21575
rect 1258 20736 15757 20761
rect 1258 20007 22141 20032
rect 1258 19193 198662 20007
rect 1258 19168 24829 19193
rect 1258 18439 21245 18464
rect 1258 17625 198662 18439
rect 1258 17600 26776 17625
rect 1258 16871 28973 16896
rect 1258 16057 198662 16871
rect 1258 16032 31549 16057
rect 1258 15303 38760 15328
rect 1258 14489 198662 15303
rect 1258 14464 49581 14489
rect 1258 13735 35469 13760
rect 1258 12921 198662 13735
rect 1258 12896 53501 12921
rect 1258 12167 43197 12192
rect 1258 11353 198662 12167
rect 1258 11328 34349 11353
rect 1258 10599 60557 10624
rect 1258 9785 198662 10599
rect 1258 9760 57869 9785
rect 1258 9031 36925 9056
rect 1258 8217 198662 9031
rect 1258 8192 37821 8217
rect 1258 7463 51709 7488
rect 1258 6649 198662 7463
rect 1258 6624 42189 6649
rect 1258 5895 51485 5920
rect 1258 5081 198662 5895
rect 1258 5056 39165 5081
rect 1258 4327 42525 4352
rect 1258 3513 198662 4327
rect 1258 3488 133064 3513
<< pwell >>
rect 1258 195648 198662 196352
rect 1258 194080 198662 194784
rect 1258 192512 198662 193216
rect 1258 190944 198662 191648
rect 1258 189376 198662 190080
rect 1258 187808 198662 188512
rect 1258 186240 198662 186944
rect 1258 184672 198662 185376
rect 1258 183104 198662 183808
rect 1258 181536 198662 182240
rect 1258 179968 198662 180672
rect 1258 178400 198662 179104
rect 1258 176832 198662 177536
rect 1258 175264 198662 175968
rect 1258 173696 198662 174400
rect 1258 172128 198662 172832
rect 1258 170560 198662 171264
rect 1258 168992 198662 169696
rect 1258 167424 198662 168128
rect 1258 165856 198662 166560
rect 1258 164288 198662 164992
rect 1258 162720 198662 163424
rect 1258 161152 198662 161856
rect 1258 159584 198662 160288
rect 1258 158016 198662 158720
rect 1258 156448 198662 157152
rect 1258 154880 198662 155584
rect 1258 153312 198662 154016
rect 1258 151744 198662 152448
rect 1258 150176 198662 150880
rect 1258 148608 198662 149312
rect 1258 147040 198662 147744
rect 1258 145472 198662 146176
rect 1258 143904 198662 144608
rect 1258 142336 198662 143040
rect 1258 140768 198662 141472
rect 1258 139200 198662 139904
rect 1258 137632 198662 138336
rect 1258 136064 198662 136768
rect 1258 134496 198662 135200
rect 1258 132928 198662 133632
rect 1258 131360 198662 132064
rect 1258 129792 198662 130496
rect 1258 128224 198662 128928
rect 1258 126656 198662 127360
rect 1258 125088 198662 125792
rect 1258 123520 198662 124224
rect 1258 121952 198662 122656
rect 1258 120384 198662 121088
rect 1258 118816 198662 119520
rect 1258 117248 198662 117952
rect 1258 115680 198662 116384
rect 1258 114112 198662 114816
rect 1258 112544 198662 113248
rect 1258 110976 198662 111680
rect 1258 109408 198662 110112
rect 1258 107840 198662 108544
rect 1258 106272 198662 106976
rect 1258 104704 198662 105408
rect 1258 103136 198662 103840
rect 1258 101568 198662 102272
rect 1258 100000 198662 100704
rect 1258 98432 198662 99136
rect 1258 96864 198662 97568
rect 1258 95296 198662 96000
rect 1258 93728 198662 94432
rect 1258 92160 198662 92864
rect 1258 90592 198662 91296
rect 1258 89024 198662 89728
rect 1258 87456 198662 88160
rect 1258 85888 198662 86592
rect 1258 84320 198662 85024
rect 1258 82752 198662 83456
rect 1258 81184 198662 81888
rect 1258 79616 198662 80320
rect 1258 78048 198662 78752
rect 1258 76480 198662 77184
rect 1258 74912 198662 75616
rect 1258 73344 198662 74048
rect 1258 71776 198662 72480
rect 1258 70208 198662 70912
rect 1258 68640 198662 69344
rect 1258 67072 198662 67776
rect 1258 65504 198662 66208
rect 1258 63936 198662 64640
rect 1258 62368 198662 63072
rect 1258 60800 198662 61504
rect 1258 59232 198662 59936
rect 1258 57664 198662 58368
rect 1258 56096 198662 56800
rect 1258 54528 198662 55232
rect 1258 52960 198662 53664
rect 1258 51392 198662 52096
rect 1258 49824 198662 50528
rect 1258 48256 198662 48960
rect 1258 46688 198662 47392
rect 1258 45120 198662 45824
rect 1258 43552 198662 44256
rect 1258 41984 198662 42688
rect 1258 40416 198662 41120
rect 1258 38848 198662 39552
rect 1258 37280 198662 37984
rect 1258 35712 198662 36416
rect 1258 34144 198662 34848
rect 1258 32576 198662 33280
rect 1258 31008 198662 31712
rect 1258 29440 198662 30144
rect 1258 27872 198662 28576
rect 1258 26304 198662 27008
rect 1258 24736 198662 25440
rect 1258 23168 198662 23872
rect 1258 21600 198662 22304
rect 1258 20032 198662 20736
rect 1258 18464 198662 19168
rect 1258 16896 198662 17600
rect 1258 15328 198662 16032
rect 1258 13760 198662 14464
rect 1258 12192 198662 12896
rect 1258 10624 198662 11328
rect 1258 9056 198662 9760
rect 1258 7488 198662 8192
rect 1258 5920 198662 6624
rect 1258 4352 198662 5056
rect 1258 3050 198662 3488
<< obsm1 >>
rect 1344 3076 198576 196844
<< metal2 >>
rect 5824 199200 5936 200000
rect 7616 199200 7728 200000
rect 9408 199200 9520 200000
rect 11200 199200 11312 200000
rect 12992 199200 13104 200000
rect 14784 199200 14896 200000
rect 16576 199200 16688 200000
rect 18368 199200 18480 200000
rect 20160 199200 20272 200000
rect 21952 199200 22064 200000
rect 23744 199200 23856 200000
rect 25536 199200 25648 200000
rect 27328 199200 27440 200000
rect 29120 199200 29232 200000
rect 30912 199200 31024 200000
rect 32704 199200 32816 200000
rect 34496 199200 34608 200000
rect 36288 199200 36400 200000
rect 38080 199200 38192 200000
rect 39872 199200 39984 200000
rect 41664 199200 41776 200000
rect 43456 199200 43568 200000
rect 45248 199200 45360 200000
rect 47040 199200 47152 200000
rect 48832 199200 48944 200000
rect 50624 199200 50736 200000
rect 52416 199200 52528 200000
rect 54208 199200 54320 200000
rect 56000 199200 56112 200000
rect 57792 199200 57904 200000
rect 59584 199200 59696 200000
rect 61376 199200 61488 200000
rect 63168 199200 63280 200000
rect 64960 199200 65072 200000
rect 66752 199200 66864 200000
rect 68544 199200 68656 200000
rect 70336 199200 70448 200000
rect 72128 199200 72240 200000
rect 73920 199200 74032 200000
rect 75712 199200 75824 200000
rect 77504 199200 77616 200000
rect 79296 199200 79408 200000
rect 81088 199200 81200 200000
rect 82880 199200 82992 200000
rect 84672 199200 84784 200000
rect 86464 199200 86576 200000
rect 88256 199200 88368 200000
rect 90048 199200 90160 200000
rect 91840 199200 91952 200000
rect 93632 199200 93744 200000
rect 95424 199200 95536 200000
rect 97216 199200 97328 200000
rect 99008 199200 99120 200000
rect 100800 199200 100912 200000
rect 102592 199200 102704 200000
rect 104384 199200 104496 200000
rect 106176 199200 106288 200000
rect 107968 199200 108080 200000
rect 109760 199200 109872 200000
rect 111552 199200 111664 200000
rect 113344 199200 113456 200000
rect 115136 199200 115248 200000
rect 116928 199200 117040 200000
rect 118720 199200 118832 200000
rect 120512 199200 120624 200000
rect 122304 199200 122416 200000
rect 124096 199200 124208 200000
rect 125888 199200 126000 200000
rect 127680 199200 127792 200000
rect 129472 199200 129584 200000
rect 131264 199200 131376 200000
rect 133056 199200 133168 200000
rect 134848 199200 134960 200000
rect 136640 199200 136752 200000
rect 138432 199200 138544 200000
rect 140224 199200 140336 200000
rect 142016 199200 142128 200000
rect 143808 199200 143920 200000
rect 145600 199200 145712 200000
rect 147392 199200 147504 200000
rect 149184 199200 149296 200000
rect 150976 199200 151088 200000
rect 152768 199200 152880 200000
rect 154560 199200 154672 200000
rect 156352 199200 156464 200000
rect 158144 199200 158256 200000
rect 159936 199200 160048 200000
rect 161728 199200 161840 200000
rect 163520 199200 163632 200000
rect 165312 199200 165424 200000
rect 167104 199200 167216 200000
rect 168896 199200 169008 200000
rect 170688 199200 170800 200000
rect 172480 199200 172592 200000
rect 174272 199200 174384 200000
rect 176064 199200 176176 200000
rect 177856 199200 177968 200000
rect 179648 199200 179760 200000
rect 181440 199200 181552 200000
rect 183232 199200 183344 200000
rect 185024 199200 185136 200000
rect 186816 199200 186928 200000
rect 188608 199200 188720 200000
rect 190400 199200 190512 200000
rect 192192 199200 192304 200000
rect 193984 199200 194096 200000
rect 3136 0 3248 800
rect 5152 0 5264 800
rect 7168 0 7280 800
rect 9184 0 9296 800
rect 11200 0 11312 800
rect 13216 0 13328 800
rect 15232 0 15344 800
rect 17248 0 17360 800
rect 19264 0 19376 800
rect 21280 0 21392 800
rect 23296 0 23408 800
rect 25312 0 25424 800
rect 27328 0 27440 800
rect 29344 0 29456 800
rect 31360 0 31472 800
rect 33376 0 33488 800
rect 35392 0 35504 800
rect 37408 0 37520 800
rect 39424 0 39536 800
rect 41440 0 41552 800
rect 43456 0 43568 800
rect 45472 0 45584 800
rect 47488 0 47600 800
rect 49504 0 49616 800
rect 51520 0 51632 800
rect 53536 0 53648 800
rect 55552 0 55664 800
rect 57568 0 57680 800
rect 59584 0 59696 800
rect 61600 0 61712 800
rect 63616 0 63728 800
rect 65632 0 65744 800
rect 67648 0 67760 800
rect 69664 0 69776 800
rect 71680 0 71792 800
rect 73696 0 73808 800
rect 75712 0 75824 800
rect 77728 0 77840 800
rect 79744 0 79856 800
rect 81760 0 81872 800
rect 83776 0 83888 800
rect 85792 0 85904 800
rect 87808 0 87920 800
rect 89824 0 89936 800
rect 91840 0 91952 800
rect 93856 0 93968 800
rect 95872 0 95984 800
rect 97888 0 98000 800
rect 99904 0 100016 800
rect 101920 0 102032 800
rect 103936 0 104048 800
rect 105952 0 106064 800
rect 107968 0 108080 800
rect 109984 0 110096 800
rect 112000 0 112112 800
rect 114016 0 114128 800
rect 116032 0 116144 800
rect 118048 0 118160 800
rect 120064 0 120176 800
rect 122080 0 122192 800
rect 124096 0 124208 800
rect 126112 0 126224 800
rect 128128 0 128240 800
rect 130144 0 130256 800
rect 132160 0 132272 800
rect 134176 0 134288 800
rect 136192 0 136304 800
rect 138208 0 138320 800
rect 140224 0 140336 800
rect 142240 0 142352 800
rect 144256 0 144368 800
rect 146272 0 146384 800
rect 148288 0 148400 800
rect 150304 0 150416 800
rect 152320 0 152432 800
rect 154336 0 154448 800
rect 156352 0 156464 800
rect 158368 0 158480 800
rect 160384 0 160496 800
rect 162400 0 162512 800
rect 164416 0 164528 800
rect 166432 0 166544 800
rect 168448 0 168560 800
rect 170464 0 170576 800
rect 172480 0 172592 800
rect 174496 0 174608 800
rect 176512 0 176624 800
rect 178528 0 178640 800
rect 180544 0 180656 800
rect 182560 0 182672 800
rect 184576 0 184688 800
rect 186592 0 186704 800
rect 188608 0 188720 800
rect 190624 0 190736 800
rect 192640 0 192752 800
rect 194656 0 194768 800
rect 196672 0 196784 800
<< obsm2 >>
rect 1596 199140 5764 199332
rect 5996 199140 7556 199332
rect 7788 199140 9348 199332
rect 9580 199140 11140 199332
rect 11372 199140 12932 199332
rect 13164 199140 14724 199332
rect 14956 199140 16516 199332
rect 16748 199140 18308 199332
rect 18540 199140 20100 199332
rect 20332 199140 21892 199332
rect 22124 199140 23684 199332
rect 23916 199140 25476 199332
rect 25708 199140 27268 199332
rect 27500 199140 29060 199332
rect 29292 199140 30852 199332
rect 31084 199140 32644 199332
rect 32876 199140 34436 199332
rect 34668 199140 36228 199332
rect 36460 199140 38020 199332
rect 38252 199140 39812 199332
rect 40044 199140 41604 199332
rect 41836 199140 43396 199332
rect 43628 199140 45188 199332
rect 45420 199140 46980 199332
rect 47212 199140 48772 199332
rect 49004 199140 50564 199332
rect 50796 199140 52356 199332
rect 52588 199140 54148 199332
rect 54380 199140 55940 199332
rect 56172 199140 57732 199332
rect 57964 199140 59524 199332
rect 59756 199140 61316 199332
rect 61548 199140 63108 199332
rect 63340 199140 64900 199332
rect 65132 199140 66692 199332
rect 66924 199140 68484 199332
rect 68716 199140 70276 199332
rect 70508 199140 72068 199332
rect 72300 199140 73860 199332
rect 74092 199140 75652 199332
rect 75884 199140 77444 199332
rect 77676 199140 79236 199332
rect 79468 199140 81028 199332
rect 81260 199140 82820 199332
rect 83052 199140 84612 199332
rect 84844 199140 86404 199332
rect 86636 199140 88196 199332
rect 88428 199140 89988 199332
rect 90220 199140 91780 199332
rect 92012 199140 93572 199332
rect 93804 199140 95364 199332
rect 95596 199140 97156 199332
rect 97388 199140 98948 199332
rect 99180 199140 100740 199332
rect 100972 199140 102532 199332
rect 102764 199140 104324 199332
rect 104556 199140 106116 199332
rect 106348 199140 107908 199332
rect 108140 199140 109700 199332
rect 109932 199140 111492 199332
rect 111724 199140 113284 199332
rect 113516 199140 115076 199332
rect 115308 199140 116868 199332
rect 117100 199140 118660 199332
rect 118892 199140 120452 199332
rect 120684 199140 122244 199332
rect 122476 199140 124036 199332
rect 124268 199140 125828 199332
rect 126060 199140 127620 199332
rect 127852 199140 129412 199332
rect 129644 199140 131204 199332
rect 131436 199140 132996 199332
rect 133228 199140 134788 199332
rect 135020 199140 136580 199332
rect 136812 199140 138372 199332
rect 138604 199140 140164 199332
rect 140396 199140 141956 199332
rect 142188 199140 143748 199332
rect 143980 199140 145540 199332
rect 145772 199140 147332 199332
rect 147564 199140 149124 199332
rect 149356 199140 150916 199332
rect 151148 199140 152708 199332
rect 152940 199140 154500 199332
rect 154732 199140 156292 199332
rect 156524 199140 158084 199332
rect 158316 199140 159876 199332
rect 160108 199140 161668 199332
rect 161900 199140 163460 199332
rect 163692 199140 165252 199332
rect 165484 199140 167044 199332
rect 167276 199140 168836 199332
rect 169068 199140 170628 199332
rect 170860 199140 172420 199332
rect 172652 199140 174212 199332
rect 174444 199140 176004 199332
rect 176236 199140 177796 199332
rect 178028 199140 179588 199332
rect 179820 199140 181380 199332
rect 181612 199140 183172 199332
rect 183404 199140 184964 199332
rect 185196 199140 186756 199332
rect 186988 199140 188548 199332
rect 188780 199140 190340 199332
rect 190572 199140 192132 199332
rect 192364 199140 193924 199332
rect 194156 199140 198436 199332
rect 1596 860 198436 199140
rect 1596 466 3076 860
rect 3308 466 5092 860
rect 5324 466 7108 860
rect 7340 466 9124 860
rect 9356 466 11140 860
rect 11372 466 13156 860
rect 13388 466 15172 860
rect 15404 466 17188 860
rect 17420 466 19204 860
rect 19436 466 21220 860
rect 21452 466 23236 860
rect 23468 466 25252 860
rect 25484 466 27268 860
rect 27500 466 29284 860
rect 29516 466 31300 860
rect 31532 466 33316 860
rect 33548 466 35332 860
rect 35564 466 37348 860
rect 37580 466 39364 860
rect 39596 466 41380 860
rect 41612 466 43396 860
rect 43628 466 45412 860
rect 45644 466 47428 860
rect 47660 466 49444 860
rect 49676 466 51460 860
rect 51692 466 53476 860
rect 53708 466 55492 860
rect 55724 466 57508 860
rect 57740 466 59524 860
rect 59756 466 61540 860
rect 61772 466 63556 860
rect 63788 466 65572 860
rect 65804 466 67588 860
rect 67820 466 69604 860
rect 69836 466 71620 860
rect 71852 466 73636 860
rect 73868 466 75652 860
rect 75884 466 77668 860
rect 77900 466 79684 860
rect 79916 466 81700 860
rect 81932 466 83716 860
rect 83948 466 85732 860
rect 85964 466 87748 860
rect 87980 466 89764 860
rect 89996 466 91780 860
rect 92012 466 93796 860
rect 94028 466 95812 860
rect 96044 466 97828 860
rect 98060 466 99844 860
rect 100076 466 101860 860
rect 102092 466 103876 860
rect 104108 466 105892 860
rect 106124 466 107908 860
rect 108140 466 109924 860
rect 110156 466 111940 860
rect 112172 466 113956 860
rect 114188 466 115972 860
rect 116204 466 117988 860
rect 118220 466 120004 860
rect 120236 466 122020 860
rect 122252 466 124036 860
rect 124268 466 126052 860
rect 126284 466 128068 860
rect 128300 466 130084 860
rect 130316 466 132100 860
rect 132332 466 134116 860
rect 134348 466 136132 860
rect 136364 466 138148 860
rect 138380 466 140164 860
rect 140396 466 142180 860
rect 142412 466 144196 860
rect 144428 466 146212 860
rect 146444 466 148228 860
rect 148460 466 150244 860
rect 150476 466 152260 860
rect 152492 466 154276 860
rect 154508 466 156292 860
rect 156524 466 158308 860
rect 158540 466 160324 860
rect 160556 466 162340 860
rect 162572 466 164356 860
rect 164588 466 166372 860
rect 166604 466 168388 860
rect 168620 466 170404 860
rect 170636 466 172420 860
rect 172652 466 174436 860
rect 174668 466 176452 860
rect 176684 466 178468 860
rect 178700 466 180484 860
rect 180716 466 182500 860
rect 182732 466 184516 860
rect 184748 466 186532 860
rect 186764 466 188548 860
rect 188780 466 190564 860
rect 190796 466 192580 860
rect 192812 466 194596 860
rect 194828 466 196612 860
rect 196844 466 198436 860
<< obsm3 >>
rect 1586 476 198446 198996
<< metal4 >>
rect 4448 3076 4768 196844
rect 19808 3076 20128 196844
rect 35168 3076 35488 196844
rect 50528 3076 50848 196844
rect 65888 3076 66208 196844
rect 81248 3076 81568 196844
rect 96608 3076 96928 196844
rect 111968 3076 112288 196844
rect 127328 3076 127648 196844
rect 142688 3076 143008 196844
rect 158048 3076 158368 196844
rect 173408 3076 173728 196844
rect 188768 3076 189088 196844
<< obsm4 >>
rect 14924 3016 19748 196206
rect 20188 3016 35108 196206
rect 35548 3016 50468 196206
rect 50908 3016 65828 196206
rect 66268 3016 81188 196206
rect 81628 3016 96548 196206
rect 96988 3016 111908 196206
rect 112348 3016 127268 196206
rect 127708 3016 142628 196206
rect 143068 3016 157988 196206
rect 158428 3016 173348 196206
rect 173788 3016 188708 196206
rect 189148 3016 191044 196206
rect 14924 578 191044 3016
<< labels >>
rlabel metal2 s 3136 0 3248 800 6 clk
port 1 nsew signal input
rlabel metal2 s 5152 0 5264 800 6 inst[0]
port 2 nsew signal input
rlabel metal2 s 25312 0 25424 800 6 inst[10]
port 3 nsew signal input
rlabel metal2 s 27328 0 27440 800 6 inst[11]
port 4 nsew signal input
rlabel metal2 s 29344 0 29456 800 6 inst[12]
port 5 nsew signal input
rlabel metal2 s 31360 0 31472 800 6 inst[13]
port 6 nsew signal input
rlabel metal2 s 33376 0 33488 800 6 inst[14]
port 7 nsew signal input
rlabel metal2 s 35392 0 35504 800 6 inst[15]
port 8 nsew signal input
rlabel metal2 s 37408 0 37520 800 6 inst[16]
port 9 nsew signal input
rlabel metal2 s 39424 0 39536 800 6 inst[17]
port 10 nsew signal input
rlabel metal2 s 41440 0 41552 800 6 inst[18]
port 11 nsew signal input
rlabel metal2 s 43456 0 43568 800 6 inst[19]
port 12 nsew signal input
rlabel metal2 s 7168 0 7280 800 6 inst[1]
port 13 nsew signal input
rlabel metal2 s 45472 0 45584 800 6 inst[20]
port 14 nsew signal input
rlabel metal2 s 47488 0 47600 800 6 inst[21]
port 15 nsew signal input
rlabel metal2 s 49504 0 49616 800 6 inst[22]
port 16 nsew signal input
rlabel metal2 s 51520 0 51632 800 6 inst[23]
port 17 nsew signal input
rlabel metal2 s 53536 0 53648 800 6 inst[24]
port 18 nsew signal input
rlabel metal2 s 55552 0 55664 800 6 inst[25]
port 19 nsew signal input
rlabel metal2 s 57568 0 57680 800 6 inst[26]
port 20 nsew signal input
rlabel metal2 s 59584 0 59696 800 6 inst[27]
port 21 nsew signal input
rlabel metal2 s 61600 0 61712 800 6 inst[28]
port 22 nsew signal input
rlabel metal2 s 63616 0 63728 800 6 inst[29]
port 23 nsew signal input
rlabel metal2 s 9184 0 9296 800 6 inst[2]
port 24 nsew signal input
rlabel metal2 s 65632 0 65744 800 6 inst[30]
port 25 nsew signal input
rlabel metal2 s 67648 0 67760 800 6 inst[31]
port 26 nsew signal input
rlabel metal2 s 11200 0 11312 800 6 inst[3]
port 27 nsew signal input
rlabel metal2 s 13216 0 13328 800 6 inst[4]
port 28 nsew signal input
rlabel metal2 s 15232 0 15344 800 6 inst[5]
port 29 nsew signal input
rlabel metal2 s 17248 0 17360 800 6 inst[6]
port 30 nsew signal input
rlabel metal2 s 19264 0 19376 800 6 inst[7]
port 31 nsew signal input
rlabel metal2 s 21280 0 21392 800 6 inst[8]
port 32 nsew signal input
rlabel metal2 s 23296 0 23408 800 6 inst[9]
port 33 nsew signal input
rlabel metal2 s 193984 199200 194096 200000 6 mem_addr[0]
port 34 nsew signal output
rlabel metal2 s 176064 199200 176176 200000 6 mem_addr[10]
port 35 nsew signal output
rlabel metal2 s 174272 199200 174384 200000 6 mem_addr[11]
port 36 nsew signal output
rlabel metal2 s 172480 199200 172592 200000 6 mem_addr[12]
port 37 nsew signal output
rlabel metal2 s 170688 199200 170800 200000 6 mem_addr[13]
port 38 nsew signal output
rlabel metal2 s 168896 199200 169008 200000 6 mem_addr[14]
port 39 nsew signal output
rlabel metal2 s 167104 199200 167216 200000 6 mem_addr[15]
port 40 nsew signal output
rlabel metal2 s 165312 199200 165424 200000 6 mem_addr[16]
port 41 nsew signal output
rlabel metal2 s 163520 199200 163632 200000 6 mem_addr[17]
port 42 nsew signal output
rlabel metal2 s 161728 199200 161840 200000 6 mem_addr[18]
port 43 nsew signal output
rlabel metal2 s 159936 199200 160048 200000 6 mem_addr[19]
port 44 nsew signal output
rlabel metal2 s 192192 199200 192304 200000 6 mem_addr[1]
port 45 nsew signal output
rlabel metal2 s 158144 199200 158256 200000 6 mem_addr[20]
port 46 nsew signal output
rlabel metal2 s 156352 199200 156464 200000 6 mem_addr[21]
port 47 nsew signal output
rlabel metal2 s 154560 199200 154672 200000 6 mem_addr[22]
port 48 nsew signal output
rlabel metal2 s 152768 199200 152880 200000 6 mem_addr[23]
port 49 nsew signal output
rlabel metal2 s 150976 199200 151088 200000 6 mem_addr[24]
port 50 nsew signal output
rlabel metal2 s 149184 199200 149296 200000 6 mem_addr[25]
port 51 nsew signal output
rlabel metal2 s 147392 199200 147504 200000 6 mem_addr[26]
port 52 nsew signal output
rlabel metal2 s 145600 199200 145712 200000 6 mem_addr[27]
port 53 nsew signal output
rlabel metal2 s 143808 199200 143920 200000 6 mem_addr[28]
port 54 nsew signal output
rlabel metal2 s 142016 199200 142128 200000 6 mem_addr[29]
port 55 nsew signal output
rlabel metal2 s 190400 199200 190512 200000 6 mem_addr[2]
port 56 nsew signal output
rlabel metal2 s 140224 199200 140336 200000 6 mem_addr[30]
port 57 nsew signal output
rlabel metal2 s 138432 199200 138544 200000 6 mem_addr[31]
port 58 nsew signal output
rlabel metal2 s 188608 199200 188720 200000 6 mem_addr[3]
port 59 nsew signal output
rlabel metal2 s 186816 199200 186928 200000 6 mem_addr[4]
port 60 nsew signal output
rlabel metal2 s 185024 199200 185136 200000 6 mem_addr[5]
port 61 nsew signal output
rlabel metal2 s 183232 199200 183344 200000 6 mem_addr[6]
port 62 nsew signal output
rlabel metal2 s 181440 199200 181552 200000 6 mem_addr[7]
port 63 nsew signal output
rlabel metal2 s 179648 199200 179760 200000 6 mem_addr[8]
port 64 nsew signal output
rlabel metal2 s 177856 199200 177968 200000 6 mem_addr[9]
port 65 nsew signal output
rlabel metal2 s 127680 199200 127792 200000 6 mem_ld_dat[0]
port 66 nsew signal input
rlabel metal2 s 109760 199200 109872 200000 6 mem_ld_dat[10]
port 67 nsew signal input
rlabel metal2 s 107968 199200 108080 200000 6 mem_ld_dat[11]
port 68 nsew signal input
rlabel metal2 s 106176 199200 106288 200000 6 mem_ld_dat[12]
port 69 nsew signal input
rlabel metal2 s 104384 199200 104496 200000 6 mem_ld_dat[13]
port 70 nsew signal input
rlabel metal2 s 102592 199200 102704 200000 6 mem_ld_dat[14]
port 71 nsew signal input
rlabel metal2 s 100800 199200 100912 200000 6 mem_ld_dat[15]
port 72 nsew signal input
rlabel metal2 s 99008 199200 99120 200000 6 mem_ld_dat[16]
port 73 nsew signal input
rlabel metal2 s 97216 199200 97328 200000 6 mem_ld_dat[17]
port 74 nsew signal input
rlabel metal2 s 95424 199200 95536 200000 6 mem_ld_dat[18]
port 75 nsew signal input
rlabel metal2 s 93632 199200 93744 200000 6 mem_ld_dat[19]
port 76 nsew signal input
rlabel metal2 s 125888 199200 126000 200000 6 mem_ld_dat[1]
port 77 nsew signal input
rlabel metal2 s 91840 199200 91952 200000 6 mem_ld_dat[20]
port 78 nsew signal input
rlabel metal2 s 90048 199200 90160 200000 6 mem_ld_dat[21]
port 79 nsew signal input
rlabel metal2 s 88256 199200 88368 200000 6 mem_ld_dat[22]
port 80 nsew signal input
rlabel metal2 s 86464 199200 86576 200000 6 mem_ld_dat[23]
port 81 nsew signal input
rlabel metal2 s 84672 199200 84784 200000 6 mem_ld_dat[24]
port 82 nsew signal input
rlabel metal2 s 82880 199200 82992 200000 6 mem_ld_dat[25]
port 83 nsew signal input
rlabel metal2 s 81088 199200 81200 200000 6 mem_ld_dat[26]
port 84 nsew signal input
rlabel metal2 s 79296 199200 79408 200000 6 mem_ld_dat[27]
port 85 nsew signal input
rlabel metal2 s 77504 199200 77616 200000 6 mem_ld_dat[28]
port 86 nsew signal input
rlabel metal2 s 75712 199200 75824 200000 6 mem_ld_dat[29]
port 87 nsew signal input
rlabel metal2 s 124096 199200 124208 200000 6 mem_ld_dat[2]
port 88 nsew signal input
rlabel metal2 s 73920 199200 74032 200000 6 mem_ld_dat[30]
port 89 nsew signal input
rlabel metal2 s 72128 199200 72240 200000 6 mem_ld_dat[31]
port 90 nsew signal input
rlabel metal2 s 122304 199200 122416 200000 6 mem_ld_dat[3]
port 91 nsew signal input
rlabel metal2 s 120512 199200 120624 200000 6 mem_ld_dat[4]
port 92 nsew signal input
rlabel metal2 s 118720 199200 118832 200000 6 mem_ld_dat[5]
port 93 nsew signal input
rlabel metal2 s 116928 199200 117040 200000 6 mem_ld_dat[6]
port 94 nsew signal input
rlabel metal2 s 115136 199200 115248 200000 6 mem_ld_dat[7]
port 95 nsew signal input
rlabel metal2 s 113344 199200 113456 200000 6 mem_ld_dat[8]
port 96 nsew signal input
rlabel metal2 s 111552 199200 111664 200000 6 mem_ld_dat[9]
port 97 nsew signal input
rlabel metal2 s 136640 199200 136752 200000 6 mem_ld_en
port 98 nsew signal output
rlabel metal2 s 134848 199200 134960 200000 6 mem_ld_mask[0]
port 99 nsew signal output
rlabel metal2 s 133056 199200 133168 200000 6 mem_ld_mask[1]
port 100 nsew signal output
rlabel metal2 s 131264 199200 131376 200000 6 mem_ld_mask[2]
port 101 nsew signal output
rlabel metal2 s 129472 199200 129584 200000 6 mem_ld_mask[3]
port 102 nsew signal output
rlabel metal2 s 61376 199200 61488 200000 6 mem_st_dat[0]
port 103 nsew signal output
rlabel metal2 s 43456 199200 43568 200000 6 mem_st_dat[10]
port 104 nsew signal output
rlabel metal2 s 41664 199200 41776 200000 6 mem_st_dat[11]
port 105 nsew signal output
rlabel metal2 s 39872 199200 39984 200000 6 mem_st_dat[12]
port 106 nsew signal output
rlabel metal2 s 38080 199200 38192 200000 6 mem_st_dat[13]
port 107 nsew signal output
rlabel metal2 s 36288 199200 36400 200000 6 mem_st_dat[14]
port 108 nsew signal output
rlabel metal2 s 34496 199200 34608 200000 6 mem_st_dat[15]
port 109 nsew signal output
rlabel metal2 s 32704 199200 32816 200000 6 mem_st_dat[16]
port 110 nsew signal output
rlabel metal2 s 30912 199200 31024 200000 6 mem_st_dat[17]
port 111 nsew signal output
rlabel metal2 s 29120 199200 29232 200000 6 mem_st_dat[18]
port 112 nsew signal output
rlabel metal2 s 27328 199200 27440 200000 6 mem_st_dat[19]
port 113 nsew signal output
rlabel metal2 s 59584 199200 59696 200000 6 mem_st_dat[1]
port 114 nsew signal output
rlabel metal2 s 25536 199200 25648 200000 6 mem_st_dat[20]
port 115 nsew signal output
rlabel metal2 s 23744 199200 23856 200000 6 mem_st_dat[21]
port 116 nsew signal output
rlabel metal2 s 21952 199200 22064 200000 6 mem_st_dat[22]
port 117 nsew signal output
rlabel metal2 s 20160 199200 20272 200000 6 mem_st_dat[23]
port 118 nsew signal output
rlabel metal2 s 18368 199200 18480 200000 6 mem_st_dat[24]
port 119 nsew signal output
rlabel metal2 s 16576 199200 16688 200000 6 mem_st_dat[25]
port 120 nsew signal output
rlabel metal2 s 14784 199200 14896 200000 6 mem_st_dat[26]
port 121 nsew signal output
rlabel metal2 s 12992 199200 13104 200000 6 mem_st_dat[27]
port 122 nsew signal output
rlabel metal2 s 11200 199200 11312 200000 6 mem_st_dat[28]
port 123 nsew signal output
rlabel metal2 s 9408 199200 9520 200000 6 mem_st_dat[29]
port 124 nsew signal output
rlabel metal2 s 57792 199200 57904 200000 6 mem_st_dat[2]
port 125 nsew signal output
rlabel metal2 s 7616 199200 7728 200000 6 mem_st_dat[30]
port 126 nsew signal output
rlabel metal2 s 5824 199200 5936 200000 6 mem_st_dat[31]
port 127 nsew signal output
rlabel metal2 s 56000 199200 56112 200000 6 mem_st_dat[3]
port 128 nsew signal output
rlabel metal2 s 54208 199200 54320 200000 6 mem_st_dat[4]
port 129 nsew signal output
rlabel metal2 s 52416 199200 52528 200000 6 mem_st_dat[5]
port 130 nsew signal output
rlabel metal2 s 50624 199200 50736 200000 6 mem_st_dat[6]
port 131 nsew signal output
rlabel metal2 s 48832 199200 48944 200000 6 mem_st_dat[7]
port 132 nsew signal output
rlabel metal2 s 47040 199200 47152 200000 6 mem_st_dat[8]
port 133 nsew signal output
rlabel metal2 s 45248 199200 45360 200000 6 mem_st_dat[9]
port 134 nsew signal output
rlabel metal2 s 70336 199200 70448 200000 6 mem_st_en
port 135 nsew signal output
rlabel metal2 s 68544 199200 68656 200000 6 mem_st_mask[0]
port 136 nsew signal output
rlabel metal2 s 66752 199200 66864 200000 6 mem_st_mask[1]
port 137 nsew signal output
rlabel metal2 s 64960 199200 65072 200000 6 mem_st_mask[2]
port 138 nsew signal output
rlabel metal2 s 63168 199200 63280 200000 6 mem_st_mask[3]
port 139 nsew signal output
rlabel metal2 s 69664 0 69776 800 6 pc[0]
port 140 nsew signal input
rlabel metal2 s 89824 0 89936 800 6 pc[10]
port 141 nsew signal input
rlabel metal2 s 91840 0 91952 800 6 pc[11]
port 142 nsew signal input
rlabel metal2 s 93856 0 93968 800 6 pc[12]
port 143 nsew signal input
rlabel metal2 s 95872 0 95984 800 6 pc[13]
port 144 nsew signal input
rlabel metal2 s 97888 0 98000 800 6 pc[14]
port 145 nsew signal input
rlabel metal2 s 99904 0 100016 800 6 pc[15]
port 146 nsew signal input
rlabel metal2 s 101920 0 102032 800 6 pc[16]
port 147 nsew signal input
rlabel metal2 s 103936 0 104048 800 6 pc[17]
port 148 nsew signal input
rlabel metal2 s 105952 0 106064 800 6 pc[18]
port 149 nsew signal input
rlabel metal2 s 107968 0 108080 800 6 pc[19]
port 150 nsew signal input
rlabel metal2 s 71680 0 71792 800 6 pc[1]
port 151 nsew signal input
rlabel metal2 s 109984 0 110096 800 6 pc[20]
port 152 nsew signal input
rlabel metal2 s 112000 0 112112 800 6 pc[21]
port 153 nsew signal input
rlabel metal2 s 114016 0 114128 800 6 pc[22]
port 154 nsew signal input
rlabel metal2 s 116032 0 116144 800 6 pc[23]
port 155 nsew signal input
rlabel metal2 s 118048 0 118160 800 6 pc[24]
port 156 nsew signal input
rlabel metal2 s 120064 0 120176 800 6 pc[25]
port 157 nsew signal input
rlabel metal2 s 122080 0 122192 800 6 pc[26]
port 158 nsew signal input
rlabel metal2 s 124096 0 124208 800 6 pc[27]
port 159 nsew signal input
rlabel metal2 s 126112 0 126224 800 6 pc[28]
port 160 nsew signal input
rlabel metal2 s 128128 0 128240 800 6 pc[29]
port 161 nsew signal input
rlabel metal2 s 73696 0 73808 800 6 pc[2]
port 162 nsew signal input
rlabel metal2 s 130144 0 130256 800 6 pc[30]
port 163 nsew signal input
rlabel metal2 s 132160 0 132272 800 6 pc[31]
port 164 nsew signal input
rlabel metal2 s 75712 0 75824 800 6 pc[3]
port 165 nsew signal input
rlabel metal2 s 77728 0 77840 800 6 pc[4]
port 166 nsew signal input
rlabel metal2 s 79744 0 79856 800 6 pc[5]
port 167 nsew signal input
rlabel metal2 s 81760 0 81872 800 6 pc[6]
port 168 nsew signal input
rlabel metal2 s 83776 0 83888 800 6 pc[7]
port 169 nsew signal input
rlabel metal2 s 85792 0 85904 800 6 pc[8]
port 170 nsew signal input
rlabel metal2 s 87808 0 87920 800 6 pc[9]
port 171 nsew signal input
rlabel metal2 s 134176 0 134288 800 6 pc_next[0]
port 172 nsew signal output
rlabel metal2 s 154336 0 154448 800 6 pc_next[10]
port 173 nsew signal output
rlabel metal2 s 156352 0 156464 800 6 pc_next[11]
port 174 nsew signal output
rlabel metal2 s 158368 0 158480 800 6 pc_next[12]
port 175 nsew signal output
rlabel metal2 s 160384 0 160496 800 6 pc_next[13]
port 176 nsew signal output
rlabel metal2 s 162400 0 162512 800 6 pc_next[14]
port 177 nsew signal output
rlabel metal2 s 164416 0 164528 800 6 pc_next[15]
port 178 nsew signal output
rlabel metal2 s 166432 0 166544 800 6 pc_next[16]
port 179 nsew signal output
rlabel metal2 s 168448 0 168560 800 6 pc_next[17]
port 180 nsew signal output
rlabel metal2 s 170464 0 170576 800 6 pc_next[18]
port 181 nsew signal output
rlabel metal2 s 172480 0 172592 800 6 pc_next[19]
port 182 nsew signal output
rlabel metal2 s 136192 0 136304 800 6 pc_next[1]
port 183 nsew signal output
rlabel metal2 s 174496 0 174608 800 6 pc_next[20]
port 184 nsew signal output
rlabel metal2 s 176512 0 176624 800 6 pc_next[21]
port 185 nsew signal output
rlabel metal2 s 178528 0 178640 800 6 pc_next[22]
port 186 nsew signal output
rlabel metal2 s 180544 0 180656 800 6 pc_next[23]
port 187 nsew signal output
rlabel metal2 s 182560 0 182672 800 6 pc_next[24]
port 188 nsew signal output
rlabel metal2 s 184576 0 184688 800 6 pc_next[25]
port 189 nsew signal output
rlabel metal2 s 186592 0 186704 800 6 pc_next[26]
port 190 nsew signal output
rlabel metal2 s 188608 0 188720 800 6 pc_next[27]
port 191 nsew signal output
rlabel metal2 s 190624 0 190736 800 6 pc_next[28]
port 192 nsew signal output
rlabel metal2 s 192640 0 192752 800 6 pc_next[29]
port 193 nsew signal output
rlabel metal2 s 138208 0 138320 800 6 pc_next[2]
port 194 nsew signal output
rlabel metal2 s 194656 0 194768 800 6 pc_next[30]
port 195 nsew signal output
rlabel metal2 s 196672 0 196784 800 6 pc_next[31]
port 196 nsew signal output
rlabel metal2 s 140224 0 140336 800 6 pc_next[3]
port 197 nsew signal output
rlabel metal2 s 142240 0 142352 800 6 pc_next[4]
port 198 nsew signal output
rlabel metal2 s 144256 0 144368 800 6 pc_next[5]
port 199 nsew signal output
rlabel metal2 s 146272 0 146384 800 6 pc_next[6]
port 200 nsew signal output
rlabel metal2 s 148288 0 148400 800 6 pc_next[7]
port 201 nsew signal output
rlabel metal2 s 150304 0 150416 800 6 pc_next[8]
port 202 nsew signal output
rlabel metal2 s 152320 0 152432 800 6 pc_next[9]
port 203 nsew signal output
rlabel metal4 s 4448 3076 4768 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 196844 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 196844 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 196844 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 196844 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 196844 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 196844 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 196844 6 vss
port 205 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27399966
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/rv_core/runs/23_11_26_16_46/results/signoff/tinyrv.magic.gds
string GDS_START 559798
<< end >>

