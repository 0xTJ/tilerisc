magic
tech gf180mcuD
magscale 1 5
timestamp 1700489575
<< obsm1 >>
rect 672 855 279328 78889
<< metal2 >>
rect 3696 79600 3752 80000
rect 5824 79600 5880 80000
rect 7952 79600 8008 80000
rect 10080 79600 10136 80000
rect 12208 79600 12264 80000
rect 14336 79600 14392 80000
rect 16464 79600 16520 80000
rect 18592 79600 18648 80000
rect 20720 79600 20776 80000
rect 22848 79600 22904 80000
rect 24976 79600 25032 80000
rect 27104 79600 27160 80000
rect 29232 79600 29288 80000
rect 31360 79600 31416 80000
rect 33488 79600 33544 80000
rect 35616 79600 35672 80000
rect 37744 79600 37800 80000
rect 39872 79600 39928 80000
rect 42000 79600 42056 80000
rect 44128 79600 44184 80000
rect 46256 79600 46312 80000
rect 48384 79600 48440 80000
rect 50512 79600 50568 80000
rect 52640 79600 52696 80000
rect 54768 79600 54824 80000
rect 56896 79600 56952 80000
rect 59024 79600 59080 80000
rect 61152 79600 61208 80000
rect 63280 79600 63336 80000
rect 65408 79600 65464 80000
rect 67536 79600 67592 80000
rect 69664 79600 69720 80000
rect 71792 79600 71848 80000
rect 73920 79600 73976 80000
rect 76048 79600 76104 80000
rect 78176 79600 78232 80000
rect 80304 79600 80360 80000
rect 82432 79600 82488 80000
rect 84560 79600 84616 80000
rect 86688 79600 86744 80000
rect 88816 79600 88872 80000
rect 90944 79600 91000 80000
rect 93072 79600 93128 80000
rect 95200 79600 95256 80000
rect 97328 79600 97384 80000
rect 99456 79600 99512 80000
rect 101584 79600 101640 80000
rect 103712 79600 103768 80000
rect 105840 79600 105896 80000
rect 107968 79600 108024 80000
rect 110096 79600 110152 80000
rect 112224 79600 112280 80000
rect 114352 79600 114408 80000
rect 116480 79600 116536 80000
rect 118608 79600 118664 80000
rect 120736 79600 120792 80000
rect 122864 79600 122920 80000
rect 124992 79600 125048 80000
rect 127120 79600 127176 80000
rect 129248 79600 129304 80000
rect 131376 79600 131432 80000
rect 133504 79600 133560 80000
rect 135632 79600 135688 80000
rect 137760 79600 137816 80000
rect 139888 79600 139944 80000
rect 142016 79600 142072 80000
rect 144144 79600 144200 80000
rect 146272 79600 146328 80000
rect 148400 79600 148456 80000
rect 150528 79600 150584 80000
rect 152656 79600 152712 80000
rect 154784 79600 154840 80000
rect 156912 79600 156968 80000
rect 159040 79600 159096 80000
rect 161168 79600 161224 80000
rect 163296 79600 163352 80000
rect 165424 79600 165480 80000
rect 167552 79600 167608 80000
rect 169680 79600 169736 80000
rect 171808 79600 171864 80000
rect 173936 79600 173992 80000
rect 176064 79600 176120 80000
rect 178192 79600 178248 80000
rect 180320 79600 180376 80000
rect 182448 79600 182504 80000
rect 184576 79600 184632 80000
rect 186704 79600 186760 80000
rect 188832 79600 188888 80000
rect 190960 79600 191016 80000
rect 193088 79600 193144 80000
rect 195216 79600 195272 80000
rect 197344 79600 197400 80000
rect 199472 79600 199528 80000
rect 201600 79600 201656 80000
rect 203728 79600 203784 80000
rect 205856 79600 205912 80000
rect 207984 79600 208040 80000
rect 210112 79600 210168 80000
rect 212240 79600 212296 80000
rect 214368 79600 214424 80000
rect 216496 79600 216552 80000
rect 218624 79600 218680 80000
rect 220752 79600 220808 80000
rect 222880 79600 222936 80000
rect 225008 79600 225064 80000
rect 227136 79600 227192 80000
rect 229264 79600 229320 80000
rect 231392 79600 231448 80000
rect 233520 79600 233576 80000
rect 235648 79600 235704 80000
rect 237776 79600 237832 80000
rect 239904 79600 239960 80000
rect 242032 79600 242088 80000
rect 244160 79600 244216 80000
rect 246288 79600 246344 80000
rect 248416 79600 248472 80000
rect 250544 79600 250600 80000
rect 252672 79600 252728 80000
rect 254800 79600 254856 80000
rect 256928 79600 256984 80000
rect 259056 79600 259112 80000
rect 261184 79600 261240 80000
rect 263312 79600 263368 80000
rect 265440 79600 265496 80000
rect 267568 79600 267624 80000
rect 269696 79600 269752 80000
rect 271824 79600 271880 80000
rect 273952 79600 274008 80000
rect 276080 79600 276136 80000
rect 3472 0 3528 400
rect 3808 0 3864 400
rect 4144 0 4200 400
rect 4480 0 4536 400
rect 4816 0 4872 400
rect 5152 0 5208 400
rect 5488 0 5544 400
rect 5824 0 5880 400
rect 6160 0 6216 400
rect 6496 0 6552 400
rect 6832 0 6888 400
rect 7168 0 7224 400
rect 7504 0 7560 400
rect 7840 0 7896 400
rect 8176 0 8232 400
rect 8512 0 8568 400
rect 8848 0 8904 400
rect 9184 0 9240 400
rect 9520 0 9576 400
rect 9856 0 9912 400
rect 10192 0 10248 400
rect 10528 0 10584 400
rect 10864 0 10920 400
rect 11200 0 11256 400
rect 11536 0 11592 400
rect 11872 0 11928 400
rect 12208 0 12264 400
rect 12544 0 12600 400
rect 12880 0 12936 400
rect 13216 0 13272 400
rect 13552 0 13608 400
rect 13888 0 13944 400
rect 14224 0 14280 400
rect 14560 0 14616 400
rect 14896 0 14952 400
rect 15232 0 15288 400
rect 15568 0 15624 400
rect 15904 0 15960 400
rect 16240 0 16296 400
rect 16576 0 16632 400
rect 16912 0 16968 400
rect 17248 0 17304 400
rect 17584 0 17640 400
rect 17920 0 17976 400
rect 18256 0 18312 400
rect 18592 0 18648 400
rect 18928 0 18984 400
rect 19264 0 19320 400
rect 19600 0 19656 400
rect 19936 0 19992 400
rect 20272 0 20328 400
rect 20608 0 20664 400
rect 20944 0 21000 400
rect 21280 0 21336 400
rect 21616 0 21672 400
rect 21952 0 22008 400
rect 22288 0 22344 400
rect 22624 0 22680 400
rect 22960 0 23016 400
rect 23296 0 23352 400
rect 23632 0 23688 400
rect 23968 0 24024 400
rect 24304 0 24360 400
rect 24640 0 24696 400
rect 24976 0 25032 400
rect 25312 0 25368 400
rect 25648 0 25704 400
rect 25984 0 26040 400
rect 26320 0 26376 400
rect 26656 0 26712 400
rect 26992 0 27048 400
rect 27328 0 27384 400
rect 27664 0 27720 400
rect 28000 0 28056 400
rect 28336 0 28392 400
rect 28672 0 28728 400
rect 29008 0 29064 400
rect 29344 0 29400 400
rect 29680 0 29736 400
rect 30016 0 30072 400
rect 30352 0 30408 400
rect 30688 0 30744 400
rect 31024 0 31080 400
rect 31360 0 31416 400
rect 31696 0 31752 400
rect 32032 0 32088 400
rect 32368 0 32424 400
rect 32704 0 32760 400
rect 33040 0 33096 400
rect 33376 0 33432 400
rect 33712 0 33768 400
rect 34048 0 34104 400
rect 34384 0 34440 400
rect 34720 0 34776 400
rect 35056 0 35112 400
rect 35392 0 35448 400
rect 35728 0 35784 400
rect 36064 0 36120 400
rect 36400 0 36456 400
rect 36736 0 36792 400
rect 37072 0 37128 400
rect 37408 0 37464 400
rect 37744 0 37800 400
rect 38080 0 38136 400
rect 38416 0 38472 400
rect 38752 0 38808 400
rect 39088 0 39144 400
rect 39424 0 39480 400
rect 39760 0 39816 400
rect 40096 0 40152 400
rect 40432 0 40488 400
rect 40768 0 40824 400
rect 41104 0 41160 400
rect 41440 0 41496 400
rect 41776 0 41832 400
rect 42112 0 42168 400
rect 42448 0 42504 400
rect 42784 0 42840 400
rect 43120 0 43176 400
rect 43456 0 43512 400
rect 43792 0 43848 400
rect 44128 0 44184 400
rect 44464 0 44520 400
rect 44800 0 44856 400
rect 45136 0 45192 400
rect 45472 0 45528 400
rect 45808 0 45864 400
rect 46144 0 46200 400
rect 46480 0 46536 400
rect 46816 0 46872 400
rect 47152 0 47208 400
rect 47488 0 47544 400
rect 47824 0 47880 400
rect 48160 0 48216 400
rect 48496 0 48552 400
rect 48832 0 48888 400
rect 49168 0 49224 400
rect 49504 0 49560 400
rect 49840 0 49896 400
rect 50176 0 50232 400
rect 50512 0 50568 400
rect 50848 0 50904 400
rect 51184 0 51240 400
rect 51520 0 51576 400
rect 51856 0 51912 400
rect 52192 0 52248 400
rect 52528 0 52584 400
rect 52864 0 52920 400
rect 53200 0 53256 400
rect 53536 0 53592 400
rect 53872 0 53928 400
rect 54208 0 54264 400
rect 54544 0 54600 400
rect 54880 0 54936 400
rect 55216 0 55272 400
rect 55552 0 55608 400
rect 55888 0 55944 400
rect 56224 0 56280 400
rect 56560 0 56616 400
rect 56896 0 56952 400
rect 57232 0 57288 400
rect 57568 0 57624 400
rect 57904 0 57960 400
rect 58240 0 58296 400
rect 58576 0 58632 400
rect 58912 0 58968 400
rect 59248 0 59304 400
rect 59584 0 59640 400
rect 59920 0 59976 400
rect 60256 0 60312 400
rect 60592 0 60648 400
rect 60928 0 60984 400
rect 61264 0 61320 400
rect 61600 0 61656 400
rect 61936 0 61992 400
rect 62272 0 62328 400
rect 62608 0 62664 400
rect 62944 0 63000 400
rect 63280 0 63336 400
rect 63616 0 63672 400
rect 63952 0 64008 400
rect 64288 0 64344 400
rect 64624 0 64680 400
rect 64960 0 65016 400
rect 65296 0 65352 400
rect 65632 0 65688 400
rect 65968 0 66024 400
rect 66304 0 66360 400
rect 66640 0 66696 400
rect 66976 0 67032 400
rect 67312 0 67368 400
rect 67648 0 67704 400
rect 67984 0 68040 400
rect 68320 0 68376 400
rect 68656 0 68712 400
rect 68992 0 69048 400
rect 69328 0 69384 400
rect 69664 0 69720 400
rect 70000 0 70056 400
rect 70336 0 70392 400
rect 70672 0 70728 400
rect 71008 0 71064 400
rect 71344 0 71400 400
rect 71680 0 71736 400
rect 72016 0 72072 400
rect 72352 0 72408 400
rect 72688 0 72744 400
rect 73024 0 73080 400
rect 73360 0 73416 400
rect 73696 0 73752 400
rect 74032 0 74088 400
rect 74368 0 74424 400
rect 74704 0 74760 400
rect 75040 0 75096 400
rect 75376 0 75432 400
rect 75712 0 75768 400
rect 76048 0 76104 400
rect 76384 0 76440 400
rect 76720 0 76776 400
rect 77056 0 77112 400
rect 77392 0 77448 400
rect 77728 0 77784 400
rect 78064 0 78120 400
rect 78400 0 78456 400
rect 78736 0 78792 400
rect 79072 0 79128 400
rect 79408 0 79464 400
rect 79744 0 79800 400
rect 80080 0 80136 400
rect 80416 0 80472 400
rect 80752 0 80808 400
rect 81088 0 81144 400
rect 81424 0 81480 400
rect 81760 0 81816 400
rect 82096 0 82152 400
rect 82432 0 82488 400
rect 82768 0 82824 400
rect 83104 0 83160 400
rect 83440 0 83496 400
rect 83776 0 83832 400
rect 84112 0 84168 400
rect 84448 0 84504 400
rect 84784 0 84840 400
rect 85120 0 85176 400
rect 85456 0 85512 400
rect 85792 0 85848 400
rect 86128 0 86184 400
rect 86464 0 86520 400
rect 86800 0 86856 400
rect 87136 0 87192 400
rect 87472 0 87528 400
rect 87808 0 87864 400
rect 88144 0 88200 400
rect 88480 0 88536 400
rect 88816 0 88872 400
rect 89152 0 89208 400
rect 89488 0 89544 400
rect 89824 0 89880 400
rect 90160 0 90216 400
rect 90496 0 90552 400
rect 90832 0 90888 400
rect 91168 0 91224 400
rect 91504 0 91560 400
rect 91840 0 91896 400
rect 92176 0 92232 400
rect 92512 0 92568 400
rect 92848 0 92904 400
rect 93184 0 93240 400
rect 93520 0 93576 400
rect 93856 0 93912 400
rect 94192 0 94248 400
rect 94528 0 94584 400
rect 94864 0 94920 400
rect 95200 0 95256 400
rect 95536 0 95592 400
rect 95872 0 95928 400
rect 96208 0 96264 400
rect 96544 0 96600 400
rect 96880 0 96936 400
rect 97216 0 97272 400
rect 97552 0 97608 400
rect 97888 0 97944 400
rect 98224 0 98280 400
rect 98560 0 98616 400
rect 98896 0 98952 400
rect 99232 0 99288 400
rect 99568 0 99624 400
rect 99904 0 99960 400
rect 100240 0 100296 400
rect 100576 0 100632 400
rect 100912 0 100968 400
rect 101248 0 101304 400
rect 101584 0 101640 400
rect 101920 0 101976 400
rect 102256 0 102312 400
rect 102592 0 102648 400
rect 102928 0 102984 400
rect 103264 0 103320 400
rect 103600 0 103656 400
rect 103936 0 103992 400
rect 104272 0 104328 400
rect 104608 0 104664 400
rect 104944 0 105000 400
rect 105280 0 105336 400
rect 105616 0 105672 400
rect 105952 0 106008 400
rect 106288 0 106344 400
rect 106624 0 106680 400
rect 106960 0 107016 400
rect 107296 0 107352 400
rect 107632 0 107688 400
rect 107968 0 108024 400
rect 108304 0 108360 400
rect 108640 0 108696 400
rect 108976 0 109032 400
rect 109312 0 109368 400
rect 109648 0 109704 400
rect 109984 0 110040 400
rect 110320 0 110376 400
rect 110656 0 110712 400
rect 110992 0 111048 400
rect 111328 0 111384 400
rect 111664 0 111720 400
rect 112000 0 112056 400
rect 112336 0 112392 400
rect 112672 0 112728 400
rect 113008 0 113064 400
rect 113344 0 113400 400
rect 113680 0 113736 400
rect 114016 0 114072 400
rect 114352 0 114408 400
rect 114688 0 114744 400
rect 115024 0 115080 400
rect 115360 0 115416 400
rect 115696 0 115752 400
rect 116032 0 116088 400
rect 116368 0 116424 400
rect 116704 0 116760 400
rect 117040 0 117096 400
rect 117376 0 117432 400
rect 117712 0 117768 400
rect 118048 0 118104 400
rect 118384 0 118440 400
rect 118720 0 118776 400
rect 119056 0 119112 400
rect 119392 0 119448 400
rect 119728 0 119784 400
rect 120064 0 120120 400
rect 120400 0 120456 400
rect 120736 0 120792 400
rect 121072 0 121128 400
rect 121408 0 121464 400
rect 121744 0 121800 400
rect 122080 0 122136 400
rect 122416 0 122472 400
rect 122752 0 122808 400
rect 123088 0 123144 400
rect 123424 0 123480 400
rect 123760 0 123816 400
rect 124096 0 124152 400
rect 124432 0 124488 400
rect 124768 0 124824 400
rect 125104 0 125160 400
rect 125440 0 125496 400
rect 125776 0 125832 400
rect 126112 0 126168 400
rect 126448 0 126504 400
rect 126784 0 126840 400
rect 127120 0 127176 400
rect 127456 0 127512 400
rect 127792 0 127848 400
rect 128128 0 128184 400
rect 128464 0 128520 400
rect 128800 0 128856 400
rect 129136 0 129192 400
rect 129472 0 129528 400
rect 129808 0 129864 400
rect 130144 0 130200 400
rect 130480 0 130536 400
rect 130816 0 130872 400
rect 131152 0 131208 400
rect 131488 0 131544 400
rect 131824 0 131880 400
rect 132160 0 132216 400
rect 132496 0 132552 400
rect 132832 0 132888 400
rect 133168 0 133224 400
rect 133504 0 133560 400
rect 133840 0 133896 400
rect 134176 0 134232 400
rect 134512 0 134568 400
rect 134848 0 134904 400
rect 135184 0 135240 400
rect 135520 0 135576 400
rect 135856 0 135912 400
rect 136192 0 136248 400
rect 136528 0 136584 400
rect 136864 0 136920 400
rect 137200 0 137256 400
rect 137536 0 137592 400
rect 137872 0 137928 400
rect 138208 0 138264 400
rect 138544 0 138600 400
rect 138880 0 138936 400
rect 139216 0 139272 400
rect 139552 0 139608 400
rect 139888 0 139944 400
rect 140224 0 140280 400
rect 140560 0 140616 400
rect 140896 0 140952 400
rect 141232 0 141288 400
rect 141568 0 141624 400
rect 141904 0 141960 400
rect 142240 0 142296 400
rect 142576 0 142632 400
rect 142912 0 142968 400
rect 143248 0 143304 400
rect 143584 0 143640 400
rect 143920 0 143976 400
rect 144256 0 144312 400
rect 144592 0 144648 400
rect 144928 0 144984 400
rect 145264 0 145320 400
rect 145600 0 145656 400
rect 145936 0 145992 400
rect 146272 0 146328 400
rect 146608 0 146664 400
rect 146944 0 147000 400
rect 147280 0 147336 400
rect 147616 0 147672 400
rect 147952 0 148008 400
rect 148288 0 148344 400
rect 148624 0 148680 400
rect 148960 0 149016 400
rect 149296 0 149352 400
rect 149632 0 149688 400
rect 149968 0 150024 400
rect 150304 0 150360 400
rect 150640 0 150696 400
rect 150976 0 151032 400
rect 151312 0 151368 400
rect 151648 0 151704 400
rect 151984 0 152040 400
rect 152320 0 152376 400
rect 152656 0 152712 400
rect 152992 0 153048 400
rect 153328 0 153384 400
rect 153664 0 153720 400
rect 154000 0 154056 400
rect 154336 0 154392 400
rect 154672 0 154728 400
rect 155008 0 155064 400
rect 155344 0 155400 400
rect 155680 0 155736 400
rect 156016 0 156072 400
rect 156352 0 156408 400
rect 156688 0 156744 400
rect 157024 0 157080 400
rect 157360 0 157416 400
rect 157696 0 157752 400
rect 158032 0 158088 400
rect 158368 0 158424 400
rect 158704 0 158760 400
rect 159040 0 159096 400
rect 159376 0 159432 400
rect 159712 0 159768 400
rect 160048 0 160104 400
rect 160384 0 160440 400
rect 160720 0 160776 400
rect 161056 0 161112 400
rect 161392 0 161448 400
rect 161728 0 161784 400
rect 162064 0 162120 400
rect 162400 0 162456 400
rect 162736 0 162792 400
rect 163072 0 163128 400
rect 163408 0 163464 400
rect 163744 0 163800 400
rect 164080 0 164136 400
rect 164416 0 164472 400
rect 164752 0 164808 400
rect 165088 0 165144 400
rect 165424 0 165480 400
rect 165760 0 165816 400
rect 166096 0 166152 400
rect 166432 0 166488 400
rect 166768 0 166824 400
rect 167104 0 167160 400
rect 167440 0 167496 400
rect 167776 0 167832 400
rect 168112 0 168168 400
rect 168448 0 168504 400
rect 168784 0 168840 400
rect 169120 0 169176 400
rect 169456 0 169512 400
rect 169792 0 169848 400
rect 170128 0 170184 400
rect 170464 0 170520 400
rect 170800 0 170856 400
rect 171136 0 171192 400
rect 171472 0 171528 400
rect 171808 0 171864 400
rect 172144 0 172200 400
rect 172480 0 172536 400
rect 172816 0 172872 400
rect 173152 0 173208 400
rect 173488 0 173544 400
rect 173824 0 173880 400
rect 174160 0 174216 400
rect 174496 0 174552 400
rect 174832 0 174888 400
rect 175168 0 175224 400
rect 175504 0 175560 400
rect 175840 0 175896 400
rect 176176 0 176232 400
rect 176512 0 176568 400
rect 176848 0 176904 400
rect 177184 0 177240 400
rect 177520 0 177576 400
rect 177856 0 177912 400
rect 178192 0 178248 400
rect 178528 0 178584 400
rect 178864 0 178920 400
rect 179200 0 179256 400
rect 179536 0 179592 400
rect 179872 0 179928 400
rect 180208 0 180264 400
rect 180544 0 180600 400
rect 180880 0 180936 400
rect 181216 0 181272 400
rect 181552 0 181608 400
rect 181888 0 181944 400
rect 182224 0 182280 400
rect 182560 0 182616 400
rect 182896 0 182952 400
rect 183232 0 183288 400
rect 183568 0 183624 400
rect 183904 0 183960 400
rect 184240 0 184296 400
rect 184576 0 184632 400
rect 184912 0 184968 400
rect 185248 0 185304 400
rect 185584 0 185640 400
rect 185920 0 185976 400
rect 186256 0 186312 400
rect 186592 0 186648 400
rect 186928 0 186984 400
rect 187264 0 187320 400
rect 187600 0 187656 400
rect 187936 0 187992 400
rect 188272 0 188328 400
rect 188608 0 188664 400
rect 188944 0 189000 400
rect 189280 0 189336 400
rect 189616 0 189672 400
rect 189952 0 190008 400
rect 190288 0 190344 400
rect 190624 0 190680 400
rect 190960 0 191016 400
rect 191296 0 191352 400
rect 191632 0 191688 400
rect 191968 0 192024 400
rect 192304 0 192360 400
rect 192640 0 192696 400
rect 192976 0 193032 400
rect 193312 0 193368 400
rect 193648 0 193704 400
rect 193984 0 194040 400
rect 194320 0 194376 400
rect 194656 0 194712 400
rect 194992 0 195048 400
rect 195328 0 195384 400
rect 195664 0 195720 400
rect 196000 0 196056 400
rect 196336 0 196392 400
rect 196672 0 196728 400
rect 197008 0 197064 400
rect 197344 0 197400 400
rect 197680 0 197736 400
rect 198016 0 198072 400
rect 198352 0 198408 400
rect 198688 0 198744 400
rect 199024 0 199080 400
rect 199360 0 199416 400
rect 199696 0 199752 400
rect 200032 0 200088 400
rect 200368 0 200424 400
rect 200704 0 200760 400
rect 201040 0 201096 400
rect 201376 0 201432 400
rect 201712 0 201768 400
rect 202048 0 202104 400
rect 202384 0 202440 400
rect 202720 0 202776 400
rect 203056 0 203112 400
rect 203392 0 203448 400
rect 203728 0 203784 400
rect 204064 0 204120 400
rect 204400 0 204456 400
rect 204736 0 204792 400
rect 205072 0 205128 400
rect 205408 0 205464 400
rect 205744 0 205800 400
rect 206080 0 206136 400
rect 206416 0 206472 400
rect 206752 0 206808 400
rect 207088 0 207144 400
rect 207424 0 207480 400
rect 207760 0 207816 400
rect 208096 0 208152 400
rect 208432 0 208488 400
rect 208768 0 208824 400
rect 209104 0 209160 400
rect 209440 0 209496 400
rect 209776 0 209832 400
rect 210112 0 210168 400
rect 210448 0 210504 400
rect 210784 0 210840 400
rect 211120 0 211176 400
rect 211456 0 211512 400
rect 211792 0 211848 400
rect 212128 0 212184 400
rect 212464 0 212520 400
rect 212800 0 212856 400
rect 213136 0 213192 400
rect 213472 0 213528 400
rect 213808 0 213864 400
rect 214144 0 214200 400
rect 214480 0 214536 400
rect 214816 0 214872 400
rect 215152 0 215208 400
rect 215488 0 215544 400
rect 215824 0 215880 400
rect 216160 0 216216 400
rect 216496 0 216552 400
rect 216832 0 216888 400
rect 217168 0 217224 400
rect 217504 0 217560 400
rect 217840 0 217896 400
rect 218176 0 218232 400
rect 218512 0 218568 400
rect 218848 0 218904 400
rect 219184 0 219240 400
rect 219520 0 219576 400
rect 219856 0 219912 400
rect 220192 0 220248 400
rect 220528 0 220584 400
rect 220864 0 220920 400
rect 221200 0 221256 400
rect 221536 0 221592 400
rect 221872 0 221928 400
rect 222208 0 222264 400
rect 222544 0 222600 400
rect 222880 0 222936 400
rect 223216 0 223272 400
rect 223552 0 223608 400
rect 223888 0 223944 400
rect 224224 0 224280 400
rect 224560 0 224616 400
rect 224896 0 224952 400
rect 225232 0 225288 400
rect 225568 0 225624 400
rect 225904 0 225960 400
rect 226240 0 226296 400
rect 226576 0 226632 400
rect 226912 0 226968 400
rect 227248 0 227304 400
rect 227584 0 227640 400
rect 227920 0 227976 400
rect 228256 0 228312 400
rect 228592 0 228648 400
rect 228928 0 228984 400
rect 229264 0 229320 400
rect 229600 0 229656 400
rect 229936 0 229992 400
rect 230272 0 230328 400
rect 230608 0 230664 400
rect 230944 0 231000 400
rect 231280 0 231336 400
rect 231616 0 231672 400
rect 231952 0 232008 400
rect 232288 0 232344 400
rect 232624 0 232680 400
rect 232960 0 233016 400
rect 233296 0 233352 400
rect 233632 0 233688 400
rect 233968 0 234024 400
rect 234304 0 234360 400
rect 234640 0 234696 400
rect 234976 0 235032 400
rect 235312 0 235368 400
rect 235648 0 235704 400
rect 235984 0 236040 400
rect 236320 0 236376 400
rect 236656 0 236712 400
rect 236992 0 237048 400
rect 237328 0 237384 400
rect 237664 0 237720 400
rect 238000 0 238056 400
rect 238336 0 238392 400
rect 238672 0 238728 400
rect 239008 0 239064 400
rect 239344 0 239400 400
rect 239680 0 239736 400
rect 240016 0 240072 400
rect 240352 0 240408 400
rect 240688 0 240744 400
rect 241024 0 241080 400
rect 241360 0 241416 400
rect 241696 0 241752 400
rect 242032 0 242088 400
rect 242368 0 242424 400
rect 242704 0 242760 400
rect 243040 0 243096 400
rect 243376 0 243432 400
rect 243712 0 243768 400
rect 244048 0 244104 400
rect 244384 0 244440 400
rect 244720 0 244776 400
rect 245056 0 245112 400
rect 245392 0 245448 400
rect 245728 0 245784 400
rect 246064 0 246120 400
rect 246400 0 246456 400
rect 246736 0 246792 400
rect 247072 0 247128 400
rect 247408 0 247464 400
rect 247744 0 247800 400
rect 248080 0 248136 400
rect 248416 0 248472 400
rect 248752 0 248808 400
rect 249088 0 249144 400
rect 249424 0 249480 400
rect 249760 0 249816 400
rect 250096 0 250152 400
rect 250432 0 250488 400
rect 250768 0 250824 400
rect 251104 0 251160 400
rect 251440 0 251496 400
rect 251776 0 251832 400
rect 252112 0 252168 400
rect 252448 0 252504 400
rect 252784 0 252840 400
rect 253120 0 253176 400
rect 253456 0 253512 400
rect 253792 0 253848 400
rect 254128 0 254184 400
rect 254464 0 254520 400
rect 254800 0 254856 400
rect 255136 0 255192 400
rect 255472 0 255528 400
rect 255808 0 255864 400
rect 256144 0 256200 400
rect 256480 0 256536 400
rect 256816 0 256872 400
rect 257152 0 257208 400
rect 257488 0 257544 400
rect 257824 0 257880 400
rect 258160 0 258216 400
rect 258496 0 258552 400
rect 258832 0 258888 400
rect 259168 0 259224 400
rect 259504 0 259560 400
rect 259840 0 259896 400
rect 260176 0 260232 400
rect 260512 0 260568 400
rect 260848 0 260904 400
rect 261184 0 261240 400
rect 261520 0 261576 400
rect 261856 0 261912 400
rect 262192 0 262248 400
rect 262528 0 262584 400
rect 262864 0 262920 400
rect 263200 0 263256 400
rect 263536 0 263592 400
rect 263872 0 263928 400
rect 264208 0 264264 400
rect 264544 0 264600 400
rect 264880 0 264936 400
rect 265216 0 265272 400
rect 265552 0 265608 400
rect 265888 0 265944 400
rect 266224 0 266280 400
rect 266560 0 266616 400
rect 266896 0 266952 400
rect 267232 0 267288 400
rect 267568 0 267624 400
rect 267904 0 267960 400
rect 268240 0 268296 400
rect 268576 0 268632 400
rect 268912 0 268968 400
rect 269248 0 269304 400
rect 269584 0 269640 400
rect 269920 0 269976 400
rect 270256 0 270312 400
rect 270592 0 270648 400
rect 270928 0 270984 400
rect 271264 0 271320 400
rect 271600 0 271656 400
rect 271936 0 271992 400
rect 272272 0 272328 400
rect 272608 0 272664 400
rect 272944 0 273000 400
rect 273280 0 273336 400
rect 273616 0 273672 400
rect 273952 0 274008 400
rect 274288 0 274344 400
rect 274624 0 274680 400
rect 274960 0 275016 400
rect 275296 0 275352 400
rect 275632 0 275688 400
rect 275968 0 276024 400
rect 276304 0 276360 400
<< obsm2 >>
rect 798 79570 3666 79600
rect 3782 79570 5794 79600
rect 5910 79570 7922 79600
rect 8038 79570 10050 79600
rect 10166 79570 12178 79600
rect 12294 79570 14306 79600
rect 14422 79570 16434 79600
rect 16550 79570 18562 79600
rect 18678 79570 20690 79600
rect 20806 79570 22818 79600
rect 22934 79570 24946 79600
rect 25062 79570 27074 79600
rect 27190 79570 29202 79600
rect 29318 79570 31330 79600
rect 31446 79570 33458 79600
rect 33574 79570 35586 79600
rect 35702 79570 37714 79600
rect 37830 79570 39842 79600
rect 39958 79570 41970 79600
rect 42086 79570 44098 79600
rect 44214 79570 46226 79600
rect 46342 79570 48354 79600
rect 48470 79570 50482 79600
rect 50598 79570 52610 79600
rect 52726 79570 54738 79600
rect 54854 79570 56866 79600
rect 56982 79570 58994 79600
rect 59110 79570 61122 79600
rect 61238 79570 63250 79600
rect 63366 79570 65378 79600
rect 65494 79570 67506 79600
rect 67622 79570 69634 79600
rect 69750 79570 71762 79600
rect 71878 79570 73890 79600
rect 74006 79570 76018 79600
rect 76134 79570 78146 79600
rect 78262 79570 80274 79600
rect 80390 79570 82402 79600
rect 82518 79570 84530 79600
rect 84646 79570 86658 79600
rect 86774 79570 88786 79600
rect 88902 79570 90914 79600
rect 91030 79570 93042 79600
rect 93158 79570 95170 79600
rect 95286 79570 97298 79600
rect 97414 79570 99426 79600
rect 99542 79570 101554 79600
rect 101670 79570 103682 79600
rect 103798 79570 105810 79600
rect 105926 79570 107938 79600
rect 108054 79570 110066 79600
rect 110182 79570 112194 79600
rect 112310 79570 114322 79600
rect 114438 79570 116450 79600
rect 116566 79570 118578 79600
rect 118694 79570 120706 79600
rect 120822 79570 122834 79600
rect 122950 79570 124962 79600
rect 125078 79570 127090 79600
rect 127206 79570 129218 79600
rect 129334 79570 131346 79600
rect 131462 79570 133474 79600
rect 133590 79570 135602 79600
rect 135718 79570 137730 79600
rect 137846 79570 139858 79600
rect 139974 79570 141986 79600
rect 142102 79570 144114 79600
rect 144230 79570 146242 79600
rect 146358 79570 148370 79600
rect 148486 79570 150498 79600
rect 150614 79570 152626 79600
rect 152742 79570 154754 79600
rect 154870 79570 156882 79600
rect 156998 79570 159010 79600
rect 159126 79570 161138 79600
rect 161254 79570 163266 79600
rect 163382 79570 165394 79600
rect 165510 79570 167522 79600
rect 167638 79570 169650 79600
rect 169766 79570 171778 79600
rect 171894 79570 173906 79600
rect 174022 79570 176034 79600
rect 176150 79570 178162 79600
rect 178278 79570 180290 79600
rect 180406 79570 182418 79600
rect 182534 79570 184546 79600
rect 184662 79570 186674 79600
rect 186790 79570 188802 79600
rect 188918 79570 190930 79600
rect 191046 79570 193058 79600
rect 193174 79570 195186 79600
rect 195302 79570 197314 79600
rect 197430 79570 199442 79600
rect 199558 79570 201570 79600
rect 201686 79570 203698 79600
rect 203814 79570 205826 79600
rect 205942 79570 207954 79600
rect 208070 79570 210082 79600
rect 210198 79570 212210 79600
rect 212326 79570 214338 79600
rect 214454 79570 216466 79600
rect 216582 79570 218594 79600
rect 218710 79570 220722 79600
rect 220838 79570 222850 79600
rect 222966 79570 224978 79600
rect 225094 79570 227106 79600
rect 227222 79570 229234 79600
rect 229350 79570 231362 79600
rect 231478 79570 233490 79600
rect 233606 79570 235618 79600
rect 235734 79570 237746 79600
rect 237862 79570 239874 79600
rect 239990 79570 242002 79600
rect 242118 79570 244130 79600
rect 244246 79570 246258 79600
rect 246374 79570 248386 79600
rect 248502 79570 250514 79600
rect 250630 79570 252642 79600
rect 252758 79570 254770 79600
rect 254886 79570 256898 79600
rect 257014 79570 259026 79600
rect 259142 79570 261154 79600
rect 261270 79570 263282 79600
rect 263398 79570 265410 79600
rect 265526 79570 267538 79600
rect 267654 79570 269666 79600
rect 269782 79570 271794 79600
rect 271910 79570 273922 79600
rect 274038 79570 276050 79600
rect 276166 79570 279146 79600
rect 798 430 279146 79570
rect 798 400 3442 430
rect 3558 400 3778 430
rect 3894 400 4114 430
rect 4230 400 4450 430
rect 4566 400 4786 430
rect 4902 400 5122 430
rect 5238 400 5458 430
rect 5574 400 5794 430
rect 5910 400 6130 430
rect 6246 400 6466 430
rect 6582 400 6802 430
rect 6918 400 7138 430
rect 7254 400 7474 430
rect 7590 400 7810 430
rect 7926 400 8146 430
rect 8262 400 8482 430
rect 8598 400 8818 430
rect 8934 400 9154 430
rect 9270 400 9490 430
rect 9606 400 9826 430
rect 9942 400 10162 430
rect 10278 400 10498 430
rect 10614 400 10834 430
rect 10950 400 11170 430
rect 11286 400 11506 430
rect 11622 400 11842 430
rect 11958 400 12178 430
rect 12294 400 12514 430
rect 12630 400 12850 430
rect 12966 400 13186 430
rect 13302 400 13522 430
rect 13638 400 13858 430
rect 13974 400 14194 430
rect 14310 400 14530 430
rect 14646 400 14866 430
rect 14982 400 15202 430
rect 15318 400 15538 430
rect 15654 400 15874 430
rect 15990 400 16210 430
rect 16326 400 16546 430
rect 16662 400 16882 430
rect 16998 400 17218 430
rect 17334 400 17554 430
rect 17670 400 17890 430
rect 18006 400 18226 430
rect 18342 400 18562 430
rect 18678 400 18898 430
rect 19014 400 19234 430
rect 19350 400 19570 430
rect 19686 400 19906 430
rect 20022 400 20242 430
rect 20358 400 20578 430
rect 20694 400 20914 430
rect 21030 400 21250 430
rect 21366 400 21586 430
rect 21702 400 21922 430
rect 22038 400 22258 430
rect 22374 400 22594 430
rect 22710 400 22930 430
rect 23046 400 23266 430
rect 23382 400 23602 430
rect 23718 400 23938 430
rect 24054 400 24274 430
rect 24390 400 24610 430
rect 24726 400 24946 430
rect 25062 400 25282 430
rect 25398 400 25618 430
rect 25734 400 25954 430
rect 26070 400 26290 430
rect 26406 400 26626 430
rect 26742 400 26962 430
rect 27078 400 27298 430
rect 27414 400 27634 430
rect 27750 400 27970 430
rect 28086 400 28306 430
rect 28422 400 28642 430
rect 28758 400 28978 430
rect 29094 400 29314 430
rect 29430 400 29650 430
rect 29766 400 29986 430
rect 30102 400 30322 430
rect 30438 400 30658 430
rect 30774 400 30994 430
rect 31110 400 31330 430
rect 31446 400 31666 430
rect 31782 400 32002 430
rect 32118 400 32338 430
rect 32454 400 32674 430
rect 32790 400 33010 430
rect 33126 400 33346 430
rect 33462 400 33682 430
rect 33798 400 34018 430
rect 34134 400 34354 430
rect 34470 400 34690 430
rect 34806 400 35026 430
rect 35142 400 35362 430
rect 35478 400 35698 430
rect 35814 400 36034 430
rect 36150 400 36370 430
rect 36486 400 36706 430
rect 36822 400 37042 430
rect 37158 400 37378 430
rect 37494 400 37714 430
rect 37830 400 38050 430
rect 38166 400 38386 430
rect 38502 400 38722 430
rect 38838 400 39058 430
rect 39174 400 39394 430
rect 39510 400 39730 430
rect 39846 400 40066 430
rect 40182 400 40402 430
rect 40518 400 40738 430
rect 40854 400 41074 430
rect 41190 400 41410 430
rect 41526 400 41746 430
rect 41862 400 42082 430
rect 42198 400 42418 430
rect 42534 400 42754 430
rect 42870 400 43090 430
rect 43206 400 43426 430
rect 43542 400 43762 430
rect 43878 400 44098 430
rect 44214 400 44434 430
rect 44550 400 44770 430
rect 44886 400 45106 430
rect 45222 400 45442 430
rect 45558 400 45778 430
rect 45894 400 46114 430
rect 46230 400 46450 430
rect 46566 400 46786 430
rect 46902 400 47122 430
rect 47238 400 47458 430
rect 47574 400 47794 430
rect 47910 400 48130 430
rect 48246 400 48466 430
rect 48582 400 48802 430
rect 48918 400 49138 430
rect 49254 400 49474 430
rect 49590 400 49810 430
rect 49926 400 50146 430
rect 50262 400 50482 430
rect 50598 400 50818 430
rect 50934 400 51154 430
rect 51270 400 51490 430
rect 51606 400 51826 430
rect 51942 400 52162 430
rect 52278 400 52498 430
rect 52614 400 52834 430
rect 52950 400 53170 430
rect 53286 400 53506 430
rect 53622 400 53842 430
rect 53958 400 54178 430
rect 54294 400 54514 430
rect 54630 400 54850 430
rect 54966 400 55186 430
rect 55302 400 55522 430
rect 55638 400 55858 430
rect 55974 400 56194 430
rect 56310 400 56530 430
rect 56646 400 56866 430
rect 56982 400 57202 430
rect 57318 400 57538 430
rect 57654 400 57874 430
rect 57990 400 58210 430
rect 58326 400 58546 430
rect 58662 400 58882 430
rect 58998 400 59218 430
rect 59334 400 59554 430
rect 59670 400 59890 430
rect 60006 400 60226 430
rect 60342 400 60562 430
rect 60678 400 60898 430
rect 61014 400 61234 430
rect 61350 400 61570 430
rect 61686 400 61906 430
rect 62022 400 62242 430
rect 62358 400 62578 430
rect 62694 400 62914 430
rect 63030 400 63250 430
rect 63366 400 63586 430
rect 63702 400 63922 430
rect 64038 400 64258 430
rect 64374 400 64594 430
rect 64710 400 64930 430
rect 65046 400 65266 430
rect 65382 400 65602 430
rect 65718 400 65938 430
rect 66054 400 66274 430
rect 66390 400 66610 430
rect 66726 400 66946 430
rect 67062 400 67282 430
rect 67398 400 67618 430
rect 67734 400 67954 430
rect 68070 400 68290 430
rect 68406 400 68626 430
rect 68742 400 68962 430
rect 69078 400 69298 430
rect 69414 400 69634 430
rect 69750 400 69970 430
rect 70086 400 70306 430
rect 70422 400 70642 430
rect 70758 400 70978 430
rect 71094 400 71314 430
rect 71430 400 71650 430
rect 71766 400 71986 430
rect 72102 400 72322 430
rect 72438 400 72658 430
rect 72774 400 72994 430
rect 73110 400 73330 430
rect 73446 400 73666 430
rect 73782 400 74002 430
rect 74118 400 74338 430
rect 74454 400 74674 430
rect 74790 400 75010 430
rect 75126 400 75346 430
rect 75462 400 75682 430
rect 75798 400 76018 430
rect 76134 400 76354 430
rect 76470 400 76690 430
rect 76806 400 77026 430
rect 77142 400 77362 430
rect 77478 400 77698 430
rect 77814 400 78034 430
rect 78150 400 78370 430
rect 78486 400 78706 430
rect 78822 400 79042 430
rect 79158 400 79378 430
rect 79494 400 79714 430
rect 79830 400 80050 430
rect 80166 400 80386 430
rect 80502 400 80722 430
rect 80838 400 81058 430
rect 81174 400 81394 430
rect 81510 400 81730 430
rect 81846 400 82066 430
rect 82182 400 82402 430
rect 82518 400 82738 430
rect 82854 400 83074 430
rect 83190 400 83410 430
rect 83526 400 83746 430
rect 83862 400 84082 430
rect 84198 400 84418 430
rect 84534 400 84754 430
rect 84870 400 85090 430
rect 85206 400 85426 430
rect 85542 400 85762 430
rect 85878 400 86098 430
rect 86214 400 86434 430
rect 86550 400 86770 430
rect 86886 400 87106 430
rect 87222 400 87442 430
rect 87558 400 87778 430
rect 87894 400 88114 430
rect 88230 400 88450 430
rect 88566 400 88786 430
rect 88902 400 89122 430
rect 89238 400 89458 430
rect 89574 400 89794 430
rect 89910 400 90130 430
rect 90246 400 90466 430
rect 90582 400 90802 430
rect 90918 400 91138 430
rect 91254 400 91474 430
rect 91590 400 91810 430
rect 91926 400 92146 430
rect 92262 400 92482 430
rect 92598 400 92818 430
rect 92934 400 93154 430
rect 93270 400 93490 430
rect 93606 400 93826 430
rect 93942 400 94162 430
rect 94278 400 94498 430
rect 94614 400 94834 430
rect 94950 400 95170 430
rect 95286 400 95506 430
rect 95622 400 95842 430
rect 95958 400 96178 430
rect 96294 400 96514 430
rect 96630 400 96850 430
rect 96966 400 97186 430
rect 97302 400 97522 430
rect 97638 400 97858 430
rect 97974 400 98194 430
rect 98310 400 98530 430
rect 98646 400 98866 430
rect 98982 400 99202 430
rect 99318 400 99538 430
rect 99654 400 99874 430
rect 99990 400 100210 430
rect 100326 400 100546 430
rect 100662 400 100882 430
rect 100998 400 101218 430
rect 101334 400 101554 430
rect 101670 400 101890 430
rect 102006 400 102226 430
rect 102342 400 102562 430
rect 102678 400 102898 430
rect 103014 400 103234 430
rect 103350 400 103570 430
rect 103686 400 103906 430
rect 104022 400 104242 430
rect 104358 400 104578 430
rect 104694 400 104914 430
rect 105030 400 105250 430
rect 105366 400 105586 430
rect 105702 400 105922 430
rect 106038 400 106258 430
rect 106374 400 106594 430
rect 106710 400 106930 430
rect 107046 400 107266 430
rect 107382 400 107602 430
rect 107718 400 107938 430
rect 108054 400 108274 430
rect 108390 400 108610 430
rect 108726 400 108946 430
rect 109062 400 109282 430
rect 109398 400 109618 430
rect 109734 400 109954 430
rect 110070 400 110290 430
rect 110406 400 110626 430
rect 110742 400 110962 430
rect 111078 400 111298 430
rect 111414 400 111634 430
rect 111750 400 111970 430
rect 112086 400 112306 430
rect 112422 400 112642 430
rect 112758 400 112978 430
rect 113094 400 113314 430
rect 113430 400 113650 430
rect 113766 400 113986 430
rect 114102 400 114322 430
rect 114438 400 114658 430
rect 114774 400 114994 430
rect 115110 400 115330 430
rect 115446 400 115666 430
rect 115782 400 116002 430
rect 116118 400 116338 430
rect 116454 400 116674 430
rect 116790 400 117010 430
rect 117126 400 117346 430
rect 117462 400 117682 430
rect 117798 400 118018 430
rect 118134 400 118354 430
rect 118470 400 118690 430
rect 118806 400 119026 430
rect 119142 400 119362 430
rect 119478 400 119698 430
rect 119814 400 120034 430
rect 120150 400 120370 430
rect 120486 400 120706 430
rect 120822 400 121042 430
rect 121158 400 121378 430
rect 121494 400 121714 430
rect 121830 400 122050 430
rect 122166 400 122386 430
rect 122502 400 122722 430
rect 122838 400 123058 430
rect 123174 400 123394 430
rect 123510 400 123730 430
rect 123846 400 124066 430
rect 124182 400 124402 430
rect 124518 400 124738 430
rect 124854 400 125074 430
rect 125190 400 125410 430
rect 125526 400 125746 430
rect 125862 400 126082 430
rect 126198 400 126418 430
rect 126534 400 126754 430
rect 126870 400 127090 430
rect 127206 400 127426 430
rect 127542 400 127762 430
rect 127878 400 128098 430
rect 128214 400 128434 430
rect 128550 400 128770 430
rect 128886 400 129106 430
rect 129222 400 129442 430
rect 129558 400 129778 430
rect 129894 400 130114 430
rect 130230 400 130450 430
rect 130566 400 130786 430
rect 130902 400 131122 430
rect 131238 400 131458 430
rect 131574 400 131794 430
rect 131910 400 132130 430
rect 132246 400 132466 430
rect 132582 400 132802 430
rect 132918 400 133138 430
rect 133254 400 133474 430
rect 133590 400 133810 430
rect 133926 400 134146 430
rect 134262 400 134482 430
rect 134598 400 134818 430
rect 134934 400 135154 430
rect 135270 400 135490 430
rect 135606 400 135826 430
rect 135942 400 136162 430
rect 136278 400 136498 430
rect 136614 400 136834 430
rect 136950 400 137170 430
rect 137286 400 137506 430
rect 137622 400 137842 430
rect 137958 400 138178 430
rect 138294 400 138514 430
rect 138630 400 138850 430
rect 138966 400 139186 430
rect 139302 400 139522 430
rect 139638 400 139858 430
rect 139974 400 140194 430
rect 140310 400 140530 430
rect 140646 400 140866 430
rect 140982 400 141202 430
rect 141318 400 141538 430
rect 141654 400 141874 430
rect 141990 400 142210 430
rect 142326 400 142546 430
rect 142662 400 142882 430
rect 142998 400 143218 430
rect 143334 400 143554 430
rect 143670 400 143890 430
rect 144006 400 144226 430
rect 144342 400 144562 430
rect 144678 400 144898 430
rect 145014 400 145234 430
rect 145350 400 145570 430
rect 145686 400 145906 430
rect 146022 400 146242 430
rect 146358 400 146578 430
rect 146694 400 146914 430
rect 147030 400 147250 430
rect 147366 400 147586 430
rect 147702 400 147922 430
rect 148038 400 148258 430
rect 148374 400 148594 430
rect 148710 400 148930 430
rect 149046 400 149266 430
rect 149382 400 149602 430
rect 149718 400 149938 430
rect 150054 400 150274 430
rect 150390 400 150610 430
rect 150726 400 150946 430
rect 151062 400 151282 430
rect 151398 400 151618 430
rect 151734 400 151954 430
rect 152070 400 152290 430
rect 152406 400 152626 430
rect 152742 400 152962 430
rect 153078 400 153298 430
rect 153414 400 153634 430
rect 153750 400 153970 430
rect 154086 400 154306 430
rect 154422 400 154642 430
rect 154758 400 154978 430
rect 155094 400 155314 430
rect 155430 400 155650 430
rect 155766 400 155986 430
rect 156102 400 156322 430
rect 156438 400 156658 430
rect 156774 400 156994 430
rect 157110 400 157330 430
rect 157446 400 157666 430
rect 157782 400 158002 430
rect 158118 400 158338 430
rect 158454 400 158674 430
rect 158790 400 159010 430
rect 159126 400 159346 430
rect 159462 400 159682 430
rect 159798 400 160018 430
rect 160134 400 160354 430
rect 160470 400 160690 430
rect 160806 400 161026 430
rect 161142 400 161362 430
rect 161478 400 161698 430
rect 161814 400 162034 430
rect 162150 400 162370 430
rect 162486 400 162706 430
rect 162822 400 163042 430
rect 163158 400 163378 430
rect 163494 400 163714 430
rect 163830 400 164050 430
rect 164166 400 164386 430
rect 164502 400 164722 430
rect 164838 400 165058 430
rect 165174 400 165394 430
rect 165510 400 165730 430
rect 165846 400 166066 430
rect 166182 400 166402 430
rect 166518 400 166738 430
rect 166854 400 167074 430
rect 167190 400 167410 430
rect 167526 400 167746 430
rect 167862 400 168082 430
rect 168198 400 168418 430
rect 168534 400 168754 430
rect 168870 400 169090 430
rect 169206 400 169426 430
rect 169542 400 169762 430
rect 169878 400 170098 430
rect 170214 400 170434 430
rect 170550 400 170770 430
rect 170886 400 171106 430
rect 171222 400 171442 430
rect 171558 400 171778 430
rect 171894 400 172114 430
rect 172230 400 172450 430
rect 172566 400 172786 430
rect 172902 400 173122 430
rect 173238 400 173458 430
rect 173574 400 173794 430
rect 173910 400 174130 430
rect 174246 400 174466 430
rect 174582 400 174802 430
rect 174918 400 175138 430
rect 175254 400 175474 430
rect 175590 400 175810 430
rect 175926 400 176146 430
rect 176262 400 176482 430
rect 176598 400 176818 430
rect 176934 400 177154 430
rect 177270 400 177490 430
rect 177606 400 177826 430
rect 177942 400 178162 430
rect 178278 400 178498 430
rect 178614 400 178834 430
rect 178950 400 179170 430
rect 179286 400 179506 430
rect 179622 400 179842 430
rect 179958 400 180178 430
rect 180294 400 180514 430
rect 180630 400 180850 430
rect 180966 400 181186 430
rect 181302 400 181522 430
rect 181638 400 181858 430
rect 181974 400 182194 430
rect 182310 400 182530 430
rect 182646 400 182866 430
rect 182982 400 183202 430
rect 183318 400 183538 430
rect 183654 400 183874 430
rect 183990 400 184210 430
rect 184326 400 184546 430
rect 184662 400 184882 430
rect 184998 400 185218 430
rect 185334 400 185554 430
rect 185670 400 185890 430
rect 186006 400 186226 430
rect 186342 400 186562 430
rect 186678 400 186898 430
rect 187014 400 187234 430
rect 187350 400 187570 430
rect 187686 400 187906 430
rect 188022 400 188242 430
rect 188358 400 188578 430
rect 188694 400 188914 430
rect 189030 400 189250 430
rect 189366 400 189586 430
rect 189702 400 189922 430
rect 190038 400 190258 430
rect 190374 400 190594 430
rect 190710 400 190930 430
rect 191046 400 191266 430
rect 191382 400 191602 430
rect 191718 400 191938 430
rect 192054 400 192274 430
rect 192390 400 192610 430
rect 192726 400 192946 430
rect 193062 400 193282 430
rect 193398 400 193618 430
rect 193734 400 193954 430
rect 194070 400 194290 430
rect 194406 400 194626 430
rect 194742 400 194962 430
rect 195078 400 195298 430
rect 195414 400 195634 430
rect 195750 400 195970 430
rect 196086 400 196306 430
rect 196422 400 196642 430
rect 196758 400 196978 430
rect 197094 400 197314 430
rect 197430 400 197650 430
rect 197766 400 197986 430
rect 198102 400 198322 430
rect 198438 400 198658 430
rect 198774 400 198994 430
rect 199110 400 199330 430
rect 199446 400 199666 430
rect 199782 400 200002 430
rect 200118 400 200338 430
rect 200454 400 200674 430
rect 200790 400 201010 430
rect 201126 400 201346 430
rect 201462 400 201682 430
rect 201798 400 202018 430
rect 202134 400 202354 430
rect 202470 400 202690 430
rect 202806 400 203026 430
rect 203142 400 203362 430
rect 203478 400 203698 430
rect 203814 400 204034 430
rect 204150 400 204370 430
rect 204486 400 204706 430
rect 204822 400 205042 430
rect 205158 400 205378 430
rect 205494 400 205714 430
rect 205830 400 206050 430
rect 206166 400 206386 430
rect 206502 400 206722 430
rect 206838 400 207058 430
rect 207174 400 207394 430
rect 207510 400 207730 430
rect 207846 400 208066 430
rect 208182 400 208402 430
rect 208518 400 208738 430
rect 208854 400 209074 430
rect 209190 400 209410 430
rect 209526 400 209746 430
rect 209862 400 210082 430
rect 210198 400 210418 430
rect 210534 400 210754 430
rect 210870 400 211090 430
rect 211206 400 211426 430
rect 211542 400 211762 430
rect 211878 400 212098 430
rect 212214 400 212434 430
rect 212550 400 212770 430
rect 212886 400 213106 430
rect 213222 400 213442 430
rect 213558 400 213778 430
rect 213894 400 214114 430
rect 214230 400 214450 430
rect 214566 400 214786 430
rect 214902 400 215122 430
rect 215238 400 215458 430
rect 215574 400 215794 430
rect 215910 400 216130 430
rect 216246 400 216466 430
rect 216582 400 216802 430
rect 216918 400 217138 430
rect 217254 400 217474 430
rect 217590 400 217810 430
rect 217926 400 218146 430
rect 218262 400 218482 430
rect 218598 400 218818 430
rect 218934 400 219154 430
rect 219270 400 219490 430
rect 219606 400 219826 430
rect 219942 400 220162 430
rect 220278 400 220498 430
rect 220614 400 220834 430
rect 220950 400 221170 430
rect 221286 400 221506 430
rect 221622 400 221842 430
rect 221958 400 222178 430
rect 222294 400 222514 430
rect 222630 400 222850 430
rect 222966 400 223186 430
rect 223302 400 223522 430
rect 223638 400 223858 430
rect 223974 400 224194 430
rect 224310 400 224530 430
rect 224646 400 224866 430
rect 224982 400 225202 430
rect 225318 400 225538 430
rect 225654 400 225874 430
rect 225990 400 226210 430
rect 226326 400 226546 430
rect 226662 400 226882 430
rect 226998 400 227218 430
rect 227334 400 227554 430
rect 227670 400 227890 430
rect 228006 400 228226 430
rect 228342 400 228562 430
rect 228678 400 228898 430
rect 229014 400 229234 430
rect 229350 400 229570 430
rect 229686 400 229906 430
rect 230022 400 230242 430
rect 230358 400 230578 430
rect 230694 400 230914 430
rect 231030 400 231250 430
rect 231366 400 231586 430
rect 231702 400 231922 430
rect 232038 400 232258 430
rect 232374 400 232594 430
rect 232710 400 232930 430
rect 233046 400 233266 430
rect 233382 400 233602 430
rect 233718 400 233938 430
rect 234054 400 234274 430
rect 234390 400 234610 430
rect 234726 400 234946 430
rect 235062 400 235282 430
rect 235398 400 235618 430
rect 235734 400 235954 430
rect 236070 400 236290 430
rect 236406 400 236626 430
rect 236742 400 236962 430
rect 237078 400 237298 430
rect 237414 400 237634 430
rect 237750 400 237970 430
rect 238086 400 238306 430
rect 238422 400 238642 430
rect 238758 400 238978 430
rect 239094 400 239314 430
rect 239430 400 239650 430
rect 239766 400 239986 430
rect 240102 400 240322 430
rect 240438 400 240658 430
rect 240774 400 240994 430
rect 241110 400 241330 430
rect 241446 400 241666 430
rect 241782 400 242002 430
rect 242118 400 242338 430
rect 242454 400 242674 430
rect 242790 400 243010 430
rect 243126 400 243346 430
rect 243462 400 243682 430
rect 243798 400 244018 430
rect 244134 400 244354 430
rect 244470 400 244690 430
rect 244806 400 245026 430
rect 245142 400 245362 430
rect 245478 400 245698 430
rect 245814 400 246034 430
rect 246150 400 246370 430
rect 246486 400 246706 430
rect 246822 400 247042 430
rect 247158 400 247378 430
rect 247494 400 247714 430
rect 247830 400 248050 430
rect 248166 400 248386 430
rect 248502 400 248722 430
rect 248838 400 249058 430
rect 249174 400 249394 430
rect 249510 400 249730 430
rect 249846 400 250066 430
rect 250182 400 250402 430
rect 250518 400 250738 430
rect 250854 400 251074 430
rect 251190 400 251410 430
rect 251526 400 251746 430
rect 251862 400 252082 430
rect 252198 400 252418 430
rect 252534 400 252754 430
rect 252870 400 253090 430
rect 253206 400 253426 430
rect 253542 400 253762 430
rect 253878 400 254098 430
rect 254214 400 254434 430
rect 254550 400 254770 430
rect 254886 400 255106 430
rect 255222 400 255442 430
rect 255558 400 255778 430
rect 255894 400 256114 430
rect 256230 400 256450 430
rect 256566 400 256786 430
rect 256902 400 257122 430
rect 257238 400 257458 430
rect 257574 400 257794 430
rect 257910 400 258130 430
rect 258246 400 258466 430
rect 258582 400 258802 430
rect 258918 400 259138 430
rect 259254 400 259474 430
rect 259590 400 259810 430
rect 259926 400 260146 430
rect 260262 400 260482 430
rect 260598 400 260818 430
rect 260934 400 261154 430
rect 261270 400 261490 430
rect 261606 400 261826 430
rect 261942 400 262162 430
rect 262278 400 262498 430
rect 262614 400 262834 430
rect 262950 400 263170 430
rect 263286 400 263506 430
rect 263622 400 263842 430
rect 263958 400 264178 430
rect 264294 400 264514 430
rect 264630 400 264850 430
rect 264966 400 265186 430
rect 265302 400 265522 430
rect 265638 400 265858 430
rect 265974 400 266194 430
rect 266310 400 266530 430
rect 266646 400 266866 430
rect 266982 400 267202 430
rect 267318 400 267538 430
rect 267654 400 267874 430
rect 267990 400 268210 430
rect 268326 400 268546 430
rect 268662 400 268882 430
rect 268998 400 269218 430
rect 269334 400 269554 430
rect 269670 400 269890 430
rect 270006 400 270226 430
rect 270342 400 270562 430
rect 270678 400 270898 430
rect 271014 400 271234 430
rect 271350 400 271570 430
rect 271686 400 271906 430
rect 272022 400 272242 430
rect 272358 400 272578 430
rect 272694 400 272914 430
rect 273030 400 273250 430
rect 273366 400 273586 430
rect 273702 400 273922 430
rect 274038 400 274258 430
rect 274374 400 274594 430
rect 274710 400 274930 430
rect 275046 400 275266 430
rect 275382 400 275602 430
rect 275718 400 275938 430
rect 276054 400 276274 430
rect 276390 400 279146 430
<< metal3 >>
rect 0 69888 400 69944
rect 0 69776 400 69832
rect 0 69664 400 69720
rect 0 69552 400 69608
rect 0 69440 400 69496
rect 0 69328 400 69384
rect 0 69216 400 69272
rect 0 69104 400 69160
rect 0 68992 400 69048
rect 0 68880 400 68936
rect 0 68768 400 68824
rect 0 68656 400 68712
rect 0 68544 400 68600
rect 0 68432 400 68488
rect 0 68320 400 68376
rect 0 68208 400 68264
rect 0 68096 400 68152
rect 0 67984 400 68040
rect 0 67872 400 67928
rect 0 67760 400 67816
rect 0 67648 400 67704
rect 0 67536 400 67592
rect 0 67424 400 67480
rect 0 67312 400 67368
rect 0 67200 400 67256
rect 0 67088 400 67144
rect 0 66976 400 67032
rect 0 66864 400 66920
rect 0 66752 400 66808
rect 0 66640 400 66696
rect 0 66528 400 66584
rect 0 66416 400 66472
rect 0 66304 400 66360
rect 0 66192 400 66248
rect 0 66080 400 66136
rect 0 65968 400 66024
rect 0 65856 400 65912
rect 0 65744 400 65800
rect 0 65632 400 65688
rect 0 65520 400 65576
rect 0 65408 400 65464
rect 0 65296 400 65352
rect 0 65184 400 65240
rect 0 65072 400 65128
rect 0 64960 400 65016
rect 0 64848 400 64904
rect 0 64736 400 64792
rect 0 64624 400 64680
rect 0 64512 400 64568
rect 0 64400 400 64456
rect 0 64288 400 64344
rect 0 64176 400 64232
rect 0 64064 400 64120
rect 0 63952 400 64008
rect 0 63840 400 63896
rect 0 63728 400 63784
rect 0 63616 400 63672
rect 0 63504 400 63560
rect 0 63392 400 63448
rect 0 63280 400 63336
rect 0 63168 400 63224
rect 0 63056 400 63112
rect 0 62944 400 63000
rect 0 62832 400 62888
rect 0 62720 400 62776
rect 0 62608 400 62664
rect 0 62496 400 62552
rect 0 62384 400 62440
rect 0 62272 400 62328
rect 0 62160 400 62216
rect 0 62048 400 62104
rect 0 61936 400 61992
rect 0 61824 400 61880
rect 0 61712 400 61768
rect 0 61600 400 61656
rect 0 61488 400 61544
rect 0 61376 400 61432
rect 0 61264 400 61320
rect 0 61152 400 61208
rect 0 61040 400 61096
rect 0 60928 400 60984
rect 0 60816 400 60872
rect 0 60704 400 60760
rect 0 60592 400 60648
rect 0 60480 400 60536
rect 0 60368 400 60424
rect 0 60256 400 60312
rect 0 60144 400 60200
rect 0 60032 400 60088
rect 0 59920 400 59976
rect 0 59808 400 59864
rect 0 59696 400 59752
rect 0 59584 400 59640
rect 0 59472 400 59528
rect 0 59360 400 59416
rect 0 59248 400 59304
rect 0 59136 400 59192
rect 0 59024 400 59080
rect 0 58912 400 58968
rect 0 58800 400 58856
rect 0 58688 400 58744
rect 0 58576 400 58632
rect 0 58464 400 58520
rect 0 58352 400 58408
rect 0 58240 400 58296
rect 0 58128 400 58184
rect 0 58016 400 58072
rect 0 57904 400 57960
rect 0 57792 400 57848
rect 0 57680 400 57736
rect 0 57568 400 57624
rect 0 57456 400 57512
rect 0 57344 400 57400
rect 0 57232 400 57288
rect 0 57120 400 57176
rect 0 57008 400 57064
rect 0 56896 400 56952
rect 0 56784 400 56840
rect 0 56672 400 56728
rect 0 56560 400 56616
rect 0 56448 400 56504
rect 0 56336 400 56392
rect 0 56224 400 56280
rect 0 56112 400 56168
rect 0 56000 400 56056
rect 0 55888 400 55944
rect 0 55776 400 55832
rect 0 55664 400 55720
rect 0 55552 400 55608
rect 0 55440 400 55496
rect 0 55328 400 55384
rect 0 55216 400 55272
rect 0 55104 400 55160
rect 0 54992 400 55048
rect 0 54880 400 54936
rect 0 54768 400 54824
rect 0 54656 400 54712
rect 0 54544 400 54600
rect 0 54432 400 54488
rect 0 54320 400 54376
rect 0 54208 400 54264
rect 0 54096 400 54152
rect 0 53984 400 54040
rect 0 53872 400 53928
rect 0 53760 400 53816
rect 0 53648 400 53704
rect 0 53536 400 53592
rect 0 53424 400 53480
rect 0 53312 400 53368
rect 0 53200 400 53256
rect 0 53088 400 53144
rect 0 52976 400 53032
rect 0 52864 400 52920
rect 0 52752 400 52808
rect 0 52640 400 52696
rect 0 52528 400 52584
rect 0 52416 400 52472
rect 0 52304 400 52360
rect 0 52192 400 52248
rect 0 52080 400 52136
rect 0 51968 400 52024
rect 0 51856 400 51912
rect 0 51744 400 51800
rect 0 51632 400 51688
rect 0 51520 400 51576
rect 0 51408 400 51464
rect 0 51296 400 51352
rect 0 51184 400 51240
rect 0 51072 400 51128
rect 0 50960 400 51016
rect 0 50848 400 50904
rect 0 50736 400 50792
rect 0 50624 400 50680
rect 0 50512 400 50568
rect 0 50400 400 50456
rect 0 50288 400 50344
rect 0 50176 400 50232
rect 0 50064 400 50120
rect 0 49952 400 50008
rect 0 49840 400 49896
rect 0 49728 400 49784
rect 0 49616 400 49672
rect 0 49504 400 49560
rect 0 49392 400 49448
rect 0 49280 400 49336
rect 0 49168 400 49224
rect 0 49056 400 49112
rect 0 48944 400 49000
rect 0 48832 400 48888
rect 0 48720 400 48776
rect 0 48608 400 48664
rect 0 48496 400 48552
rect 0 48384 400 48440
rect 0 48272 400 48328
rect 0 48160 400 48216
rect 0 48048 400 48104
rect 0 47936 400 47992
rect 0 47824 400 47880
rect 0 47712 400 47768
rect 0 47600 400 47656
rect 0 47488 400 47544
rect 0 47376 400 47432
rect 0 47264 400 47320
rect 0 47152 400 47208
rect 0 47040 400 47096
rect 0 46928 400 46984
rect 0 46816 400 46872
rect 0 46704 400 46760
rect 0 46592 400 46648
rect 0 46480 400 46536
rect 0 46368 400 46424
rect 0 46256 400 46312
rect 0 46144 400 46200
rect 0 46032 400 46088
rect 0 45920 400 45976
rect 0 45808 400 45864
rect 0 45696 400 45752
rect 0 45584 400 45640
rect 0 45472 400 45528
rect 0 45360 400 45416
rect 0 45248 400 45304
rect 0 45136 400 45192
rect 0 45024 400 45080
rect 0 44912 400 44968
rect 0 44800 400 44856
rect 0 44688 400 44744
rect 0 44576 400 44632
rect 0 44464 400 44520
rect 0 44352 400 44408
rect 0 44240 400 44296
rect 0 44128 400 44184
rect 0 44016 400 44072
rect 0 43904 400 43960
rect 0 43792 400 43848
rect 0 43680 400 43736
rect 0 43568 400 43624
rect 0 43456 400 43512
rect 0 43344 400 43400
rect 0 43232 400 43288
rect 0 43120 400 43176
rect 0 43008 400 43064
rect 0 42896 400 42952
rect 0 42784 400 42840
rect 0 42672 400 42728
rect 0 42560 400 42616
rect 0 42448 400 42504
rect 0 42336 400 42392
rect 0 42224 400 42280
rect 0 42112 400 42168
rect 0 42000 400 42056
rect 0 41888 400 41944
rect 0 41776 400 41832
rect 0 41664 400 41720
rect 0 41552 400 41608
rect 0 41440 400 41496
rect 0 41328 400 41384
rect 0 41216 400 41272
rect 0 41104 400 41160
rect 0 40992 400 41048
rect 0 40880 400 40936
rect 0 40768 400 40824
rect 0 40656 400 40712
rect 0 40544 400 40600
rect 0 40432 400 40488
rect 0 40320 400 40376
rect 0 40208 400 40264
rect 0 40096 400 40152
rect 0 39984 400 40040
rect 0 39872 400 39928
rect 0 39760 400 39816
rect 0 39648 400 39704
rect 0 39536 400 39592
rect 0 39424 400 39480
rect 0 39312 400 39368
rect 0 39200 400 39256
rect 0 39088 400 39144
rect 0 38976 400 39032
rect 0 38864 400 38920
rect 0 38752 400 38808
rect 0 38640 400 38696
rect 0 38528 400 38584
rect 0 38416 400 38472
rect 0 38304 400 38360
rect 0 38192 400 38248
rect 0 38080 400 38136
rect 0 37968 400 38024
rect 0 37856 400 37912
rect 0 37744 400 37800
rect 0 37632 400 37688
rect 0 37520 400 37576
rect 0 37408 400 37464
rect 0 37296 400 37352
rect 0 37184 400 37240
rect 0 37072 400 37128
rect 0 36960 400 37016
rect 0 36848 400 36904
rect 0 36736 400 36792
rect 0 36624 400 36680
rect 0 36512 400 36568
rect 0 36400 400 36456
rect 0 36288 400 36344
rect 0 36176 400 36232
rect 0 36064 400 36120
rect 0 35952 400 36008
rect 0 35840 400 35896
rect 0 35728 400 35784
rect 0 35616 400 35672
rect 0 35504 400 35560
rect 0 35392 400 35448
rect 0 35280 400 35336
rect 0 35168 400 35224
rect 0 35056 400 35112
rect 0 34944 400 35000
rect 0 34832 400 34888
rect 0 34720 400 34776
rect 0 34608 400 34664
rect 0 34496 400 34552
rect 0 34384 400 34440
rect 0 34272 400 34328
rect 0 34160 400 34216
rect 0 34048 400 34104
rect 0 33936 400 33992
rect 0 33824 400 33880
rect 0 33712 400 33768
rect 0 33600 400 33656
rect 0 33488 400 33544
rect 0 33376 400 33432
rect 0 33264 400 33320
rect 0 33152 400 33208
rect 0 33040 400 33096
rect 0 32928 400 32984
rect 0 32816 400 32872
rect 0 32704 400 32760
rect 0 32592 400 32648
rect 0 32480 400 32536
rect 0 32368 400 32424
rect 0 32256 400 32312
rect 0 32144 400 32200
rect 0 32032 400 32088
rect 0 31920 400 31976
rect 0 31808 400 31864
rect 0 31696 400 31752
rect 0 31584 400 31640
rect 0 31472 400 31528
rect 0 31360 400 31416
rect 0 31248 400 31304
rect 0 31136 400 31192
rect 0 31024 400 31080
rect 0 30912 400 30968
rect 0 30800 400 30856
rect 0 30688 400 30744
rect 0 30576 400 30632
rect 0 30464 400 30520
rect 0 30352 400 30408
rect 0 30240 400 30296
rect 0 30128 400 30184
rect 0 30016 400 30072
rect 0 29904 400 29960
rect 0 29792 400 29848
rect 0 29680 400 29736
rect 0 29568 400 29624
rect 0 29456 400 29512
rect 0 29344 400 29400
rect 0 29232 400 29288
rect 0 29120 400 29176
rect 0 29008 400 29064
rect 0 28896 400 28952
rect 0 28784 400 28840
rect 0 28672 400 28728
rect 0 28560 400 28616
rect 0 28448 400 28504
rect 0 28336 400 28392
rect 0 28224 400 28280
rect 0 28112 400 28168
rect 0 28000 400 28056
rect 0 27888 400 27944
rect 0 27776 400 27832
rect 0 27664 400 27720
rect 0 27552 400 27608
rect 0 27440 400 27496
rect 0 27328 400 27384
rect 0 27216 400 27272
rect 0 27104 400 27160
rect 0 26992 400 27048
rect 0 26880 400 26936
rect 0 26768 400 26824
rect 0 26656 400 26712
rect 0 26544 400 26600
rect 0 26432 400 26488
rect 0 26320 400 26376
rect 0 26208 400 26264
rect 0 26096 400 26152
rect 0 25984 400 26040
rect 0 25872 400 25928
rect 0 25760 400 25816
rect 0 25648 400 25704
rect 0 25536 400 25592
rect 0 25424 400 25480
rect 0 25312 400 25368
rect 0 25200 400 25256
rect 0 25088 400 25144
rect 0 24976 400 25032
rect 0 24864 400 24920
rect 0 24752 400 24808
rect 0 24640 400 24696
rect 0 24528 400 24584
rect 0 24416 400 24472
rect 0 24304 400 24360
rect 0 24192 400 24248
rect 0 24080 400 24136
rect 0 23968 400 24024
rect 0 23856 400 23912
rect 0 23744 400 23800
rect 0 23632 400 23688
rect 0 23520 400 23576
rect 0 23408 400 23464
rect 0 23296 400 23352
rect 0 23184 400 23240
rect 0 23072 400 23128
rect 0 22960 400 23016
rect 0 22848 400 22904
rect 0 22736 400 22792
rect 0 22624 400 22680
rect 0 22512 400 22568
rect 0 22400 400 22456
rect 0 22288 400 22344
rect 0 22176 400 22232
rect 0 22064 400 22120
rect 0 21952 400 22008
rect 0 21840 400 21896
rect 0 21728 400 21784
rect 0 21616 400 21672
rect 0 21504 400 21560
rect 0 21392 400 21448
rect 0 21280 400 21336
rect 0 21168 400 21224
rect 0 21056 400 21112
rect 0 20944 400 21000
rect 0 20832 400 20888
rect 0 20720 400 20776
rect 0 20608 400 20664
rect 0 20496 400 20552
rect 0 20384 400 20440
rect 0 20272 400 20328
rect 0 20160 400 20216
rect 0 20048 400 20104
rect 0 19936 400 19992
rect 0 19824 400 19880
rect 0 19712 400 19768
rect 0 19600 400 19656
rect 0 19488 400 19544
rect 0 19376 400 19432
rect 0 19264 400 19320
rect 0 19152 400 19208
rect 0 19040 400 19096
rect 0 18928 400 18984
rect 0 18816 400 18872
rect 0 18704 400 18760
rect 0 18592 400 18648
rect 0 18480 400 18536
rect 0 18368 400 18424
rect 0 18256 400 18312
rect 0 18144 400 18200
rect 0 18032 400 18088
rect 0 17920 400 17976
rect 0 17808 400 17864
rect 0 17696 400 17752
rect 0 17584 400 17640
rect 0 17472 400 17528
rect 0 17360 400 17416
rect 0 17248 400 17304
rect 0 17136 400 17192
rect 0 17024 400 17080
rect 0 16912 400 16968
rect 0 16800 400 16856
rect 0 16688 400 16744
rect 0 16576 400 16632
rect 0 16464 400 16520
rect 0 16352 400 16408
rect 0 16240 400 16296
rect 0 16128 400 16184
rect 0 16016 400 16072
rect 0 15904 400 15960
rect 0 15792 400 15848
rect 0 15680 400 15736
rect 0 15568 400 15624
rect 0 15456 400 15512
rect 0 15344 400 15400
rect 0 15232 400 15288
rect 0 15120 400 15176
rect 0 15008 400 15064
rect 0 14896 400 14952
rect 0 14784 400 14840
rect 0 14672 400 14728
rect 0 14560 400 14616
rect 0 14448 400 14504
rect 0 14336 400 14392
rect 0 14224 400 14280
rect 0 14112 400 14168
rect 0 14000 400 14056
rect 0 13888 400 13944
rect 0 13776 400 13832
rect 0 13664 400 13720
rect 0 13552 400 13608
rect 0 13440 400 13496
rect 0 13328 400 13384
rect 0 13216 400 13272
rect 0 13104 400 13160
rect 0 12992 400 13048
rect 0 12880 400 12936
rect 0 12768 400 12824
rect 0 12656 400 12712
rect 0 12544 400 12600
rect 0 12432 400 12488
rect 0 12320 400 12376
rect 0 12208 400 12264
rect 0 12096 400 12152
rect 0 11984 400 12040
rect 0 11872 400 11928
rect 0 11760 400 11816
rect 0 11648 400 11704
rect 0 11536 400 11592
rect 0 11424 400 11480
rect 0 11312 400 11368
rect 0 11200 400 11256
rect 0 11088 400 11144
rect 0 10976 400 11032
rect 0 10864 400 10920
rect 0 10752 400 10808
rect 0 10640 400 10696
rect 0 10528 400 10584
rect 0 10416 400 10472
rect 0 10304 400 10360
rect 0 10192 400 10248
rect 0 10080 400 10136
rect 0 9968 400 10024
rect 279600 69888 280000 69944
rect 279600 69776 280000 69832
rect 279600 69664 280000 69720
rect 279600 69552 280000 69608
rect 279600 69440 280000 69496
rect 279600 69328 280000 69384
rect 279600 69216 280000 69272
rect 279600 69104 280000 69160
rect 279600 68992 280000 69048
rect 279600 68880 280000 68936
rect 279600 68768 280000 68824
rect 279600 68656 280000 68712
rect 279600 68544 280000 68600
rect 279600 68432 280000 68488
rect 279600 68320 280000 68376
rect 279600 68208 280000 68264
rect 279600 68096 280000 68152
rect 279600 67984 280000 68040
rect 279600 67872 280000 67928
rect 279600 67760 280000 67816
rect 279600 67648 280000 67704
rect 279600 67536 280000 67592
rect 279600 67424 280000 67480
rect 279600 67312 280000 67368
rect 279600 67200 280000 67256
rect 279600 67088 280000 67144
rect 279600 66976 280000 67032
rect 279600 66864 280000 66920
rect 279600 66752 280000 66808
rect 279600 66640 280000 66696
rect 279600 66528 280000 66584
rect 279600 66416 280000 66472
rect 279600 66304 280000 66360
rect 279600 66192 280000 66248
rect 279600 66080 280000 66136
rect 279600 65968 280000 66024
rect 279600 65856 280000 65912
rect 279600 65744 280000 65800
rect 279600 65632 280000 65688
rect 279600 65520 280000 65576
rect 279600 65408 280000 65464
rect 279600 65296 280000 65352
rect 279600 65184 280000 65240
rect 279600 65072 280000 65128
rect 279600 64960 280000 65016
rect 279600 64848 280000 64904
rect 279600 64736 280000 64792
rect 279600 64624 280000 64680
rect 279600 64512 280000 64568
rect 279600 64400 280000 64456
rect 279600 64288 280000 64344
rect 279600 64176 280000 64232
rect 279600 64064 280000 64120
rect 279600 63952 280000 64008
rect 279600 63840 280000 63896
rect 279600 63728 280000 63784
rect 279600 63616 280000 63672
rect 279600 63504 280000 63560
rect 279600 63392 280000 63448
rect 279600 63280 280000 63336
rect 279600 63168 280000 63224
rect 279600 63056 280000 63112
rect 279600 62944 280000 63000
rect 279600 62832 280000 62888
rect 279600 62720 280000 62776
rect 279600 62608 280000 62664
rect 279600 62496 280000 62552
rect 279600 62384 280000 62440
rect 279600 62272 280000 62328
rect 279600 62160 280000 62216
rect 279600 62048 280000 62104
rect 279600 61936 280000 61992
rect 279600 61824 280000 61880
rect 279600 61712 280000 61768
rect 279600 61600 280000 61656
rect 279600 61488 280000 61544
rect 279600 61376 280000 61432
rect 279600 61264 280000 61320
rect 279600 61152 280000 61208
rect 279600 61040 280000 61096
rect 279600 60928 280000 60984
rect 279600 60816 280000 60872
rect 279600 60704 280000 60760
rect 279600 60592 280000 60648
rect 279600 60480 280000 60536
rect 279600 60368 280000 60424
rect 279600 60256 280000 60312
rect 279600 60144 280000 60200
rect 279600 60032 280000 60088
rect 279600 59920 280000 59976
rect 279600 59808 280000 59864
rect 279600 59696 280000 59752
rect 279600 59584 280000 59640
rect 279600 59472 280000 59528
rect 279600 59360 280000 59416
rect 279600 59248 280000 59304
rect 279600 59136 280000 59192
rect 279600 59024 280000 59080
rect 279600 58912 280000 58968
rect 279600 58800 280000 58856
rect 279600 58688 280000 58744
rect 279600 58576 280000 58632
rect 279600 58464 280000 58520
rect 279600 58352 280000 58408
rect 279600 58240 280000 58296
rect 279600 58128 280000 58184
rect 279600 58016 280000 58072
rect 279600 57904 280000 57960
rect 279600 57792 280000 57848
rect 279600 57680 280000 57736
rect 279600 57568 280000 57624
rect 279600 57456 280000 57512
rect 279600 57344 280000 57400
rect 279600 57232 280000 57288
rect 279600 57120 280000 57176
rect 279600 57008 280000 57064
rect 279600 56896 280000 56952
rect 279600 56784 280000 56840
rect 279600 56672 280000 56728
rect 279600 56560 280000 56616
rect 279600 56448 280000 56504
rect 279600 56336 280000 56392
rect 279600 56224 280000 56280
rect 279600 56112 280000 56168
rect 279600 56000 280000 56056
rect 279600 55888 280000 55944
rect 279600 55776 280000 55832
rect 279600 55664 280000 55720
rect 279600 55552 280000 55608
rect 279600 55440 280000 55496
rect 279600 55328 280000 55384
rect 279600 55216 280000 55272
rect 279600 55104 280000 55160
rect 279600 54992 280000 55048
rect 279600 54880 280000 54936
rect 279600 54768 280000 54824
rect 279600 54656 280000 54712
rect 279600 54544 280000 54600
rect 279600 54432 280000 54488
rect 279600 54320 280000 54376
rect 279600 54208 280000 54264
rect 279600 54096 280000 54152
rect 279600 53984 280000 54040
rect 279600 53872 280000 53928
rect 279600 53760 280000 53816
rect 279600 53648 280000 53704
rect 279600 53536 280000 53592
rect 279600 53424 280000 53480
rect 279600 53312 280000 53368
rect 279600 53200 280000 53256
rect 279600 53088 280000 53144
rect 279600 52976 280000 53032
rect 279600 52864 280000 52920
rect 279600 52752 280000 52808
rect 279600 52640 280000 52696
rect 279600 52528 280000 52584
rect 279600 52416 280000 52472
rect 279600 52304 280000 52360
rect 279600 52192 280000 52248
rect 279600 52080 280000 52136
rect 279600 51968 280000 52024
rect 279600 51856 280000 51912
rect 279600 51744 280000 51800
rect 279600 51632 280000 51688
rect 279600 51520 280000 51576
rect 279600 51408 280000 51464
rect 279600 51296 280000 51352
rect 279600 51184 280000 51240
rect 279600 51072 280000 51128
rect 279600 50960 280000 51016
rect 279600 50848 280000 50904
rect 279600 50736 280000 50792
rect 279600 50624 280000 50680
rect 279600 50512 280000 50568
rect 279600 50400 280000 50456
rect 279600 50288 280000 50344
rect 279600 50176 280000 50232
rect 279600 50064 280000 50120
rect 279600 49952 280000 50008
rect 279600 49840 280000 49896
rect 279600 49728 280000 49784
rect 279600 49616 280000 49672
rect 279600 49504 280000 49560
rect 279600 49392 280000 49448
rect 279600 49280 280000 49336
rect 279600 49168 280000 49224
rect 279600 49056 280000 49112
rect 279600 48944 280000 49000
rect 279600 48832 280000 48888
rect 279600 48720 280000 48776
rect 279600 48608 280000 48664
rect 279600 48496 280000 48552
rect 279600 48384 280000 48440
rect 279600 48272 280000 48328
rect 279600 48160 280000 48216
rect 279600 48048 280000 48104
rect 279600 47936 280000 47992
rect 279600 47824 280000 47880
rect 279600 47712 280000 47768
rect 279600 47600 280000 47656
rect 279600 47488 280000 47544
rect 279600 47376 280000 47432
rect 279600 47264 280000 47320
rect 279600 47152 280000 47208
rect 279600 47040 280000 47096
rect 279600 46928 280000 46984
rect 279600 46816 280000 46872
rect 279600 46704 280000 46760
rect 279600 46592 280000 46648
rect 279600 46480 280000 46536
rect 279600 46368 280000 46424
rect 279600 46256 280000 46312
rect 279600 46144 280000 46200
rect 279600 46032 280000 46088
rect 279600 45920 280000 45976
rect 279600 45808 280000 45864
rect 279600 45696 280000 45752
rect 279600 45584 280000 45640
rect 279600 45472 280000 45528
rect 279600 45360 280000 45416
rect 279600 45248 280000 45304
rect 279600 45136 280000 45192
rect 279600 45024 280000 45080
rect 279600 44912 280000 44968
rect 279600 44800 280000 44856
rect 279600 44688 280000 44744
rect 279600 44576 280000 44632
rect 279600 44464 280000 44520
rect 279600 44352 280000 44408
rect 279600 44240 280000 44296
rect 279600 44128 280000 44184
rect 279600 44016 280000 44072
rect 279600 43904 280000 43960
rect 279600 43792 280000 43848
rect 279600 43680 280000 43736
rect 279600 43568 280000 43624
rect 279600 43456 280000 43512
rect 279600 43344 280000 43400
rect 279600 43232 280000 43288
rect 279600 43120 280000 43176
rect 279600 43008 280000 43064
rect 279600 42896 280000 42952
rect 279600 42784 280000 42840
rect 279600 42672 280000 42728
rect 279600 42560 280000 42616
rect 279600 42448 280000 42504
rect 279600 42336 280000 42392
rect 279600 42224 280000 42280
rect 279600 42112 280000 42168
rect 279600 42000 280000 42056
rect 279600 41888 280000 41944
rect 279600 41776 280000 41832
rect 279600 41664 280000 41720
rect 279600 41552 280000 41608
rect 279600 41440 280000 41496
rect 279600 41328 280000 41384
rect 279600 41216 280000 41272
rect 279600 41104 280000 41160
rect 279600 40992 280000 41048
rect 279600 40880 280000 40936
rect 279600 40768 280000 40824
rect 279600 40656 280000 40712
rect 279600 40544 280000 40600
rect 279600 40432 280000 40488
rect 279600 40320 280000 40376
rect 279600 40208 280000 40264
rect 279600 40096 280000 40152
rect 279600 39984 280000 40040
rect 279600 39872 280000 39928
rect 279600 39760 280000 39816
rect 279600 39648 280000 39704
rect 279600 39536 280000 39592
rect 279600 39424 280000 39480
rect 279600 39312 280000 39368
rect 279600 39200 280000 39256
rect 279600 39088 280000 39144
rect 279600 38976 280000 39032
rect 279600 38864 280000 38920
rect 279600 38752 280000 38808
rect 279600 38640 280000 38696
rect 279600 38528 280000 38584
rect 279600 38416 280000 38472
rect 279600 38304 280000 38360
rect 279600 38192 280000 38248
rect 279600 38080 280000 38136
rect 279600 37968 280000 38024
rect 279600 37856 280000 37912
rect 279600 37744 280000 37800
rect 279600 37632 280000 37688
rect 279600 37520 280000 37576
rect 279600 37408 280000 37464
rect 279600 37296 280000 37352
rect 279600 37184 280000 37240
rect 279600 37072 280000 37128
rect 279600 36960 280000 37016
rect 279600 36848 280000 36904
rect 279600 36736 280000 36792
rect 279600 36624 280000 36680
rect 279600 36512 280000 36568
rect 279600 36400 280000 36456
rect 279600 36288 280000 36344
rect 279600 36176 280000 36232
rect 279600 36064 280000 36120
rect 279600 35952 280000 36008
rect 279600 35840 280000 35896
rect 279600 35728 280000 35784
rect 279600 35616 280000 35672
rect 279600 35504 280000 35560
rect 279600 35392 280000 35448
rect 279600 35280 280000 35336
rect 279600 35168 280000 35224
rect 279600 35056 280000 35112
rect 279600 34944 280000 35000
rect 279600 34832 280000 34888
rect 279600 34720 280000 34776
rect 279600 34608 280000 34664
rect 279600 34496 280000 34552
rect 279600 34384 280000 34440
rect 279600 34272 280000 34328
rect 279600 34160 280000 34216
rect 279600 34048 280000 34104
rect 279600 33936 280000 33992
rect 279600 33824 280000 33880
rect 279600 33712 280000 33768
rect 279600 33600 280000 33656
rect 279600 33488 280000 33544
rect 279600 33376 280000 33432
rect 279600 33264 280000 33320
rect 279600 33152 280000 33208
rect 279600 33040 280000 33096
rect 279600 32928 280000 32984
rect 279600 32816 280000 32872
rect 279600 32704 280000 32760
rect 279600 32592 280000 32648
rect 279600 32480 280000 32536
rect 279600 32368 280000 32424
rect 279600 32256 280000 32312
rect 279600 32144 280000 32200
rect 279600 32032 280000 32088
rect 279600 31920 280000 31976
rect 279600 31808 280000 31864
rect 279600 31696 280000 31752
rect 279600 31584 280000 31640
rect 279600 31472 280000 31528
rect 279600 31360 280000 31416
rect 279600 31248 280000 31304
rect 279600 31136 280000 31192
rect 279600 31024 280000 31080
rect 279600 30912 280000 30968
rect 279600 30800 280000 30856
rect 279600 30688 280000 30744
rect 279600 30576 280000 30632
rect 279600 30464 280000 30520
rect 279600 30352 280000 30408
rect 279600 30240 280000 30296
rect 279600 30128 280000 30184
rect 279600 30016 280000 30072
rect 279600 29904 280000 29960
rect 279600 29792 280000 29848
rect 279600 29680 280000 29736
rect 279600 29568 280000 29624
rect 279600 29456 280000 29512
rect 279600 29344 280000 29400
rect 279600 29232 280000 29288
rect 279600 29120 280000 29176
rect 279600 29008 280000 29064
rect 279600 28896 280000 28952
rect 279600 28784 280000 28840
rect 279600 28672 280000 28728
rect 279600 28560 280000 28616
rect 279600 28448 280000 28504
rect 279600 28336 280000 28392
rect 279600 28224 280000 28280
rect 279600 28112 280000 28168
rect 279600 28000 280000 28056
rect 279600 27888 280000 27944
rect 279600 27776 280000 27832
rect 279600 27664 280000 27720
rect 279600 27552 280000 27608
rect 279600 27440 280000 27496
rect 279600 27328 280000 27384
rect 279600 27216 280000 27272
rect 279600 27104 280000 27160
rect 279600 26992 280000 27048
rect 279600 26880 280000 26936
rect 279600 26768 280000 26824
rect 279600 26656 280000 26712
rect 279600 26544 280000 26600
rect 279600 26432 280000 26488
rect 279600 26320 280000 26376
rect 279600 26208 280000 26264
rect 279600 26096 280000 26152
rect 279600 25984 280000 26040
rect 279600 25872 280000 25928
rect 279600 25760 280000 25816
rect 279600 25648 280000 25704
rect 279600 25536 280000 25592
rect 279600 25424 280000 25480
rect 279600 25312 280000 25368
rect 279600 25200 280000 25256
rect 279600 25088 280000 25144
rect 279600 24976 280000 25032
rect 279600 24864 280000 24920
rect 279600 24752 280000 24808
rect 279600 24640 280000 24696
rect 279600 24528 280000 24584
rect 279600 24416 280000 24472
rect 279600 24304 280000 24360
rect 279600 24192 280000 24248
rect 279600 24080 280000 24136
rect 279600 23968 280000 24024
rect 279600 23856 280000 23912
rect 279600 23744 280000 23800
rect 279600 23632 280000 23688
rect 279600 23520 280000 23576
rect 279600 23408 280000 23464
rect 279600 23296 280000 23352
rect 279600 23184 280000 23240
rect 279600 23072 280000 23128
rect 279600 22960 280000 23016
rect 279600 22848 280000 22904
rect 279600 22736 280000 22792
rect 279600 22624 280000 22680
rect 279600 22512 280000 22568
rect 279600 22400 280000 22456
rect 279600 22288 280000 22344
rect 279600 22176 280000 22232
rect 279600 22064 280000 22120
rect 279600 21952 280000 22008
rect 279600 21840 280000 21896
rect 279600 21728 280000 21784
rect 279600 21616 280000 21672
rect 279600 21504 280000 21560
rect 279600 21392 280000 21448
rect 279600 21280 280000 21336
rect 279600 21168 280000 21224
rect 279600 21056 280000 21112
rect 279600 20944 280000 21000
rect 279600 20832 280000 20888
rect 279600 20720 280000 20776
rect 279600 20608 280000 20664
rect 279600 20496 280000 20552
rect 279600 20384 280000 20440
rect 279600 20272 280000 20328
rect 279600 20160 280000 20216
rect 279600 20048 280000 20104
rect 279600 19936 280000 19992
rect 279600 19824 280000 19880
rect 279600 19712 280000 19768
rect 279600 19600 280000 19656
rect 279600 19488 280000 19544
rect 279600 19376 280000 19432
rect 279600 19264 280000 19320
rect 279600 19152 280000 19208
rect 279600 19040 280000 19096
rect 279600 18928 280000 18984
rect 279600 18816 280000 18872
rect 279600 18704 280000 18760
rect 279600 18592 280000 18648
rect 279600 18480 280000 18536
rect 279600 18368 280000 18424
rect 279600 18256 280000 18312
rect 279600 18144 280000 18200
rect 279600 18032 280000 18088
rect 279600 17920 280000 17976
rect 279600 17808 280000 17864
rect 279600 17696 280000 17752
rect 279600 17584 280000 17640
rect 279600 17472 280000 17528
rect 279600 17360 280000 17416
rect 279600 17248 280000 17304
rect 279600 17136 280000 17192
rect 279600 17024 280000 17080
rect 279600 16912 280000 16968
rect 279600 16800 280000 16856
rect 279600 16688 280000 16744
rect 279600 16576 280000 16632
rect 279600 16464 280000 16520
rect 279600 16352 280000 16408
rect 279600 16240 280000 16296
rect 279600 16128 280000 16184
rect 279600 16016 280000 16072
rect 279600 15904 280000 15960
rect 279600 15792 280000 15848
rect 279600 15680 280000 15736
rect 279600 15568 280000 15624
rect 279600 15456 280000 15512
rect 279600 15344 280000 15400
rect 279600 15232 280000 15288
rect 279600 15120 280000 15176
rect 279600 15008 280000 15064
rect 279600 14896 280000 14952
rect 279600 14784 280000 14840
rect 279600 14672 280000 14728
rect 279600 14560 280000 14616
rect 279600 14448 280000 14504
rect 279600 14336 280000 14392
rect 279600 14224 280000 14280
rect 279600 14112 280000 14168
rect 279600 14000 280000 14056
rect 279600 13888 280000 13944
rect 279600 13776 280000 13832
rect 279600 13664 280000 13720
rect 279600 13552 280000 13608
rect 279600 13440 280000 13496
rect 279600 13328 280000 13384
rect 279600 13216 280000 13272
rect 279600 13104 280000 13160
rect 279600 12992 280000 13048
rect 279600 12880 280000 12936
rect 279600 12768 280000 12824
rect 279600 12656 280000 12712
rect 279600 12544 280000 12600
rect 279600 12432 280000 12488
rect 279600 12320 280000 12376
rect 279600 12208 280000 12264
rect 279600 12096 280000 12152
rect 279600 11984 280000 12040
rect 279600 11872 280000 11928
rect 279600 11760 280000 11816
rect 279600 11648 280000 11704
rect 279600 11536 280000 11592
rect 279600 11424 280000 11480
rect 279600 11312 280000 11368
rect 279600 11200 280000 11256
rect 279600 11088 280000 11144
rect 279600 10976 280000 11032
rect 279600 10864 280000 10920
rect 279600 10752 280000 10808
rect 279600 10640 280000 10696
rect 279600 10528 280000 10584
rect 279600 10416 280000 10472
rect 279600 10304 280000 10360
rect 279600 10192 280000 10248
rect 279600 10080 280000 10136
rect 279600 9968 280000 10024
<< obsm3 >>
rect 400 69974 279600 79338
rect 430 9938 279570 69974
rect 400 1554 279600 9938
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
rect 71344 1538 71504 78430
rect 79024 1538 79184 78430
rect 86704 1538 86864 78430
rect 94384 1538 94544 78430
rect 102064 1538 102224 78430
rect 109744 1538 109904 78430
rect 117424 1538 117584 78430
rect 125104 1538 125264 78430
rect 132784 1538 132944 78430
rect 140464 1538 140624 78430
rect 148144 1538 148304 78430
rect 155824 1538 155984 78430
rect 163504 1538 163664 78430
rect 171184 1538 171344 78430
rect 178864 1538 179024 78430
rect 186544 1538 186704 78430
rect 194224 1538 194384 78430
rect 201904 1538 202064 78430
rect 209584 1538 209744 78430
rect 217264 1538 217424 78430
rect 224944 1538 225104 78430
rect 232624 1538 232784 78430
rect 240304 1538 240464 78430
rect 247984 1538 248144 78430
rect 255664 1538 255824 78430
rect 263344 1538 263504 78430
rect 271024 1538 271184 78430
rect 278704 1538 278864 78430
<< obsm4 >>
rect 77742 76393 78994 77439
rect 79214 76393 86674 77439
rect 86894 76393 94354 77439
rect 94574 76393 102034 77439
rect 102254 76393 109714 77439
rect 109934 76393 117394 77439
rect 117614 76393 125074 77439
rect 125294 76393 132754 77439
rect 132974 76393 140434 77439
rect 140654 76393 148114 77439
rect 148334 76393 155794 77439
rect 156014 76393 163474 77439
rect 163694 76393 171154 77439
rect 171374 76393 174762 77439
<< labels >>
rlabel metal2 s 276080 79600 276136 80000 6 gpu_clk
port 1 nsew signal input
rlabel metal3 s 279600 9968 280000 10024 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 69216 400 69272 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 0 68880 400 68936 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 0 68544 400 68600 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 0 68208 400 68264 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 0 67872 400 67928 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 0 67536 400 67592 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 279600 10304 280000 10360 6 io_in[1]
port 9 nsew signal input
rlabel metal3 s 279600 10640 280000 10696 6 io_in[2]
port 10 nsew signal input
rlabel metal3 s 279600 10976 280000 11032 6 io_in[3]
port 11 nsew signal input
rlabel metal3 s 279600 11312 280000 11368 6 io_in[4]
port 12 nsew signal input
rlabel metal3 s 279600 11648 280000 11704 6 io_in[5]
port 13 nsew signal input
rlabel metal3 s 279600 11984 280000 12040 6 io_in[6]
port 14 nsew signal input
rlabel metal3 s 279600 12320 280000 12376 6 io_in[7]
port 15 nsew signal input
rlabel metal3 s 0 69888 400 69944 6 io_in[8]
port 16 nsew signal input
rlabel metal3 s 0 69552 400 69608 6 io_in[9]
port 17 nsew signal input
rlabel metal3 s 279600 10192 280000 10248 6 io_oeb[0]
port 18 nsew signal output
rlabel metal3 s 0 68992 400 69048 6 io_oeb[10]
port 19 nsew signal output
rlabel metal3 s 0 68656 400 68712 6 io_oeb[11]
port 20 nsew signal output
rlabel metal3 s 0 68320 400 68376 6 io_oeb[12]
port 21 nsew signal output
rlabel metal3 s 0 67984 400 68040 6 io_oeb[13]
port 22 nsew signal output
rlabel metal3 s 0 67648 400 67704 6 io_oeb[14]
port 23 nsew signal output
rlabel metal3 s 0 67312 400 67368 6 io_oeb[15]
port 24 nsew signal output
rlabel metal3 s 279600 10528 280000 10584 6 io_oeb[1]
port 25 nsew signal output
rlabel metal3 s 279600 10864 280000 10920 6 io_oeb[2]
port 26 nsew signal output
rlabel metal3 s 279600 11200 280000 11256 6 io_oeb[3]
port 27 nsew signal output
rlabel metal3 s 279600 11536 280000 11592 6 io_oeb[4]
port 28 nsew signal output
rlabel metal3 s 279600 11872 280000 11928 6 io_oeb[5]
port 29 nsew signal output
rlabel metal3 s 279600 12208 280000 12264 6 io_oeb[6]
port 30 nsew signal output
rlabel metal3 s 279600 12544 280000 12600 6 io_oeb[7]
port 31 nsew signal output
rlabel metal3 s 0 69664 400 69720 6 io_oeb[8]
port 32 nsew signal output
rlabel metal3 s 0 69328 400 69384 6 io_oeb[9]
port 33 nsew signal output
rlabel metal3 s 279600 10080 280000 10136 6 io_out[0]
port 34 nsew signal output
rlabel metal3 s 0 69104 400 69160 6 io_out[10]
port 35 nsew signal output
rlabel metal3 s 0 68768 400 68824 6 io_out[11]
port 36 nsew signal output
rlabel metal3 s 0 68432 400 68488 6 io_out[12]
port 37 nsew signal output
rlabel metal3 s 0 68096 400 68152 6 io_out[13]
port 38 nsew signal output
rlabel metal3 s 0 67760 400 67816 6 io_out[14]
port 39 nsew signal output
rlabel metal3 s 0 67424 400 67480 6 io_out[15]
port 40 nsew signal output
rlabel metal3 s 279600 10416 280000 10472 6 io_out[1]
port 41 nsew signal output
rlabel metal3 s 279600 10752 280000 10808 6 io_out[2]
port 42 nsew signal output
rlabel metal3 s 279600 11088 280000 11144 6 io_out[3]
port 43 nsew signal output
rlabel metal3 s 279600 11424 280000 11480 6 io_out[4]
port 44 nsew signal output
rlabel metal3 s 279600 11760 280000 11816 6 io_out[5]
port 45 nsew signal output
rlabel metal3 s 279600 12096 280000 12152 6 io_out[6]
port 46 nsew signal output
rlabel metal3 s 279600 12432 280000 12488 6 io_out[7]
port 47 nsew signal output
rlabel metal3 s 0 69776 400 69832 6 io_out[8]
port 48 nsew signal output
rlabel metal3 s 0 69440 400 69496 6 io_out[9]
port 49 nsew signal output
rlabel metal2 s 103600 0 103656 400 6 irq[0]
port 50 nsew signal output
rlabel metal2 s 103936 0 103992 400 6 irq[1]
port 51 nsew signal output
rlabel metal2 s 104272 0 104328 400 6 irq[2]
port 52 nsew signal output
rlabel metal2 s 39088 0 39144 400 6 la_data_in[0]
port 53 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 la_data_in[10]
port 54 nsew signal input
rlabel metal2 s 50176 0 50232 400 6 la_data_in[11]
port 55 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 la_data_in[12]
port 56 nsew signal input
rlabel metal2 s 52192 0 52248 400 6 la_data_in[13]
port 57 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 la_data_in[14]
port 58 nsew signal input
rlabel metal2 s 54208 0 54264 400 6 la_data_in[15]
port 59 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 la_data_in[16]
port 60 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 la_data_in[17]
port 61 nsew signal input
rlabel metal2 s 57232 0 57288 400 6 la_data_in[18]
port 62 nsew signal input
rlabel metal2 s 58240 0 58296 400 6 la_data_in[19]
port 63 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 la_data_in[1]
port 64 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_data_in[20]
port 65 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 la_data_in[21]
port 66 nsew signal input
rlabel metal2 s 61264 0 61320 400 6 la_data_in[22]
port 67 nsew signal input
rlabel metal2 s 62272 0 62328 400 6 la_data_in[23]
port 68 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 la_data_in[24]
port 69 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 la_data_in[25]
port 70 nsew signal input
rlabel metal2 s 65296 0 65352 400 6 la_data_in[26]
port 71 nsew signal input
rlabel metal2 s 66304 0 66360 400 6 la_data_in[27]
port 72 nsew signal input
rlabel metal2 s 67312 0 67368 400 6 la_data_in[28]
port 73 nsew signal input
rlabel metal2 s 68320 0 68376 400 6 la_data_in[29]
port 74 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 la_data_in[2]
port 75 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_data_in[30]
port 76 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 la_data_in[31]
port 77 nsew signal input
rlabel metal2 s 71344 0 71400 400 6 la_data_in[32]
port 78 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 la_data_in[33]
port 79 nsew signal input
rlabel metal2 s 73360 0 73416 400 6 la_data_in[34]
port 80 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 la_data_in[35]
port 81 nsew signal input
rlabel metal2 s 75376 0 75432 400 6 la_data_in[36]
port 82 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 la_data_in[37]
port 83 nsew signal input
rlabel metal2 s 77392 0 77448 400 6 la_data_in[38]
port 84 nsew signal input
rlabel metal2 s 78400 0 78456 400 6 la_data_in[39]
port 85 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 la_data_in[3]
port 86 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_data_in[40]
port 87 nsew signal input
rlabel metal2 s 80416 0 80472 400 6 la_data_in[41]
port 88 nsew signal input
rlabel metal2 s 81424 0 81480 400 6 la_data_in[42]
port 89 nsew signal input
rlabel metal2 s 82432 0 82488 400 6 la_data_in[43]
port 90 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 la_data_in[44]
port 91 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 la_data_in[45]
port 92 nsew signal input
rlabel metal2 s 85456 0 85512 400 6 la_data_in[46]
port 93 nsew signal input
rlabel metal2 s 86464 0 86520 400 6 la_data_in[47]
port 94 nsew signal input
rlabel metal2 s 87472 0 87528 400 6 la_data_in[48]
port 95 nsew signal input
rlabel metal2 s 88480 0 88536 400 6 la_data_in[49]
port 96 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 la_data_in[4]
port 97 nsew signal input
rlabel metal2 s 89488 0 89544 400 6 la_data_in[50]
port 98 nsew signal input
rlabel metal2 s 90496 0 90552 400 6 la_data_in[51]
port 99 nsew signal input
rlabel metal2 s 91504 0 91560 400 6 la_data_in[52]
port 100 nsew signal input
rlabel metal2 s 92512 0 92568 400 6 la_data_in[53]
port 101 nsew signal input
rlabel metal2 s 93520 0 93576 400 6 la_data_in[54]
port 102 nsew signal input
rlabel metal2 s 94528 0 94584 400 6 la_data_in[55]
port 103 nsew signal input
rlabel metal2 s 95536 0 95592 400 6 la_data_in[56]
port 104 nsew signal input
rlabel metal2 s 96544 0 96600 400 6 la_data_in[57]
port 105 nsew signal input
rlabel metal2 s 97552 0 97608 400 6 la_data_in[58]
port 106 nsew signal input
rlabel metal2 s 98560 0 98616 400 6 la_data_in[59]
port 107 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 la_data_in[5]
port 108 nsew signal input
rlabel metal2 s 99568 0 99624 400 6 la_data_in[60]
port 109 nsew signal input
rlabel metal2 s 100576 0 100632 400 6 la_data_in[61]
port 110 nsew signal input
rlabel metal2 s 101584 0 101640 400 6 la_data_in[62]
port 111 nsew signal input
rlabel metal2 s 102592 0 102648 400 6 la_data_in[63]
port 112 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 la_data_in[6]
port 113 nsew signal input
rlabel metal2 s 46144 0 46200 400 6 la_data_in[7]
port 114 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 la_data_in[8]
port 115 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 la_data_in[9]
port 116 nsew signal input
rlabel metal2 s 39424 0 39480 400 6 la_data_out[0]
port 117 nsew signal output
rlabel metal2 s 49504 0 49560 400 6 la_data_out[10]
port 118 nsew signal output
rlabel metal2 s 50512 0 50568 400 6 la_data_out[11]
port 119 nsew signal output
rlabel metal2 s 51520 0 51576 400 6 la_data_out[12]
port 120 nsew signal output
rlabel metal2 s 52528 0 52584 400 6 la_data_out[13]
port 121 nsew signal output
rlabel metal2 s 53536 0 53592 400 6 la_data_out[14]
port 122 nsew signal output
rlabel metal2 s 54544 0 54600 400 6 la_data_out[15]
port 123 nsew signal output
rlabel metal2 s 55552 0 55608 400 6 la_data_out[16]
port 124 nsew signal output
rlabel metal2 s 56560 0 56616 400 6 la_data_out[17]
port 125 nsew signal output
rlabel metal2 s 57568 0 57624 400 6 la_data_out[18]
port 126 nsew signal output
rlabel metal2 s 58576 0 58632 400 6 la_data_out[19]
port 127 nsew signal output
rlabel metal2 s 40432 0 40488 400 6 la_data_out[1]
port 128 nsew signal output
rlabel metal2 s 59584 0 59640 400 6 la_data_out[20]
port 129 nsew signal output
rlabel metal2 s 60592 0 60648 400 6 la_data_out[21]
port 130 nsew signal output
rlabel metal2 s 61600 0 61656 400 6 la_data_out[22]
port 131 nsew signal output
rlabel metal2 s 62608 0 62664 400 6 la_data_out[23]
port 132 nsew signal output
rlabel metal2 s 63616 0 63672 400 6 la_data_out[24]
port 133 nsew signal output
rlabel metal2 s 64624 0 64680 400 6 la_data_out[25]
port 134 nsew signal output
rlabel metal2 s 65632 0 65688 400 6 la_data_out[26]
port 135 nsew signal output
rlabel metal2 s 66640 0 66696 400 6 la_data_out[27]
port 136 nsew signal output
rlabel metal2 s 67648 0 67704 400 6 la_data_out[28]
port 137 nsew signal output
rlabel metal2 s 68656 0 68712 400 6 la_data_out[29]
port 138 nsew signal output
rlabel metal2 s 41440 0 41496 400 6 la_data_out[2]
port 139 nsew signal output
rlabel metal2 s 69664 0 69720 400 6 la_data_out[30]
port 140 nsew signal output
rlabel metal2 s 70672 0 70728 400 6 la_data_out[31]
port 141 nsew signal output
rlabel metal2 s 71680 0 71736 400 6 la_data_out[32]
port 142 nsew signal output
rlabel metal2 s 72688 0 72744 400 6 la_data_out[33]
port 143 nsew signal output
rlabel metal2 s 73696 0 73752 400 6 la_data_out[34]
port 144 nsew signal output
rlabel metal2 s 74704 0 74760 400 6 la_data_out[35]
port 145 nsew signal output
rlabel metal2 s 75712 0 75768 400 6 la_data_out[36]
port 146 nsew signal output
rlabel metal2 s 76720 0 76776 400 6 la_data_out[37]
port 147 nsew signal output
rlabel metal2 s 77728 0 77784 400 6 la_data_out[38]
port 148 nsew signal output
rlabel metal2 s 78736 0 78792 400 6 la_data_out[39]
port 149 nsew signal output
rlabel metal2 s 42448 0 42504 400 6 la_data_out[3]
port 150 nsew signal output
rlabel metal2 s 79744 0 79800 400 6 la_data_out[40]
port 151 nsew signal output
rlabel metal2 s 80752 0 80808 400 6 la_data_out[41]
port 152 nsew signal output
rlabel metal2 s 81760 0 81816 400 6 la_data_out[42]
port 153 nsew signal output
rlabel metal2 s 82768 0 82824 400 6 la_data_out[43]
port 154 nsew signal output
rlabel metal2 s 83776 0 83832 400 6 la_data_out[44]
port 155 nsew signal output
rlabel metal2 s 84784 0 84840 400 6 la_data_out[45]
port 156 nsew signal output
rlabel metal2 s 85792 0 85848 400 6 la_data_out[46]
port 157 nsew signal output
rlabel metal2 s 86800 0 86856 400 6 la_data_out[47]
port 158 nsew signal output
rlabel metal2 s 87808 0 87864 400 6 la_data_out[48]
port 159 nsew signal output
rlabel metal2 s 88816 0 88872 400 6 la_data_out[49]
port 160 nsew signal output
rlabel metal2 s 43456 0 43512 400 6 la_data_out[4]
port 161 nsew signal output
rlabel metal2 s 89824 0 89880 400 6 la_data_out[50]
port 162 nsew signal output
rlabel metal2 s 90832 0 90888 400 6 la_data_out[51]
port 163 nsew signal output
rlabel metal2 s 91840 0 91896 400 6 la_data_out[52]
port 164 nsew signal output
rlabel metal2 s 92848 0 92904 400 6 la_data_out[53]
port 165 nsew signal output
rlabel metal2 s 93856 0 93912 400 6 la_data_out[54]
port 166 nsew signal output
rlabel metal2 s 94864 0 94920 400 6 la_data_out[55]
port 167 nsew signal output
rlabel metal2 s 95872 0 95928 400 6 la_data_out[56]
port 168 nsew signal output
rlabel metal2 s 96880 0 96936 400 6 la_data_out[57]
port 169 nsew signal output
rlabel metal2 s 97888 0 97944 400 6 la_data_out[58]
port 170 nsew signal output
rlabel metal2 s 98896 0 98952 400 6 la_data_out[59]
port 171 nsew signal output
rlabel metal2 s 44464 0 44520 400 6 la_data_out[5]
port 172 nsew signal output
rlabel metal2 s 99904 0 99960 400 6 la_data_out[60]
port 173 nsew signal output
rlabel metal2 s 100912 0 100968 400 6 la_data_out[61]
port 174 nsew signal output
rlabel metal2 s 101920 0 101976 400 6 la_data_out[62]
port 175 nsew signal output
rlabel metal2 s 102928 0 102984 400 6 la_data_out[63]
port 176 nsew signal output
rlabel metal2 s 45472 0 45528 400 6 la_data_out[6]
port 177 nsew signal output
rlabel metal2 s 46480 0 46536 400 6 la_data_out[7]
port 178 nsew signal output
rlabel metal2 s 47488 0 47544 400 6 la_data_out[8]
port 179 nsew signal output
rlabel metal2 s 48496 0 48552 400 6 la_data_out[9]
port 180 nsew signal output
rlabel metal2 s 39760 0 39816 400 6 la_oenb[0]
port 181 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 la_oenb[10]
port 182 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 la_oenb[11]
port 183 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 la_oenb[12]
port 184 nsew signal input
rlabel metal2 s 52864 0 52920 400 6 la_oenb[13]
port 185 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 la_oenb[14]
port 186 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 la_oenb[15]
port 187 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 la_oenb[16]
port 188 nsew signal input
rlabel metal2 s 56896 0 56952 400 6 la_oenb[17]
port 189 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 la_oenb[18]
port 190 nsew signal input
rlabel metal2 s 58912 0 58968 400 6 la_oenb[19]
port 191 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 la_oenb[1]
port 192 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 la_oenb[20]
port 193 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 la_oenb[21]
port 194 nsew signal input
rlabel metal2 s 61936 0 61992 400 6 la_oenb[22]
port 195 nsew signal input
rlabel metal2 s 62944 0 63000 400 6 la_oenb[23]
port 196 nsew signal input
rlabel metal2 s 63952 0 64008 400 6 la_oenb[24]
port 197 nsew signal input
rlabel metal2 s 64960 0 65016 400 6 la_oenb[25]
port 198 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 la_oenb[26]
port 199 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 la_oenb[27]
port 200 nsew signal input
rlabel metal2 s 67984 0 68040 400 6 la_oenb[28]
port 201 nsew signal input
rlabel metal2 s 68992 0 69048 400 6 la_oenb[29]
port 202 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 la_oenb[2]
port 203 nsew signal input
rlabel metal2 s 70000 0 70056 400 6 la_oenb[30]
port 204 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 la_oenb[31]
port 205 nsew signal input
rlabel metal2 s 72016 0 72072 400 6 la_oenb[32]
port 206 nsew signal input
rlabel metal2 s 73024 0 73080 400 6 la_oenb[33]
port 207 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 la_oenb[34]
port 208 nsew signal input
rlabel metal2 s 75040 0 75096 400 6 la_oenb[35]
port 209 nsew signal input
rlabel metal2 s 76048 0 76104 400 6 la_oenb[36]
port 210 nsew signal input
rlabel metal2 s 77056 0 77112 400 6 la_oenb[37]
port 211 nsew signal input
rlabel metal2 s 78064 0 78120 400 6 la_oenb[38]
port 212 nsew signal input
rlabel metal2 s 79072 0 79128 400 6 la_oenb[39]
port 213 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 la_oenb[3]
port 214 nsew signal input
rlabel metal2 s 80080 0 80136 400 6 la_oenb[40]
port 215 nsew signal input
rlabel metal2 s 81088 0 81144 400 6 la_oenb[41]
port 216 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 la_oenb[42]
port 217 nsew signal input
rlabel metal2 s 83104 0 83160 400 6 la_oenb[43]
port 218 nsew signal input
rlabel metal2 s 84112 0 84168 400 6 la_oenb[44]
port 219 nsew signal input
rlabel metal2 s 85120 0 85176 400 6 la_oenb[45]
port 220 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 la_oenb[46]
port 221 nsew signal input
rlabel metal2 s 87136 0 87192 400 6 la_oenb[47]
port 222 nsew signal input
rlabel metal2 s 88144 0 88200 400 6 la_oenb[48]
port 223 nsew signal input
rlabel metal2 s 89152 0 89208 400 6 la_oenb[49]
port 224 nsew signal input
rlabel metal2 s 43792 0 43848 400 6 la_oenb[4]
port 225 nsew signal input
rlabel metal2 s 90160 0 90216 400 6 la_oenb[50]
port 226 nsew signal input
rlabel metal2 s 91168 0 91224 400 6 la_oenb[51]
port 227 nsew signal input
rlabel metal2 s 92176 0 92232 400 6 la_oenb[52]
port 228 nsew signal input
rlabel metal2 s 93184 0 93240 400 6 la_oenb[53]
port 229 nsew signal input
rlabel metal2 s 94192 0 94248 400 6 la_oenb[54]
port 230 nsew signal input
rlabel metal2 s 95200 0 95256 400 6 la_oenb[55]
port 231 nsew signal input
rlabel metal2 s 96208 0 96264 400 6 la_oenb[56]
port 232 nsew signal input
rlabel metal2 s 97216 0 97272 400 6 la_oenb[57]
port 233 nsew signal input
rlabel metal2 s 98224 0 98280 400 6 la_oenb[58]
port 234 nsew signal input
rlabel metal2 s 99232 0 99288 400 6 la_oenb[59]
port 235 nsew signal input
rlabel metal2 s 44800 0 44856 400 6 la_oenb[5]
port 236 nsew signal input
rlabel metal2 s 100240 0 100296 400 6 la_oenb[60]
port 237 nsew signal input
rlabel metal2 s 101248 0 101304 400 6 la_oenb[61]
port 238 nsew signal input
rlabel metal2 s 102256 0 102312 400 6 la_oenb[62]
port 239 nsew signal input
rlabel metal2 s 103264 0 103320 400 6 la_oenb[63]
port 240 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 la_oenb[6]
port 241 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 la_oenb[7]
port 242 nsew signal input
rlabel metal2 s 47824 0 47880 400 6 la_oenb[8]
port 243 nsew signal input
rlabel metal2 s 48832 0 48888 400 6 la_oenb[9]
port 244 nsew signal input
rlabel metal2 s 137760 79600 137816 80000 6 tri_wbs_ack_o[0]
port 245 nsew signal input
rlabel metal2 s 116480 79600 116536 80000 6 tri_wbs_ack_o[10]
port 246 nsew signal input
rlabel metal2 s 114352 79600 114408 80000 6 tri_wbs_ack_o[11]
port 247 nsew signal input
rlabel metal2 s 112224 79600 112280 80000 6 tri_wbs_ack_o[12]
port 248 nsew signal input
rlabel metal2 s 110096 79600 110152 80000 6 tri_wbs_ack_o[13]
port 249 nsew signal input
rlabel metal2 s 107968 79600 108024 80000 6 tri_wbs_ack_o[14]
port 250 nsew signal input
rlabel metal2 s 105840 79600 105896 80000 6 tri_wbs_ack_o[15]
port 251 nsew signal input
rlabel metal2 s 103712 79600 103768 80000 6 tri_wbs_ack_o[16]
port 252 nsew signal input
rlabel metal2 s 101584 79600 101640 80000 6 tri_wbs_ack_o[17]
port 253 nsew signal input
rlabel metal2 s 99456 79600 99512 80000 6 tri_wbs_ack_o[18]
port 254 nsew signal input
rlabel metal2 s 97328 79600 97384 80000 6 tri_wbs_ack_o[19]
port 255 nsew signal input
rlabel metal2 s 135632 79600 135688 80000 6 tri_wbs_ack_o[1]
port 256 nsew signal input
rlabel metal2 s 95200 79600 95256 80000 6 tri_wbs_ack_o[20]
port 257 nsew signal input
rlabel metal2 s 93072 79600 93128 80000 6 tri_wbs_ack_o[21]
port 258 nsew signal input
rlabel metal2 s 90944 79600 91000 80000 6 tri_wbs_ack_o[22]
port 259 nsew signal input
rlabel metal2 s 88816 79600 88872 80000 6 tri_wbs_ack_o[23]
port 260 nsew signal input
rlabel metal2 s 86688 79600 86744 80000 6 tri_wbs_ack_o[24]
port 261 nsew signal input
rlabel metal2 s 84560 79600 84616 80000 6 tri_wbs_ack_o[25]
port 262 nsew signal input
rlabel metal2 s 82432 79600 82488 80000 6 tri_wbs_ack_o[26]
port 263 nsew signal input
rlabel metal2 s 80304 79600 80360 80000 6 tri_wbs_ack_o[27]
port 264 nsew signal input
rlabel metal2 s 78176 79600 78232 80000 6 tri_wbs_ack_o[28]
port 265 nsew signal input
rlabel metal2 s 76048 79600 76104 80000 6 tri_wbs_ack_o[29]
port 266 nsew signal input
rlabel metal2 s 133504 79600 133560 80000 6 tri_wbs_ack_o[2]
port 267 nsew signal input
rlabel metal2 s 73920 79600 73976 80000 6 tri_wbs_ack_o[30]
port 268 nsew signal input
rlabel metal2 s 71792 79600 71848 80000 6 tri_wbs_ack_o[31]
port 269 nsew signal input
rlabel metal2 s 69664 79600 69720 80000 6 tri_wbs_ack_o[32]
port 270 nsew signal input
rlabel metal2 s 67536 79600 67592 80000 6 tri_wbs_ack_o[33]
port 271 nsew signal input
rlabel metal2 s 65408 79600 65464 80000 6 tri_wbs_ack_o[34]
port 272 nsew signal input
rlabel metal2 s 63280 79600 63336 80000 6 tri_wbs_ack_o[35]
port 273 nsew signal input
rlabel metal2 s 61152 79600 61208 80000 6 tri_wbs_ack_o[36]
port 274 nsew signal input
rlabel metal2 s 59024 79600 59080 80000 6 tri_wbs_ack_o[37]
port 275 nsew signal input
rlabel metal2 s 56896 79600 56952 80000 6 tri_wbs_ack_o[38]
port 276 nsew signal input
rlabel metal2 s 54768 79600 54824 80000 6 tri_wbs_ack_o[39]
port 277 nsew signal input
rlabel metal2 s 131376 79600 131432 80000 6 tri_wbs_ack_o[3]
port 278 nsew signal input
rlabel metal2 s 52640 79600 52696 80000 6 tri_wbs_ack_o[40]
port 279 nsew signal input
rlabel metal2 s 50512 79600 50568 80000 6 tri_wbs_ack_o[41]
port 280 nsew signal input
rlabel metal2 s 48384 79600 48440 80000 6 tri_wbs_ack_o[42]
port 281 nsew signal input
rlabel metal2 s 46256 79600 46312 80000 6 tri_wbs_ack_o[43]
port 282 nsew signal input
rlabel metal2 s 44128 79600 44184 80000 6 tri_wbs_ack_o[44]
port 283 nsew signal input
rlabel metal2 s 42000 79600 42056 80000 6 tri_wbs_ack_o[45]
port 284 nsew signal input
rlabel metal2 s 39872 79600 39928 80000 6 tri_wbs_ack_o[46]
port 285 nsew signal input
rlabel metal2 s 37744 79600 37800 80000 6 tri_wbs_ack_o[47]
port 286 nsew signal input
rlabel metal2 s 35616 79600 35672 80000 6 tri_wbs_ack_o[48]
port 287 nsew signal input
rlabel metal2 s 33488 79600 33544 80000 6 tri_wbs_ack_o[49]
port 288 nsew signal input
rlabel metal2 s 129248 79600 129304 80000 6 tri_wbs_ack_o[4]
port 289 nsew signal input
rlabel metal2 s 31360 79600 31416 80000 6 tri_wbs_ack_o[50]
port 290 nsew signal input
rlabel metal2 s 29232 79600 29288 80000 6 tri_wbs_ack_o[51]
port 291 nsew signal input
rlabel metal2 s 27104 79600 27160 80000 6 tri_wbs_ack_o[52]
port 292 nsew signal input
rlabel metal2 s 24976 79600 25032 80000 6 tri_wbs_ack_o[53]
port 293 nsew signal input
rlabel metal2 s 22848 79600 22904 80000 6 tri_wbs_ack_o[54]
port 294 nsew signal input
rlabel metal2 s 20720 79600 20776 80000 6 tri_wbs_ack_o[55]
port 295 nsew signal input
rlabel metal2 s 18592 79600 18648 80000 6 tri_wbs_ack_o[56]
port 296 nsew signal input
rlabel metal2 s 16464 79600 16520 80000 6 tri_wbs_ack_o[57]
port 297 nsew signal input
rlabel metal2 s 14336 79600 14392 80000 6 tri_wbs_ack_o[58]
port 298 nsew signal input
rlabel metal2 s 12208 79600 12264 80000 6 tri_wbs_ack_o[59]
port 299 nsew signal input
rlabel metal2 s 127120 79600 127176 80000 6 tri_wbs_ack_o[5]
port 300 nsew signal input
rlabel metal2 s 10080 79600 10136 80000 6 tri_wbs_ack_o[60]
port 301 nsew signal input
rlabel metal2 s 7952 79600 8008 80000 6 tri_wbs_ack_o[61]
port 302 nsew signal input
rlabel metal2 s 5824 79600 5880 80000 6 tri_wbs_ack_o[62]
port 303 nsew signal input
rlabel metal2 s 3696 79600 3752 80000 6 tri_wbs_ack_o[63]
port 304 nsew signal input
rlabel metal2 s 124992 79600 125048 80000 6 tri_wbs_ack_o[6]
port 305 nsew signal input
rlabel metal2 s 122864 79600 122920 80000 6 tri_wbs_ack_o[7]
port 306 nsew signal input
rlabel metal2 s 120736 79600 120792 80000 6 tri_wbs_ack_o[8]
port 307 nsew signal input
rlabel metal2 s 118608 79600 118664 80000 6 tri_wbs_ack_o[9]
port 308 nsew signal input
rlabel metal2 s 273952 79600 274008 80000 6 tri_wbs_stb_i[0]
port 309 nsew signal output
rlabel metal2 s 252672 79600 252728 80000 6 tri_wbs_stb_i[10]
port 310 nsew signal output
rlabel metal2 s 250544 79600 250600 80000 6 tri_wbs_stb_i[11]
port 311 nsew signal output
rlabel metal2 s 248416 79600 248472 80000 6 tri_wbs_stb_i[12]
port 312 nsew signal output
rlabel metal2 s 246288 79600 246344 80000 6 tri_wbs_stb_i[13]
port 313 nsew signal output
rlabel metal2 s 244160 79600 244216 80000 6 tri_wbs_stb_i[14]
port 314 nsew signal output
rlabel metal2 s 242032 79600 242088 80000 6 tri_wbs_stb_i[15]
port 315 nsew signal output
rlabel metal2 s 239904 79600 239960 80000 6 tri_wbs_stb_i[16]
port 316 nsew signal output
rlabel metal2 s 237776 79600 237832 80000 6 tri_wbs_stb_i[17]
port 317 nsew signal output
rlabel metal2 s 235648 79600 235704 80000 6 tri_wbs_stb_i[18]
port 318 nsew signal output
rlabel metal2 s 233520 79600 233576 80000 6 tri_wbs_stb_i[19]
port 319 nsew signal output
rlabel metal2 s 271824 79600 271880 80000 6 tri_wbs_stb_i[1]
port 320 nsew signal output
rlabel metal2 s 231392 79600 231448 80000 6 tri_wbs_stb_i[20]
port 321 nsew signal output
rlabel metal2 s 229264 79600 229320 80000 6 tri_wbs_stb_i[21]
port 322 nsew signal output
rlabel metal2 s 227136 79600 227192 80000 6 tri_wbs_stb_i[22]
port 323 nsew signal output
rlabel metal2 s 225008 79600 225064 80000 6 tri_wbs_stb_i[23]
port 324 nsew signal output
rlabel metal2 s 222880 79600 222936 80000 6 tri_wbs_stb_i[24]
port 325 nsew signal output
rlabel metal2 s 220752 79600 220808 80000 6 tri_wbs_stb_i[25]
port 326 nsew signal output
rlabel metal2 s 218624 79600 218680 80000 6 tri_wbs_stb_i[26]
port 327 nsew signal output
rlabel metal2 s 216496 79600 216552 80000 6 tri_wbs_stb_i[27]
port 328 nsew signal output
rlabel metal2 s 214368 79600 214424 80000 6 tri_wbs_stb_i[28]
port 329 nsew signal output
rlabel metal2 s 212240 79600 212296 80000 6 tri_wbs_stb_i[29]
port 330 nsew signal output
rlabel metal2 s 269696 79600 269752 80000 6 tri_wbs_stb_i[2]
port 331 nsew signal output
rlabel metal2 s 210112 79600 210168 80000 6 tri_wbs_stb_i[30]
port 332 nsew signal output
rlabel metal2 s 207984 79600 208040 80000 6 tri_wbs_stb_i[31]
port 333 nsew signal output
rlabel metal2 s 205856 79600 205912 80000 6 tri_wbs_stb_i[32]
port 334 nsew signal output
rlabel metal2 s 203728 79600 203784 80000 6 tri_wbs_stb_i[33]
port 335 nsew signal output
rlabel metal2 s 201600 79600 201656 80000 6 tri_wbs_stb_i[34]
port 336 nsew signal output
rlabel metal2 s 199472 79600 199528 80000 6 tri_wbs_stb_i[35]
port 337 nsew signal output
rlabel metal2 s 197344 79600 197400 80000 6 tri_wbs_stb_i[36]
port 338 nsew signal output
rlabel metal2 s 195216 79600 195272 80000 6 tri_wbs_stb_i[37]
port 339 nsew signal output
rlabel metal2 s 193088 79600 193144 80000 6 tri_wbs_stb_i[38]
port 340 nsew signal output
rlabel metal2 s 190960 79600 191016 80000 6 tri_wbs_stb_i[39]
port 341 nsew signal output
rlabel metal2 s 267568 79600 267624 80000 6 tri_wbs_stb_i[3]
port 342 nsew signal output
rlabel metal2 s 188832 79600 188888 80000 6 tri_wbs_stb_i[40]
port 343 nsew signal output
rlabel metal2 s 186704 79600 186760 80000 6 tri_wbs_stb_i[41]
port 344 nsew signal output
rlabel metal2 s 184576 79600 184632 80000 6 tri_wbs_stb_i[42]
port 345 nsew signal output
rlabel metal2 s 182448 79600 182504 80000 6 tri_wbs_stb_i[43]
port 346 nsew signal output
rlabel metal2 s 180320 79600 180376 80000 6 tri_wbs_stb_i[44]
port 347 nsew signal output
rlabel metal2 s 178192 79600 178248 80000 6 tri_wbs_stb_i[45]
port 348 nsew signal output
rlabel metal2 s 176064 79600 176120 80000 6 tri_wbs_stb_i[46]
port 349 nsew signal output
rlabel metal2 s 173936 79600 173992 80000 6 tri_wbs_stb_i[47]
port 350 nsew signal output
rlabel metal2 s 171808 79600 171864 80000 6 tri_wbs_stb_i[48]
port 351 nsew signal output
rlabel metal2 s 169680 79600 169736 80000 6 tri_wbs_stb_i[49]
port 352 nsew signal output
rlabel metal2 s 265440 79600 265496 80000 6 tri_wbs_stb_i[4]
port 353 nsew signal output
rlabel metal2 s 167552 79600 167608 80000 6 tri_wbs_stb_i[50]
port 354 nsew signal output
rlabel metal2 s 165424 79600 165480 80000 6 tri_wbs_stb_i[51]
port 355 nsew signal output
rlabel metal2 s 163296 79600 163352 80000 6 tri_wbs_stb_i[52]
port 356 nsew signal output
rlabel metal2 s 161168 79600 161224 80000 6 tri_wbs_stb_i[53]
port 357 nsew signal output
rlabel metal2 s 159040 79600 159096 80000 6 tri_wbs_stb_i[54]
port 358 nsew signal output
rlabel metal2 s 156912 79600 156968 80000 6 tri_wbs_stb_i[55]
port 359 nsew signal output
rlabel metal2 s 154784 79600 154840 80000 6 tri_wbs_stb_i[56]
port 360 nsew signal output
rlabel metal2 s 152656 79600 152712 80000 6 tri_wbs_stb_i[57]
port 361 nsew signal output
rlabel metal2 s 150528 79600 150584 80000 6 tri_wbs_stb_i[58]
port 362 nsew signal output
rlabel metal2 s 148400 79600 148456 80000 6 tri_wbs_stb_i[59]
port 363 nsew signal output
rlabel metal2 s 263312 79600 263368 80000 6 tri_wbs_stb_i[5]
port 364 nsew signal output
rlabel metal2 s 146272 79600 146328 80000 6 tri_wbs_stb_i[60]
port 365 nsew signal output
rlabel metal2 s 144144 79600 144200 80000 6 tri_wbs_stb_i[61]
port 366 nsew signal output
rlabel metal2 s 142016 79600 142072 80000 6 tri_wbs_stb_i[62]
port 367 nsew signal output
rlabel metal2 s 139888 79600 139944 80000 6 tri_wbs_stb_i[63]
port 368 nsew signal output
rlabel metal2 s 261184 79600 261240 80000 6 tri_wbs_stb_i[6]
port 369 nsew signal output
rlabel metal2 s 259056 79600 259112 80000 6 tri_wbs_stb_i[7]
port 370 nsew signal output
rlabel metal2 s 256928 79600 256984 80000 6 tri_wbs_stb_i[8]
port 371 nsew signal output
rlabel metal2 s 254800 79600 254856 80000 6 tri_wbs_stb_i[9]
port 372 nsew signal output
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 78430 6 vdd
port 373 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 78430 6 vss
port 374 nsew ground bidirectional
rlabel metal2 s 3472 0 3528 400 6 wb_clk_i
port 375 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wb_rst_i
port 376 nsew signal input
rlabel metal2 s 4144 0 4200 400 6 wbs_ack_o
port 377 nsew signal output
rlabel metal2 s 5488 0 5544 400 6 wbs_adr_i[0]
port 378 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 wbs_adr_i[10]
port 379 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 wbs_adr_i[11]
port 380 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_adr_i[12]
port 381 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_adr_i[13]
port 382 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 wbs_adr_i[14]
port 383 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 wbs_adr_i[15]
port 384 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 wbs_adr_i[16]
port 385 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 wbs_adr_i[17]
port 386 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 wbs_adr_i[18]
port 387 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 wbs_adr_i[19]
port 388 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 wbs_adr_i[1]
port 389 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_adr_i[20]
port 390 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 wbs_adr_i[21]
port 391 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 wbs_adr_i[22]
port 392 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 wbs_adr_i[23]
port 393 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 wbs_adr_i[24]
port 394 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 wbs_adr_i[25]
port 395 nsew signal input
rlabel metal2 s 33040 0 33096 400 6 wbs_adr_i[26]
port 396 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 wbs_adr_i[27]
port 397 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 wbs_adr_i[28]
port 398 nsew signal input
rlabel metal2 s 36064 0 36120 400 6 wbs_adr_i[29]
port 399 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_adr_i[2]
port 400 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 wbs_adr_i[30]
port 401 nsew signal input
rlabel metal2 s 38080 0 38136 400 6 wbs_adr_i[31]
port 402 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_adr_i[3]
port 403 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_adr_i[4]
port 404 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_adr_i[5]
port 405 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_adr_i[6]
port 406 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 wbs_adr_i[7]
port 407 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_adr_i[8]
port 408 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_adr_i[9]
port 409 nsew signal input
rlabel metal2 s 4480 0 4536 400 6 wbs_cyc_i
port 410 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 wbs_dat_i[0]
port 411 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_dat_i[10]
port 412 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 wbs_dat_i[11]
port 413 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 wbs_dat_i[12]
port 414 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_dat_i[13]
port 415 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 wbs_dat_i[14]
port 416 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_i[15]
port 417 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 wbs_dat_i[16]
port 418 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_dat_i[17]
port 419 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 wbs_dat_i[18]
port 420 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 wbs_dat_i[19]
port 421 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 wbs_dat_i[1]
port 422 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 wbs_dat_i[20]
port 423 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_dat_i[21]
port 424 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 wbs_dat_i[22]
port 425 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 wbs_dat_i[23]
port 426 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 wbs_dat_i[24]
port 427 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 wbs_dat_i[25]
port 428 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 wbs_dat_i[26]
port 429 nsew signal input
rlabel metal2 s 34384 0 34440 400 6 wbs_dat_i[27]
port 430 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 wbs_dat_i[28]
port 431 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 wbs_dat_i[29]
port 432 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 wbs_dat_i[2]
port 433 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 wbs_dat_i[30]
port 434 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 wbs_dat_i[31]
port 435 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 wbs_dat_i[3]
port 436 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 wbs_dat_i[4]
port 437 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_dat_i[5]
port 438 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_dat_i[6]
port 439 nsew signal input
rlabel metal2 s 14224 0 14280 400 6 wbs_dat_i[7]
port 440 nsew signal input
rlabel metal2 s 15232 0 15288 400 6 wbs_dat_i[8]
port 441 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_i[9]
port 442 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 wbs_dat_o[0]
port 443 nsew signal output
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_o[10]
port 444 nsew signal output
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_o[11]
port 445 nsew signal output
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_o[12]
port 446 nsew signal output
rlabel metal2 s 20608 0 20664 400 6 wbs_dat_o[13]
port 447 nsew signal output
rlabel metal2 s 21616 0 21672 400 6 wbs_dat_o[14]
port 448 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 wbs_dat_o[15]
port 449 nsew signal output
rlabel metal2 s 23632 0 23688 400 6 wbs_dat_o[16]
port 450 nsew signal output
rlabel metal2 s 24640 0 24696 400 6 wbs_dat_o[17]
port 451 nsew signal output
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_o[18]
port 452 nsew signal output
rlabel metal2 s 26656 0 26712 400 6 wbs_dat_o[19]
port 453 nsew signal output
rlabel metal2 s 7504 0 7560 400 6 wbs_dat_o[1]
port 454 nsew signal output
rlabel metal2 s 27664 0 27720 400 6 wbs_dat_o[20]
port 455 nsew signal output
rlabel metal2 s 28672 0 28728 400 6 wbs_dat_o[21]
port 456 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 wbs_dat_o[22]
port 457 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 wbs_dat_o[23]
port 458 nsew signal output
rlabel metal2 s 31696 0 31752 400 6 wbs_dat_o[24]
port 459 nsew signal output
rlabel metal2 s 32704 0 32760 400 6 wbs_dat_o[25]
port 460 nsew signal output
rlabel metal2 s 33712 0 33768 400 6 wbs_dat_o[26]
port 461 nsew signal output
rlabel metal2 s 34720 0 34776 400 6 wbs_dat_o[27]
port 462 nsew signal output
rlabel metal2 s 35728 0 35784 400 6 wbs_dat_o[28]
port 463 nsew signal output
rlabel metal2 s 36736 0 36792 400 6 wbs_dat_o[29]
port 464 nsew signal output
rlabel metal2 s 8848 0 8904 400 6 wbs_dat_o[2]
port 465 nsew signal output
rlabel metal2 s 37744 0 37800 400 6 wbs_dat_o[30]
port 466 nsew signal output
rlabel metal2 s 38752 0 38808 400 6 wbs_dat_o[31]
port 467 nsew signal output
rlabel metal2 s 10192 0 10248 400 6 wbs_dat_o[3]
port 468 nsew signal output
rlabel metal2 s 11536 0 11592 400 6 wbs_dat_o[4]
port 469 nsew signal output
rlabel metal2 s 12544 0 12600 400 6 wbs_dat_o[5]
port 470 nsew signal output
rlabel metal2 s 13552 0 13608 400 6 wbs_dat_o[6]
port 471 nsew signal output
rlabel metal2 s 14560 0 14616 400 6 wbs_dat_o[7]
port 472 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 wbs_dat_o[8]
port 473 nsew signal output
rlabel metal2 s 16576 0 16632 400 6 wbs_dat_o[9]
port 474 nsew signal output
rlabel metal2 s 6496 0 6552 400 6 wbs_sel_i[0]
port 475 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_sel_i[1]
port 476 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 wbs_sel_i[2]
port 477 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 wbs_sel_i[3]
port 478 nsew signal input
rlabel metal2 s 4816 0 4872 400 6 wbs_stb_i
port 479 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 wbs_we_i
port 480 nsew signal input
rlabel metal3 s 0 67200 400 67256 6 x_end[0]
port 481 nsew signal input
rlabel metal3 s 0 56000 400 56056 6 x_end[100]
port 482 nsew signal input
rlabel metal3 s 0 55888 400 55944 6 x_end[101]
port 483 nsew signal input
rlabel metal3 s 0 55776 400 55832 6 x_end[102]
port 484 nsew signal input
rlabel metal3 s 0 55664 400 55720 6 x_end[103]
port 485 nsew signal input
rlabel metal3 s 0 55552 400 55608 6 x_end[104]
port 486 nsew signal input
rlabel metal3 s 0 55440 400 55496 6 x_end[105]
port 487 nsew signal input
rlabel metal3 s 0 55328 400 55384 6 x_end[106]
port 488 nsew signal input
rlabel metal3 s 0 55216 400 55272 6 x_end[107]
port 489 nsew signal input
rlabel metal3 s 0 55104 400 55160 6 x_end[108]
port 490 nsew signal input
rlabel metal3 s 0 54992 400 55048 6 x_end[109]
port 491 nsew signal input
rlabel metal3 s 0 66080 400 66136 6 x_end[10]
port 492 nsew signal input
rlabel metal3 s 0 54880 400 54936 6 x_end[110]
port 493 nsew signal input
rlabel metal3 s 0 54768 400 54824 6 x_end[111]
port 494 nsew signal input
rlabel metal3 s 0 54656 400 54712 6 x_end[112]
port 495 nsew signal input
rlabel metal3 s 0 54544 400 54600 6 x_end[113]
port 496 nsew signal input
rlabel metal3 s 0 54432 400 54488 6 x_end[114]
port 497 nsew signal input
rlabel metal3 s 0 54320 400 54376 6 x_end[115]
port 498 nsew signal input
rlabel metal3 s 0 54208 400 54264 6 x_end[116]
port 499 nsew signal input
rlabel metal3 s 0 54096 400 54152 6 x_end[117]
port 500 nsew signal input
rlabel metal3 s 0 53984 400 54040 6 x_end[118]
port 501 nsew signal input
rlabel metal3 s 0 53872 400 53928 6 x_end[119]
port 502 nsew signal input
rlabel metal3 s 0 65968 400 66024 6 x_end[11]
port 503 nsew signal input
rlabel metal3 s 0 53760 400 53816 6 x_end[120]
port 504 nsew signal input
rlabel metal3 s 0 53648 400 53704 6 x_end[121]
port 505 nsew signal input
rlabel metal3 s 0 53536 400 53592 6 x_end[122]
port 506 nsew signal input
rlabel metal3 s 0 53424 400 53480 6 x_end[123]
port 507 nsew signal input
rlabel metal3 s 0 53312 400 53368 6 x_end[124]
port 508 nsew signal input
rlabel metal3 s 0 53200 400 53256 6 x_end[125]
port 509 nsew signal input
rlabel metal3 s 0 53088 400 53144 6 x_end[126]
port 510 nsew signal input
rlabel metal3 s 0 52976 400 53032 6 x_end[127]
port 511 nsew signal input
rlabel metal3 s 0 52864 400 52920 6 x_end[128]
port 512 nsew signal input
rlabel metal3 s 0 52752 400 52808 6 x_end[129]
port 513 nsew signal input
rlabel metal3 s 0 65856 400 65912 6 x_end[12]
port 514 nsew signal input
rlabel metal3 s 0 52640 400 52696 6 x_end[130]
port 515 nsew signal input
rlabel metal3 s 0 52528 400 52584 6 x_end[131]
port 516 nsew signal input
rlabel metal3 s 0 52416 400 52472 6 x_end[132]
port 517 nsew signal input
rlabel metal3 s 0 52304 400 52360 6 x_end[133]
port 518 nsew signal input
rlabel metal3 s 0 52192 400 52248 6 x_end[134]
port 519 nsew signal input
rlabel metal3 s 0 52080 400 52136 6 x_end[135]
port 520 nsew signal input
rlabel metal3 s 0 51968 400 52024 6 x_end[136]
port 521 nsew signal input
rlabel metal3 s 0 51856 400 51912 6 x_end[137]
port 522 nsew signal input
rlabel metal3 s 0 51744 400 51800 6 x_end[138]
port 523 nsew signal input
rlabel metal3 s 0 51632 400 51688 6 x_end[139]
port 524 nsew signal input
rlabel metal3 s 0 65744 400 65800 6 x_end[13]
port 525 nsew signal input
rlabel metal3 s 0 51520 400 51576 6 x_end[140]
port 526 nsew signal input
rlabel metal3 s 0 51408 400 51464 6 x_end[141]
port 527 nsew signal input
rlabel metal3 s 0 51296 400 51352 6 x_end[142]
port 528 nsew signal input
rlabel metal3 s 0 51184 400 51240 6 x_end[143]
port 529 nsew signal input
rlabel metal3 s 0 51072 400 51128 6 x_end[144]
port 530 nsew signal input
rlabel metal3 s 0 50960 400 51016 6 x_end[145]
port 531 nsew signal input
rlabel metal3 s 0 50848 400 50904 6 x_end[146]
port 532 nsew signal input
rlabel metal3 s 0 50736 400 50792 6 x_end[147]
port 533 nsew signal input
rlabel metal3 s 0 50624 400 50680 6 x_end[148]
port 534 nsew signal input
rlabel metal3 s 0 50512 400 50568 6 x_end[149]
port 535 nsew signal input
rlabel metal3 s 0 65632 400 65688 6 x_end[14]
port 536 nsew signal input
rlabel metal3 s 0 50400 400 50456 6 x_end[150]
port 537 nsew signal input
rlabel metal3 s 0 50288 400 50344 6 x_end[151]
port 538 nsew signal input
rlabel metal3 s 0 50176 400 50232 6 x_end[152]
port 539 nsew signal input
rlabel metal3 s 0 50064 400 50120 6 x_end[153]
port 540 nsew signal input
rlabel metal3 s 0 49952 400 50008 6 x_end[154]
port 541 nsew signal input
rlabel metal3 s 0 49840 400 49896 6 x_end[155]
port 542 nsew signal input
rlabel metal3 s 0 49728 400 49784 6 x_end[156]
port 543 nsew signal input
rlabel metal3 s 0 49616 400 49672 6 x_end[157]
port 544 nsew signal input
rlabel metal3 s 0 49504 400 49560 6 x_end[158]
port 545 nsew signal input
rlabel metal3 s 0 49392 400 49448 6 x_end[159]
port 546 nsew signal input
rlabel metal3 s 0 65520 400 65576 6 x_end[15]
port 547 nsew signal input
rlabel metal3 s 0 49280 400 49336 6 x_end[160]
port 548 nsew signal input
rlabel metal3 s 0 49168 400 49224 6 x_end[161]
port 549 nsew signal input
rlabel metal3 s 0 49056 400 49112 6 x_end[162]
port 550 nsew signal input
rlabel metal3 s 0 48944 400 49000 6 x_end[163]
port 551 nsew signal input
rlabel metal3 s 0 48832 400 48888 6 x_end[164]
port 552 nsew signal input
rlabel metal3 s 0 48720 400 48776 6 x_end[165]
port 553 nsew signal input
rlabel metal3 s 0 48608 400 48664 6 x_end[166]
port 554 nsew signal input
rlabel metal3 s 0 48496 400 48552 6 x_end[167]
port 555 nsew signal input
rlabel metal3 s 0 48384 400 48440 6 x_end[168]
port 556 nsew signal input
rlabel metal3 s 0 48272 400 48328 6 x_end[169]
port 557 nsew signal input
rlabel metal3 s 0 65408 400 65464 6 x_end[16]
port 558 nsew signal input
rlabel metal3 s 0 48160 400 48216 6 x_end[170]
port 559 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 x_end[171]
port 560 nsew signal input
rlabel metal3 s 0 47936 400 47992 6 x_end[172]
port 561 nsew signal input
rlabel metal3 s 0 47824 400 47880 6 x_end[173]
port 562 nsew signal input
rlabel metal3 s 0 47712 400 47768 6 x_end[174]
port 563 nsew signal input
rlabel metal3 s 0 47600 400 47656 6 x_end[175]
port 564 nsew signal input
rlabel metal3 s 0 47488 400 47544 6 x_end[176]
port 565 nsew signal input
rlabel metal3 s 0 47376 400 47432 6 x_end[177]
port 566 nsew signal input
rlabel metal3 s 0 47264 400 47320 6 x_end[178]
port 567 nsew signal input
rlabel metal3 s 0 47152 400 47208 6 x_end[179]
port 568 nsew signal input
rlabel metal3 s 0 65296 400 65352 6 x_end[17]
port 569 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 x_end[180]
port 570 nsew signal input
rlabel metal3 s 0 46928 400 46984 6 x_end[181]
port 571 nsew signal input
rlabel metal3 s 0 46816 400 46872 6 x_end[182]
port 572 nsew signal input
rlabel metal3 s 0 46704 400 46760 6 x_end[183]
port 573 nsew signal input
rlabel metal3 s 0 46592 400 46648 6 x_end[184]
port 574 nsew signal input
rlabel metal3 s 0 46480 400 46536 6 x_end[185]
port 575 nsew signal input
rlabel metal3 s 0 46368 400 46424 6 x_end[186]
port 576 nsew signal input
rlabel metal3 s 0 46256 400 46312 6 x_end[187]
port 577 nsew signal input
rlabel metal3 s 0 46144 400 46200 6 x_end[188]
port 578 nsew signal input
rlabel metal3 s 0 46032 400 46088 6 x_end[189]
port 579 nsew signal input
rlabel metal3 s 0 65184 400 65240 6 x_end[18]
port 580 nsew signal input
rlabel metal3 s 0 45920 400 45976 6 x_end[190]
port 581 nsew signal input
rlabel metal3 s 0 45808 400 45864 6 x_end[191]
port 582 nsew signal input
rlabel metal3 s 0 45696 400 45752 6 x_end[192]
port 583 nsew signal input
rlabel metal3 s 0 45584 400 45640 6 x_end[193]
port 584 nsew signal input
rlabel metal3 s 0 45472 400 45528 6 x_end[194]
port 585 nsew signal input
rlabel metal3 s 0 45360 400 45416 6 x_end[195]
port 586 nsew signal input
rlabel metal3 s 0 45248 400 45304 6 x_end[196]
port 587 nsew signal input
rlabel metal3 s 0 45136 400 45192 6 x_end[197]
port 588 nsew signal input
rlabel metal3 s 0 45024 400 45080 6 x_end[198]
port 589 nsew signal input
rlabel metal3 s 0 44912 400 44968 6 x_end[199]
port 590 nsew signal input
rlabel metal3 s 0 65072 400 65128 6 x_end[19]
port 591 nsew signal input
rlabel metal3 s 0 67088 400 67144 6 x_end[1]
port 592 nsew signal input
rlabel metal3 s 0 44800 400 44856 6 x_end[200]
port 593 nsew signal input
rlabel metal3 s 0 44688 400 44744 6 x_end[201]
port 594 nsew signal input
rlabel metal3 s 0 44576 400 44632 6 x_end[202]
port 595 nsew signal input
rlabel metal3 s 0 44464 400 44520 6 x_end[203]
port 596 nsew signal input
rlabel metal3 s 0 44352 400 44408 6 x_end[204]
port 597 nsew signal input
rlabel metal3 s 0 44240 400 44296 6 x_end[205]
port 598 nsew signal input
rlabel metal3 s 0 44128 400 44184 6 x_end[206]
port 599 nsew signal input
rlabel metal3 s 0 44016 400 44072 6 x_end[207]
port 600 nsew signal input
rlabel metal3 s 0 43904 400 43960 6 x_end[208]
port 601 nsew signal input
rlabel metal3 s 0 43792 400 43848 6 x_end[209]
port 602 nsew signal input
rlabel metal3 s 0 64960 400 65016 6 x_end[20]
port 603 nsew signal input
rlabel metal3 s 0 43680 400 43736 6 x_end[210]
port 604 nsew signal input
rlabel metal3 s 0 43568 400 43624 6 x_end[211]
port 605 nsew signal input
rlabel metal3 s 0 43456 400 43512 6 x_end[212]
port 606 nsew signal input
rlabel metal3 s 0 43344 400 43400 6 x_end[213]
port 607 nsew signal input
rlabel metal3 s 0 43232 400 43288 6 x_end[214]
port 608 nsew signal input
rlabel metal3 s 0 43120 400 43176 6 x_end[215]
port 609 nsew signal input
rlabel metal3 s 0 43008 400 43064 6 x_end[216]
port 610 nsew signal input
rlabel metal3 s 0 42896 400 42952 6 x_end[217]
port 611 nsew signal input
rlabel metal3 s 0 42784 400 42840 6 x_end[218]
port 612 nsew signal input
rlabel metal3 s 0 42672 400 42728 6 x_end[219]
port 613 nsew signal input
rlabel metal3 s 0 64848 400 64904 6 x_end[21]
port 614 nsew signal input
rlabel metal3 s 0 42560 400 42616 6 x_end[220]
port 615 nsew signal input
rlabel metal3 s 0 42448 400 42504 6 x_end[221]
port 616 nsew signal input
rlabel metal3 s 0 42336 400 42392 6 x_end[222]
port 617 nsew signal input
rlabel metal3 s 0 42224 400 42280 6 x_end[223]
port 618 nsew signal input
rlabel metal3 s 0 42112 400 42168 6 x_end[224]
port 619 nsew signal input
rlabel metal3 s 0 42000 400 42056 6 x_end[225]
port 620 nsew signal input
rlabel metal3 s 0 41888 400 41944 6 x_end[226]
port 621 nsew signal input
rlabel metal3 s 0 41776 400 41832 6 x_end[227]
port 622 nsew signal input
rlabel metal3 s 0 41664 400 41720 6 x_end[228]
port 623 nsew signal input
rlabel metal3 s 0 41552 400 41608 6 x_end[229]
port 624 nsew signal input
rlabel metal3 s 0 64736 400 64792 6 x_end[22]
port 625 nsew signal input
rlabel metal3 s 0 41440 400 41496 6 x_end[230]
port 626 nsew signal input
rlabel metal3 s 0 41328 400 41384 6 x_end[231]
port 627 nsew signal input
rlabel metal3 s 0 41216 400 41272 6 x_end[232]
port 628 nsew signal input
rlabel metal3 s 0 41104 400 41160 6 x_end[233]
port 629 nsew signal input
rlabel metal3 s 0 40992 400 41048 6 x_end[234]
port 630 nsew signal input
rlabel metal3 s 0 40880 400 40936 6 x_end[235]
port 631 nsew signal input
rlabel metal3 s 0 40768 400 40824 6 x_end[236]
port 632 nsew signal input
rlabel metal3 s 0 40656 400 40712 6 x_end[237]
port 633 nsew signal input
rlabel metal3 s 0 40544 400 40600 6 x_end[238]
port 634 nsew signal input
rlabel metal3 s 0 40432 400 40488 6 x_end[239]
port 635 nsew signal input
rlabel metal3 s 0 64624 400 64680 6 x_end[23]
port 636 nsew signal input
rlabel metal3 s 0 40320 400 40376 6 x_end[240]
port 637 nsew signal input
rlabel metal3 s 0 40208 400 40264 6 x_end[241]
port 638 nsew signal input
rlabel metal3 s 0 40096 400 40152 6 x_end[242]
port 639 nsew signal input
rlabel metal3 s 0 39984 400 40040 6 x_end[243]
port 640 nsew signal input
rlabel metal3 s 0 39872 400 39928 6 x_end[244]
port 641 nsew signal input
rlabel metal3 s 0 39760 400 39816 6 x_end[245]
port 642 nsew signal input
rlabel metal3 s 0 39648 400 39704 6 x_end[246]
port 643 nsew signal input
rlabel metal3 s 0 39536 400 39592 6 x_end[247]
port 644 nsew signal input
rlabel metal3 s 0 39424 400 39480 6 x_end[248]
port 645 nsew signal input
rlabel metal3 s 0 39312 400 39368 6 x_end[249]
port 646 nsew signal input
rlabel metal3 s 0 64512 400 64568 6 x_end[24]
port 647 nsew signal input
rlabel metal3 s 0 39200 400 39256 6 x_end[250]
port 648 nsew signal input
rlabel metal3 s 0 39088 400 39144 6 x_end[251]
port 649 nsew signal input
rlabel metal3 s 0 38976 400 39032 6 x_end[252]
port 650 nsew signal input
rlabel metal3 s 0 38864 400 38920 6 x_end[253]
port 651 nsew signal input
rlabel metal3 s 0 38752 400 38808 6 x_end[254]
port 652 nsew signal input
rlabel metal3 s 0 38640 400 38696 6 x_end[255]
port 653 nsew signal input
rlabel metal3 s 0 38528 400 38584 6 x_end[256]
port 654 nsew signal input
rlabel metal3 s 0 38416 400 38472 6 x_end[257]
port 655 nsew signal input
rlabel metal3 s 0 38304 400 38360 6 x_end[258]
port 656 nsew signal input
rlabel metal3 s 0 38192 400 38248 6 x_end[259]
port 657 nsew signal input
rlabel metal3 s 0 64400 400 64456 6 x_end[25]
port 658 nsew signal input
rlabel metal3 s 0 38080 400 38136 6 x_end[260]
port 659 nsew signal input
rlabel metal3 s 0 37968 400 38024 6 x_end[261]
port 660 nsew signal input
rlabel metal3 s 0 37856 400 37912 6 x_end[262]
port 661 nsew signal input
rlabel metal3 s 0 37744 400 37800 6 x_end[263]
port 662 nsew signal input
rlabel metal3 s 0 37632 400 37688 6 x_end[264]
port 663 nsew signal input
rlabel metal3 s 0 37520 400 37576 6 x_end[265]
port 664 nsew signal input
rlabel metal3 s 0 37408 400 37464 6 x_end[266]
port 665 nsew signal input
rlabel metal3 s 0 37296 400 37352 6 x_end[267]
port 666 nsew signal input
rlabel metal3 s 0 37184 400 37240 6 x_end[268]
port 667 nsew signal input
rlabel metal3 s 0 37072 400 37128 6 x_end[269]
port 668 nsew signal input
rlabel metal3 s 0 64288 400 64344 6 x_end[26]
port 669 nsew signal input
rlabel metal3 s 0 36960 400 37016 6 x_end[270]
port 670 nsew signal input
rlabel metal3 s 0 36848 400 36904 6 x_end[271]
port 671 nsew signal input
rlabel metal3 s 0 36736 400 36792 6 x_end[272]
port 672 nsew signal input
rlabel metal3 s 0 36624 400 36680 6 x_end[273]
port 673 nsew signal input
rlabel metal3 s 0 36512 400 36568 6 x_end[274]
port 674 nsew signal input
rlabel metal3 s 0 36400 400 36456 6 x_end[275]
port 675 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 x_end[276]
port 676 nsew signal input
rlabel metal3 s 0 36176 400 36232 6 x_end[277]
port 677 nsew signal input
rlabel metal3 s 0 36064 400 36120 6 x_end[278]
port 678 nsew signal input
rlabel metal3 s 0 35952 400 36008 6 x_end[279]
port 679 nsew signal input
rlabel metal3 s 0 64176 400 64232 6 x_end[27]
port 680 nsew signal input
rlabel metal3 s 0 35840 400 35896 6 x_end[280]
port 681 nsew signal input
rlabel metal3 s 0 35728 400 35784 6 x_end[281]
port 682 nsew signal input
rlabel metal3 s 0 35616 400 35672 6 x_end[282]
port 683 nsew signal input
rlabel metal3 s 0 35504 400 35560 6 x_end[283]
port 684 nsew signal input
rlabel metal3 s 0 35392 400 35448 6 x_end[284]
port 685 nsew signal input
rlabel metal3 s 0 35280 400 35336 6 x_end[285]
port 686 nsew signal input
rlabel metal3 s 0 35168 400 35224 6 x_end[286]
port 687 nsew signal input
rlabel metal3 s 0 35056 400 35112 6 x_end[287]
port 688 nsew signal input
rlabel metal3 s 0 34944 400 35000 6 x_end[288]
port 689 nsew signal input
rlabel metal3 s 0 34832 400 34888 6 x_end[289]
port 690 nsew signal input
rlabel metal3 s 0 64064 400 64120 6 x_end[28]
port 691 nsew signal input
rlabel metal3 s 0 34720 400 34776 6 x_end[290]
port 692 nsew signal input
rlabel metal3 s 0 34608 400 34664 6 x_end[291]
port 693 nsew signal input
rlabel metal3 s 0 34496 400 34552 6 x_end[292]
port 694 nsew signal input
rlabel metal3 s 0 34384 400 34440 6 x_end[293]
port 695 nsew signal input
rlabel metal3 s 0 34272 400 34328 6 x_end[294]
port 696 nsew signal input
rlabel metal3 s 0 34160 400 34216 6 x_end[295]
port 697 nsew signal input
rlabel metal3 s 0 34048 400 34104 6 x_end[296]
port 698 nsew signal input
rlabel metal3 s 0 33936 400 33992 6 x_end[297]
port 699 nsew signal input
rlabel metal3 s 0 33824 400 33880 6 x_end[298]
port 700 nsew signal input
rlabel metal3 s 0 33712 400 33768 6 x_end[299]
port 701 nsew signal input
rlabel metal3 s 0 63952 400 64008 6 x_end[29]
port 702 nsew signal input
rlabel metal3 s 0 66976 400 67032 6 x_end[2]
port 703 nsew signal input
rlabel metal3 s 0 33600 400 33656 6 x_end[300]
port 704 nsew signal input
rlabel metal3 s 0 33488 400 33544 6 x_end[301]
port 705 nsew signal input
rlabel metal3 s 0 33376 400 33432 6 x_end[302]
port 706 nsew signal input
rlabel metal3 s 0 33264 400 33320 6 x_end[303]
port 707 nsew signal input
rlabel metal3 s 0 33152 400 33208 6 x_end[304]
port 708 nsew signal input
rlabel metal3 s 0 33040 400 33096 6 x_end[305]
port 709 nsew signal input
rlabel metal3 s 0 32928 400 32984 6 x_end[306]
port 710 nsew signal input
rlabel metal3 s 0 32816 400 32872 6 x_end[307]
port 711 nsew signal input
rlabel metal3 s 0 32704 400 32760 6 x_end[308]
port 712 nsew signal input
rlabel metal3 s 0 32592 400 32648 6 x_end[309]
port 713 nsew signal input
rlabel metal3 s 0 63840 400 63896 6 x_end[30]
port 714 nsew signal input
rlabel metal3 s 0 32480 400 32536 6 x_end[310]
port 715 nsew signal input
rlabel metal3 s 0 32368 400 32424 6 x_end[311]
port 716 nsew signal input
rlabel metal3 s 0 32256 400 32312 6 x_end[312]
port 717 nsew signal input
rlabel metal3 s 0 32144 400 32200 6 x_end[313]
port 718 nsew signal input
rlabel metal3 s 0 32032 400 32088 6 x_end[314]
port 719 nsew signal input
rlabel metal3 s 0 31920 400 31976 6 x_end[315]
port 720 nsew signal input
rlabel metal3 s 0 31808 400 31864 6 x_end[316]
port 721 nsew signal input
rlabel metal3 s 0 31696 400 31752 6 x_end[317]
port 722 nsew signal input
rlabel metal3 s 0 31584 400 31640 6 x_end[318]
port 723 nsew signal input
rlabel metal3 s 0 31472 400 31528 6 x_end[319]
port 724 nsew signal input
rlabel metal3 s 0 63728 400 63784 6 x_end[31]
port 725 nsew signal input
rlabel metal3 s 0 31360 400 31416 6 x_end[320]
port 726 nsew signal input
rlabel metal3 s 0 31248 400 31304 6 x_end[321]
port 727 nsew signal input
rlabel metal3 s 0 31136 400 31192 6 x_end[322]
port 728 nsew signal input
rlabel metal3 s 0 31024 400 31080 6 x_end[323]
port 729 nsew signal input
rlabel metal3 s 0 30912 400 30968 6 x_end[324]
port 730 nsew signal input
rlabel metal3 s 0 30800 400 30856 6 x_end[325]
port 731 nsew signal input
rlabel metal3 s 0 30688 400 30744 6 x_end[326]
port 732 nsew signal input
rlabel metal3 s 0 30576 400 30632 6 x_end[327]
port 733 nsew signal input
rlabel metal3 s 0 30464 400 30520 6 x_end[328]
port 734 nsew signal input
rlabel metal3 s 0 30352 400 30408 6 x_end[329]
port 735 nsew signal input
rlabel metal3 s 0 63616 400 63672 6 x_end[32]
port 736 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 x_end[330]
port 737 nsew signal input
rlabel metal3 s 0 30128 400 30184 6 x_end[331]
port 738 nsew signal input
rlabel metal3 s 0 30016 400 30072 6 x_end[332]
port 739 nsew signal input
rlabel metal3 s 0 29904 400 29960 6 x_end[333]
port 740 nsew signal input
rlabel metal3 s 0 29792 400 29848 6 x_end[334]
port 741 nsew signal input
rlabel metal3 s 0 29680 400 29736 6 x_end[335]
port 742 nsew signal input
rlabel metal3 s 0 29568 400 29624 6 x_end[336]
port 743 nsew signal input
rlabel metal3 s 0 29456 400 29512 6 x_end[337]
port 744 nsew signal input
rlabel metal3 s 0 29344 400 29400 6 x_end[338]
port 745 nsew signal input
rlabel metal3 s 0 29232 400 29288 6 x_end[339]
port 746 nsew signal input
rlabel metal3 s 0 63504 400 63560 6 x_end[33]
port 747 nsew signal input
rlabel metal3 s 0 29120 400 29176 6 x_end[340]
port 748 nsew signal input
rlabel metal3 s 0 29008 400 29064 6 x_end[341]
port 749 nsew signal input
rlabel metal3 s 0 28896 400 28952 6 x_end[342]
port 750 nsew signal input
rlabel metal3 s 0 28784 400 28840 6 x_end[343]
port 751 nsew signal input
rlabel metal3 s 0 28672 400 28728 6 x_end[344]
port 752 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 x_end[345]
port 753 nsew signal input
rlabel metal3 s 0 28448 400 28504 6 x_end[346]
port 754 nsew signal input
rlabel metal3 s 0 28336 400 28392 6 x_end[347]
port 755 nsew signal input
rlabel metal3 s 0 28224 400 28280 6 x_end[348]
port 756 nsew signal input
rlabel metal3 s 0 28112 400 28168 6 x_end[349]
port 757 nsew signal input
rlabel metal3 s 0 63392 400 63448 6 x_end[34]
port 758 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 x_end[350]
port 759 nsew signal input
rlabel metal3 s 0 27888 400 27944 6 x_end[351]
port 760 nsew signal input
rlabel metal3 s 0 27776 400 27832 6 x_end[352]
port 761 nsew signal input
rlabel metal3 s 0 27664 400 27720 6 x_end[353]
port 762 nsew signal input
rlabel metal3 s 0 27552 400 27608 6 x_end[354]
port 763 nsew signal input
rlabel metal3 s 0 27440 400 27496 6 x_end[355]
port 764 nsew signal input
rlabel metal3 s 0 27328 400 27384 6 x_end[356]
port 765 nsew signal input
rlabel metal3 s 0 27216 400 27272 6 x_end[357]
port 766 nsew signal input
rlabel metal3 s 0 27104 400 27160 6 x_end[358]
port 767 nsew signal input
rlabel metal3 s 0 26992 400 27048 6 x_end[359]
port 768 nsew signal input
rlabel metal3 s 0 63280 400 63336 6 x_end[35]
port 769 nsew signal input
rlabel metal3 s 0 26880 400 26936 6 x_end[360]
port 770 nsew signal input
rlabel metal3 s 0 26768 400 26824 6 x_end[361]
port 771 nsew signal input
rlabel metal3 s 0 26656 400 26712 6 x_end[362]
port 772 nsew signal input
rlabel metal3 s 0 26544 400 26600 6 x_end[363]
port 773 nsew signal input
rlabel metal3 s 0 26432 400 26488 6 x_end[364]
port 774 nsew signal input
rlabel metal3 s 0 26320 400 26376 6 x_end[365]
port 775 nsew signal input
rlabel metal3 s 0 26208 400 26264 6 x_end[366]
port 776 nsew signal input
rlabel metal3 s 0 26096 400 26152 6 x_end[367]
port 777 nsew signal input
rlabel metal3 s 0 25984 400 26040 6 x_end[368]
port 778 nsew signal input
rlabel metal3 s 0 25872 400 25928 6 x_end[369]
port 779 nsew signal input
rlabel metal3 s 0 63168 400 63224 6 x_end[36]
port 780 nsew signal input
rlabel metal3 s 0 25760 400 25816 6 x_end[370]
port 781 nsew signal input
rlabel metal3 s 0 25648 400 25704 6 x_end[371]
port 782 nsew signal input
rlabel metal3 s 0 25536 400 25592 6 x_end[372]
port 783 nsew signal input
rlabel metal3 s 0 25424 400 25480 6 x_end[373]
port 784 nsew signal input
rlabel metal3 s 0 25312 400 25368 6 x_end[374]
port 785 nsew signal input
rlabel metal3 s 0 25200 400 25256 6 x_end[375]
port 786 nsew signal input
rlabel metal3 s 0 25088 400 25144 6 x_end[376]
port 787 nsew signal input
rlabel metal3 s 0 24976 400 25032 6 x_end[377]
port 788 nsew signal input
rlabel metal3 s 0 24864 400 24920 6 x_end[378]
port 789 nsew signal input
rlabel metal3 s 0 24752 400 24808 6 x_end[379]
port 790 nsew signal input
rlabel metal3 s 0 63056 400 63112 6 x_end[37]
port 791 nsew signal input
rlabel metal3 s 0 24640 400 24696 6 x_end[380]
port 792 nsew signal input
rlabel metal3 s 0 24528 400 24584 6 x_end[381]
port 793 nsew signal input
rlabel metal3 s 0 24416 400 24472 6 x_end[382]
port 794 nsew signal input
rlabel metal3 s 0 24304 400 24360 6 x_end[383]
port 795 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 x_end[384]
port 796 nsew signal input
rlabel metal3 s 0 24080 400 24136 6 x_end[385]
port 797 nsew signal input
rlabel metal3 s 0 23968 400 24024 6 x_end[386]
port 798 nsew signal input
rlabel metal3 s 0 23856 400 23912 6 x_end[387]
port 799 nsew signal input
rlabel metal3 s 0 23744 400 23800 6 x_end[388]
port 800 nsew signal input
rlabel metal3 s 0 23632 400 23688 6 x_end[389]
port 801 nsew signal input
rlabel metal3 s 0 62944 400 63000 6 x_end[38]
port 802 nsew signal input
rlabel metal3 s 0 23520 400 23576 6 x_end[390]
port 803 nsew signal input
rlabel metal3 s 0 23408 400 23464 6 x_end[391]
port 804 nsew signal input
rlabel metal3 s 0 23296 400 23352 6 x_end[392]
port 805 nsew signal input
rlabel metal3 s 0 23184 400 23240 6 x_end[393]
port 806 nsew signal input
rlabel metal3 s 0 23072 400 23128 6 x_end[394]
port 807 nsew signal input
rlabel metal3 s 0 22960 400 23016 6 x_end[395]
port 808 nsew signal input
rlabel metal3 s 0 22848 400 22904 6 x_end[396]
port 809 nsew signal input
rlabel metal3 s 0 22736 400 22792 6 x_end[397]
port 810 nsew signal input
rlabel metal3 s 0 22624 400 22680 6 x_end[398]
port 811 nsew signal input
rlabel metal3 s 0 22512 400 22568 6 x_end[399]
port 812 nsew signal input
rlabel metal3 s 0 62832 400 62888 6 x_end[39]
port 813 nsew signal input
rlabel metal3 s 0 66864 400 66920 6 x_end[3]
port 814 nsew signal input
rlabel metal3 s 0 22400 400 22456 6 x_end[400]
port 815 nsew signal input
rlabel metal3 s 0 22288 400 22344 6 x_end[401]
port 816 nsew signal input
rlabel metal3 s 0 22176 400 22232 6 x_end[402]
port 817 nsew signal input
rlabel metal3 s 0 22064 400 22120 6 x_end[403]
port 818 nsew signal input
rlabel metal3 s 0 21952 400 22008 6 x_end[404]
port 819 nsew signal input
rlabel metal3 s 0 21840 400 21896 6 x_end[405]
port 820 nsew signal input
rlabel metal3 s 0 21728 400 21784 6 x_end[406]
port 821 nsew signal input
rlabel metal3 s 0 21616 400 21672 6 x_end[407]
port 822 nsew signal input
rlabel metal3 s 0 21504 400 21560 6 x_end[408]
port 823 nsew signal input
rlabel metal3 s 0 21392 400 21448 6 x_end[409]
port 824 nsew signal input
rlabel metal3 s 0 62720 400 62776 6 x_end[40]
port 825 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 x_end[410]
port 826 nsew signal input
rlabel metal3 s 0 21168 400 21224 6 x_end[411]
port 827 nsew signal input
rlabel metal3 s 0 21056 400 21112 6 x_end[412]
port 828 nsew signal input
rlabel metal3 s 0 20944 400 21000 6 x_end[413]
port 829 nsew signal input
rlabel metal3 s 0 20832 400 20888 6 x_end[414]
port 830 nsew signal input
rlabel metal3 s 0 20720 400 20776 6 x_end[415]
port 831 nsew signal input
rlabel metal3 s 0 20608 400 20664 6 x_end[416]
port 832 nsew signal input
rlabel metal3 s 0 20496 400 20552 6 x_end[417]
port 833 nsew signal input
rlabel metal3 s 0 20384 400 20440 6 x_end[418]
port 834 nsew signal input
rlabel metal3 s 0 20272 400 20328 6 x_end[419]
port 835 nsew signal input
rlabel metal3 s 0 62608 400 62664 6 x_end[41]
port 836 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 x_end[420]
port 837 nsew signal input
rlabel metal3 s 0 20048 400 20104 6 x_end[421]
port 838 nsew signal input
rlabel metal3 s 0 19936 400 19992 6 x_end[422]
port 839 nsew signal input
rlabel metal3 s 0 19824 400 19880 6 x_end[423]
port 840 nsew signal input
rlabel metal3 s 0 19712 400 19768 6 x_end[424]
port 841 nsew signal input
rlabel metal3 s 0 19600 400 19656 6 x_end[425]
port 842 nsew signal input
rlabel metal3 s 0 19488 400 19544 6 x_end[426]
port 843 nsew signal input
rlabel metal3 s 0 19376 400 19432 6 x_end[427]
port 844 nsew signal input
rlabel metal3 s 0 19264 400 19320 6 x_end[428]
port 845 nsew signal input
rlabel metal3 s 0 19152 400 19208 6 x_end[429]
port 846 nsew signal input
rlabel metal3 s 0 62496 400 62552 6 x_end[42]
port 847 nsew signal input
rlabel metal3 s 0 19040 400 19096 6 x_end[430]
port 848 nsew signal input
rlabel metal3 s 0 18928 400 18984 6 x_end[431]
port 849 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 x_end[432]
port 850 nsew signal input
rlabel metal3 s 0 18704 400 18760 6 x_end[433]
port 851 nsew signal input
rlabel metal3 s 0 18592 400 18648 6 x_end[434]
port 852 nsew signal input
rlabel metal3 s 0 18480 400 18536 6 x_end[435]
port 853 nsew signal input
rlabel metal3 s 0 18368 400 18424 6 x_end[436]
port 854 nsew signal input
rlabel metal3 s 0 18256 400 18312 6 x_end[437]
port 855 nsew signal input
rlabel metal3 s 0 18144 400 18200 6 x_end[438]
port 856 nsew signal input
rlabel metal3 s 0 18032 400 18088 6 x_end[439]
port 857 nsew signal input
rlabel metal3 s 0 62384 400 62440 6 x_end[43]
port 858 nsew signal input
rlabel metal3 s 0 17920 400 17976 6 x_end[440]
port 859 nsew signal input
rlabel metal3 s 0 17808 400 17864 6 x_end[441]
port 860 nsew signal input
rlabel metal3 s 0 17696 400 17752 6 x_end[442]
port 861 nsew signal input
rlabel metal3 s 0 17584 400 17640 6 x_end[443]
port 862 nsew signal input
rlabel metal3 s 0 17472 400 17528 6 x_end[444]
port 863 nsew signal input
rlabel metal3 s 0 17360 400 17416 6 x_end[445]
port 864 nsew signal input
rlabel metal3 s 0 17248 400 17304 6 x_end[446]
port 865 nsew signal input
rlabel metal3 s 0 17136 400 17192 6 x_end[447]
port 866 nsew signal input
rlabel metal3 s 0 17024 400 17080 6 x_end[448]
port 867 nsew signal input
rlabel metal3 s 0 16912 400 16968 6 x_end[449]
port 868 nsew signal input
rlabel metal3 s 0 62272 400 62328 6 x_end[44]
port 869 nsew signal input
rlabel metal3 s 0 16800 400 16856 6 x_end[450]
port 870 nsew signal input
rlabel metal3 s 0 16688 400 16744 6 x_end[451]
port 871 nsew signal input
rlabel metal3 s 0 16576 400 16632 6 x_end[452]
port 872 nsew signal input
rlabel metal3 s 0 16464 400 16520 6 x_end[453]
port 873 nsew signal input
rlabel metal3 s 0 16352 400 16408 6 x_end[454]
port 874 nsew signal input
rlabel metal3 s 0 16240 400 16296 6 x_end[455]
port 875 nsew signal input
rlabel metal3 s 0 16128 400 16184 6 x_end[456]
port 876 nsew signal input
rlabel metal3 s 0 16016 400 16072 6 x_end[457]
port 877 nsew signal input
rlabel metal3 s 0 15904 400 15960 6 x_end[458]
port 878 nsew signal input
rlabel metal3 s 0 15792 400 15848 6 x_end[459]
port 879 nsew signal input
rlabel metal3 s 0 62160 400 62216 6 x_end[45]
port 880 nsew signal input
rlabel metal3 s 0 15680 400 15736 6 x_end[460]
port 881 nsew signal input
rlabel metal3 s 0 15568 400 15624 6 x_end[461]
port 882 nsew signal input
rlabel metal3 s 0 15456 400 15512 6 x_end[462]
port 883 nsew signal input
rlabel metal3 s 0 15344 400 15400 6 x_end[463]
port 884 nsew signal input
rlabel metal3 s 0 15232 400 15288 6 x_end[464]
port 885 nsew signal input
rlabel metal3 s 0 15120 400 15176 6 x_end[465]
port 886 nsew signal input
rlabel metal3 s 0 15008 400 15064 6 x_end[466]
port 887 nsew signal input
rlabel metal3 s 0 14896 400 14952 6 x_end[467]
port 888 nsew signal input
rlabel metal3 s 0 14784 400 14840 6 x_end[468]
port 889 nsew signal input
rlabel metal3 s 0 14672 400 14728 6 x_end[469]
port 890 nsew signal input
rlabel metal3 s 0 62048 400 62104 6 x_end[46]
port 891 nsew signal input
rlabel metal3 s 0 14560 400 14616 6 x_end[470]
port 892 nsew signal input
rlabel metal3 s 0 14448 400 14504 6 x_end[471]
port 893 nsew signal input
rlabel metal3 s 0 14336 400 14392 6 x_end[472]
port 894 nsew signal input
rlabel metal3 s 0 14224 400 14280 6 x_end[473]
port 895 nsew signal input
rlabel metal3 s 0 14112 400 14168 6 x_end[474]
port 896 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 x_end[475]
port 897 nsew signal input
rlabel metal3 s 0 13888 400 13944 6 x_end[476]
port 898 nsew signal input
rlabel metal3 s 0 13776 400 13832 6 x_end[477]
port 899 nsew signal input
rlabel metal3 s 0 13664 400 13720 6 x_end[478]
port 900 nsew signal input
rlabel metal3 s 0 13552 400 13608 6 x_end[479]
port 901 nsew signal input
rlabel metal3 s 0 61936 400 61992 6 x_end[47]
port 902 nsew signal input
rlabel metal3 s 0 13440 400 13496 6 x_end[480]
port 903 nsew signal input
rlabel metal3 s 0 13328 400 13384 6 x_end[481]
port 904 nsew signal input
rlabel metal3 s 0 13216 400 13272 6 x_end[482]
port 905 nsew signal input
rlabel metal3 s 0 13104 400 13160 6 x_end[483]
port 906 nsew signal input
rlabel metal3 s 0 12992 400 13048 6 x_end[484]
port 907 nsew signal input
rlabel metal3 s 0 12880 400 12936 6 x_end[485]
port 908 nsew signal input
rlabel metal3 s 0 12768 400 12824 6 x_end[486]
port 909 nsew signal input
rlabel metal3 s 0 12656 400 12712 6 x_end[487]
port 910 nsew signal input
rlabel metal3 s 0 12544 400 12600 6 x_end[488]
port 911 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 x_end[489]
port 912 nsew signal input
rlabel metal3 s 0 61824 400 61880 6 x_end[48]
port 913 nsew signal input
rlabel metal3 s 0 12320 400 12376 6 x_end[490]
port 914 nsew signal input
rlabel metal3 s 0 12208 400 12264 6 x_end[491]
port 915 nsew signal input
rlabel metal3 s 0 12096 400 12152 6 x_end[492]
port 916 nsew signal input
rlabel metal3 s 0 11984 400 12040 6 x_end[493]
port 917 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 x_end[494]
port 918 nsew signal input
rlabel metal3 s 0 11760 400 11816 6 x_end[495]
port 919 nsew signal input
rlabel metal3 s 0 11648 400 11704 6 x_end[496]
port 920 nsew signal input
rlabel metal3 s 0 11536 400 11592 6 x_end[497]
port 921 nsew signal input
rlabel metal3 s 0 11424 400 11480 6 x_end[498]
port 922 nsew signal input
rlabel metal3 s 0 11312 400 11368 6 x_end[499]
port 923 nsew signal input
rlabel metal3 s 0 61712 400 61768 6 x_end[49]
port 924 nsew signal input
rlabel metal3 s 0 66752 400 66808 6 x_end[4]
port 925 nsew signal input
rlabel metal3 s 0 11200 400 11256 6 x_end[500]
port 926 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 x_end[501]
port 927 nsew signal input
rlabel metal3 s 0 10976 400 11032 6 x_end[502]
port 928 nsew signal input
rlabel metal3 s 0 10864 400 10920 6 x_end[503]
port 929 nsew signal input
rlabel metal3 s 0 10752 400 10808 6 x_end[504]
port 930 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 x_end[505]
port 931 nsew signal input
rlabel metal3 s 0 10528 400 10584 6 x_end[506]
port 932 nsew signal input
rlabel metal3 s 0 10416 400 10472 6 x_end[507]
port 933 nsew signal input
rlabel metal3 s 0 10304 400 10360 6 x_end[508]
port 934 nsew signal input
rlabel metal3 s 0 10192 400 10248 6 x_end[509]
port 935 nsew signal input
rlabel metal3 s 0 61600 400 61656 6 x_end[50]
port 936 nsew signal input
rlabel metal3 s 0 10080 400 10136 6 x_end[510]
port 937 nsew signal input
rlabel metal3 s 0 9968 400 10024 6 x_end[511]
port 938 nsew signal input
rlabel metal3 s 0 61488 400 61544 6 x_end[51]
port 939 nsew signal input
rlabel metal3 s 0 61376 400 61432 6 x_end[52]
port 940 nsew signal input
rlabel metal3 s 0 61264 400 61320 6 x_end[53]
port 941 nsew signal input
rlabel metal3 s 0 61152 400 61208 6 x_end[54]
port 942 nsew signal input
rlabel metal3 s 0 61040 400 61096 6 x_end[55]
port 943 nsew signal input
rlabel metal3 s 0 60928 400 60984 6 x_end[56]
port 944 nsew signal input
rlabel metal3 s 0 60816 400 60872 6 x_end[57]
port 945 nsew signal input
rlabel metal3 s 0 60704 400 60760 6 x_end[58]
port 946 nsew signal input
rlabel metal3 s 0 60592 400 60648 6 x_end[59]
port 947 nsew signal input
rlabel metal3 s 0 66640 400 66696 6 x_end[5]
port 948 nsew signal input
rlabel metal3 s 0 60480 400 60536 6 x_end[60]
port 949 nsew signal input
rlabel metal3 s 0 60368 400 60424 6 x_end[61]
port 950 nsew signal input
rlabel metal3 s 0 60256 400 60312 6 x_end[62]
port 951 nsew signal input
rlabel metal3 s 0 60144 400 60200 6 x_end[63]
port 952 nsew signal input
rlabel metal3 s 0 60032 400 60088 6 x_end[64]
port 953 nsew signal input
rlabel metal3 s 0 59920 400 59976 6 x_end[65]
port 954 nsew signal input
rlabel metal3 s 0 59808 400 59864 6 x_end[66]
port 955 nsew signal input
rlabel metal3 s 0 59696 400 59752 6 x_end[67]
port 956 nsew signal input
rlabel metal3 s 0 59584 400 59640 6 x_end[68]
port 957 nsew signal input
rlabel metal3 s 0 59472 400 59528 6 x_end[69]
port 958 nsew signal input
rlabel metal3 s 0 66528 400 66584 6 x_end[6]
port 959 nsew signal input
rlabel metal3 s 0 59360 400 59416 6 x_end[70]
port 960 nsew signal input
rlabel metal3 s 0 59248 400 59304 6 x_end[71]
port 961 nsew signal input
rlabel metal3 s 0 59136 400 59192 6 x_end[72]
port 962 nsew signal input
rlabel metal3 s 0 59024 400 59080 6 x_end[73]
port 963 nsew signal input
rlabel metal3 s 0 58912 400 58968 6 x_end[74]
port 964 nsew signal input
rlabel metal3 s 0 58800 400 58856 6 x_end[75]
port 965 nsew signal input
rlabel metal3 s 0 58688 400 58744 6 x_end[76]
port 966 nsew signal input
rlabel metal3 s 0 58576 400 58632 6 x_end[77]
port 967 nsew signal input
rlabel metal3 s 0 58464 400 58520 6 x_end[78]
port 968 nsew signal input
rlabel metal3 s 0 58352 400 58408 6 x_end[79]
port 969 nsew signal input
rlabel metal3 s 0 66416 400 66472 6 x_end[7]
port 970 nsew signal input
rlabel metal3 s 0 58240 400 58296 6 x_end[80]
port 971 nsew signal input
rlabel metal3 s 0 58128 400 58184 6 x_end[81]
port 972 nsew signal input
rlabel metal3 s 0 58016 400 58072 6 x_end[82]
port 973 nsew signal input
rlabel metal3 s 0 57904 400 57960 6 x_end[83]
port 974 nsew signal input
rlabel metal3 s 0 57792 400 57848 6 x_end[84]
port 975 nsew signal input
rlabel metal3 s 0 57680 400 57736 6 x_end[85]
port 976 nsew signal input
rlabel metal3 s 0 57568 400 57624 6 x_end[86]
port 977 nsew signal input
rlabel metal3 s 0 57456 400 57512 6 x_end[87]
port 978 nsew signal input
rlabel metal3 s 0 57344 400 57400 6 x_end[88]
port 979 nsew signal input
rlabel metal3 s 0 57232 400 57288 6 x_end[89]
port 980 nsew signal input
rlabel metal3 s 0 66304 400 66360 6 x_end[8]
port 981 nsew signal input
rlabel metal3 s 0 57120 400 57176 6 x_end[90]
port 982 nsew signal input
rlabel metal3 s 0 57008 400 57064 6 x_end[91]
port 983 nsew signal input
rlabel metal3 s 0 56896 400 56952 6 x_end[92]
port 984 nsew signal input
rlabel metal3 s 0 56784 400 56840 6 x_end[93]
port 985 nsew signal input
rlabel metal3 s 0 56672 400 56728 6 x_end[94]
port 986 nsew signal input
rlabel metal3 s 0 56560 400 56616 6 x_end[95]
port 987 nsew signal input
rlabel metal3 s 0 56448 400 56504 6 x_end[96]
port 988 nsew signal input
rlabel metal3 s 0 56336 400 56392 6 x_end[97]
port 989 nsew signal input
rlabel metal3 s 0 56224 400 56280 6 x_end[98]
port 990 nsew signal input
rlabel metal3 s 0 56112 400 56168 6 x_end[99]
port 991 nsew signal input
rlabel metal3 s 0 66192 400 66248 6 x_end[9]
port 992 nsew signal input
rlabel metal3 s 279600 12656 280000 12712 6 x_start[0]
port 993 nsew signal input
rlabel metal3 s 279600 23856 280000 23912 6 x_start[100]
port 994 nsew signal input
rlabel metal3 s 279600 23968 280000 24024 6 x_start[101]
port 995 nsew signal input
rlabel metal3 s 279600 24080 280000 24136 6 x_start[102]
port 996 nsew signal input
rlabel metal3 s 279600 24192 280000 24248 6 x_start[103]
port 997 nsew signal input
rlabel metal3 s 279600 24304 280000 24360 6 x_start[104]
port 998 nsew signal input
rlabel metal3 s 279600 24416 280000 24472 6 x_start[105]
port 999 nsew signal input
rlabel metal3 s 279600 24528 280000 24584 6 x_start[106]
port 1000 nsew signal input
rlabel metal3 s 279600 24640 280000 24696 6 x_start[107]
port 1001 nsew signal input
rlabel metal3 s 279600 24752 280000 24808 6 x_start[108]
port 1002 nsew signal input
rlabel metal3 s 279600 24864 280000 24920 6 x_start[109]
port 1003 nsew signal input
rlabel metal3 s 279600 13776 280000 13832 6 x_start[10]
port 1004 nsew signal input
rlabel metal3 s 279600 24976 280000 25032 6 x_start[110]
port 1005 nsew signal input
rlabel metal3 s 279600 25088 280000 25144 6 x_start[111]
port 1006 nsew signal input
rlabel metal3 s 279600 25200 280000 25256 6 x_start[112]
port 1007 nsew signal input
rlabel metal3 s 279600 25312 280000 25368 6 x_start[113]
port 1008 nsew signal input
rlabel metal3 s 279600 25424 280000 25480 6 x_start[114]
port 1009 nsew signal input
rlabel metal3 s 279600 25536 280000 25592 6 x_start[115]
port 1010 nsew signal input
rlabel metal3 s 279600 25648 280000 25704 6 x_start[116]
port 1011 nsew signal input
rlabel metal3 s 279600 25760 280000 25816 6 x_start[117]
port 1012 nsew signal input
rlabel metal3 s 279600 25872 280000 25928 6 x_start[118]
port 1013 nsew signal input
rlabel metal3 s 279600 25984 280000 26040 6 x_start[119]
port 1014 nsew signal input
rlabel metal3 s 279600 13888 280000 13944 6 x_start[11]
port 1015 nsew signal input
rlabel metal3 s 279600 26096 280000 26152 6 x_start[120]
port 1016 nsew signal input
rlabel metal3 s 279600 26208 280000 26264 6 x_start[121]
port 1017 nsew signal input
rlabel metal3 s 279600 26320 280000 26376 6 x_start[122]
port 1018 nsew signal input
rlabel metal3 s 279600 26432 280000 26488 6 x_start[123]
port 1019 nsew signal input
rlabel metal3 s 279600 26544 280000 26600 6 x_start[124]
port 1020 nsew signal input
rlabel metal3 s 279600 26656 280000 26712 6 x_start[125]
port 1021 nsew signal input
rlabel metal3 s 279600 26768 280000 26824 6 x_start[126]
port 1022 nsew signal input
rlabel metal3 s 279600 26880 280000 26936 6 x_start[127]
port 1023 nsew signal input
rlabel metal3 s 279600 26992 280000 27048 6 x_start[128]
port 1024 nsew signal input
rlabel metal3 s 279600 27104 280000 27160 6 x_start[129]
port 1025 nsew signal input
rlabel metal3 s 279600 14000 280000 14056 6 x_start[12]
port 1026 nsew signal input
rlabel metal3 s 279600 27216 280000 27272 6 x_start[130]
port 1027 nsew signal input
rlabel metal3 s 279600 27328 280000 27384 6 x_start[131]
port 1028 nsew signal input
rlabel metal3 s 279600 27440 280000 27496 6 x_start[132]
port 1029 nsew signal input
rlabel metal3 s 279600 27552 280000 27608 6 x_start[133]
port 1030 nsew signal input
rlabel metal3 s 279600 27664 280000 27720 6 x_start[134]
port 1031 nsew signal input
rlabel metal3 s 279600 27776 280000 27832 6 x_start[135]
port 1032 nsew signal input
rlabel metal3 s 279600 27888 280000 27944 6 x_start[136]
port 1033 nsew signal input
rlabel metal3 s 279600 28000 280000 28056 6 x_start[137]
port 1034 nsew signal input
rlabel metal3 s 279600 28112 280000 28168 6 x_start[138]
port 1035 nsew signal input
rlabel metal3 s 279600 28224 280000 28280 6 x_start[139]
port 1036 nsew signal input
rlabel metal3 s 279600 14112 280000 14168 6 x_start[13]
port 1037 nsew signal input
rlabel metal3 s 279600 28336 280000 28392 6 x_start[140]
port 1038 nsew signal input
rlabel metal3 s 279600 28448 280000 28504 6 x_start[141]
port 1039 nsew signal input
rlabel metal3 s 279600 28560 280000 28616 6 x_start[142]
port 1040 nsew signal input
rlabel metal3 s 279600 28672 280000 28728 6 x_start[143]
port 1041 nsew signal input
rlabel metal3 s 279600 28784 280000 28840 6 x_start[144]
port 1042 nsew signal input
rlabel metal3 s 279600 28896 280000 28952 6 x_start[145]
port 1043 nsew signal input
rlabel metal3 s 279600 29008 280000 29064 6 x_start[146]
port 1044 nsew signal input
rlabel metal3 s 279600 29120 280000 29176 6 x_start[147]
port 1045 nsew signal input
rlabel metal3 s 279600 29232 280000 29288 6 x_start[148]
port 1046 nsew signal input
rlabel metal3 s 279600 29344 280000 29400 6 x_start[149]
port 1047 nsew signal input
rlabel metal3 s 279600 14224 280000 14280 6 x_start[14]
port 1048 nsew signal input
rlabel metal3 s 279600 29456 280000 29512 6 x_start[150]
port 1049 nsew signal input
rlabel metal3 s 279600 29568 280000 29624 6 x_start[151]
port 1050 nsew signal input
rlabel metal3 s 279600 29680 280000 29736 6 x_start[152]
port 1051 nsew signal input
rlabel metal3 s 279600 29792 280000 29848 6 x_start[153]
port 1052 nsew signal input
rlabel metal3 s 279600 29904 280000 29960 6 x_start[154]
port 1053 nsew signal input
rlabel metal3 s 279600 30016 280000 30072 6 x_start[155]
port 1054 nsew signal input
rlabel metal3 s 279600 30128 280000 30184 6 x_start[156]
port 1055 nsew signal input
rlabel metal3 s 279600 30240 280000 30296 6 x_start[157]
port 1056 nsew signal input
rlabel metal3 s 279600 30352 280000 30408 6 x_start[158]
port 1057 nsew signal input
rlabel metal3 s 279600 30464 280000 30520 6 x_start[159]
port 1058 nsew signal input
rlabel metal3 s 279600 14336 280000 14392 6 x_start[15]
port 1059 nsew signal input
rlabel metal3 s 279600 30576 280000 30632 6 x_start[160]
port 1060 nsew signal input
rlabel metal3 s 279600 30688 280000 30744 6 x_start[161]
port 1061 nsew signal input
rlabel metal3 s 279600 30800 280000 30856 6 x_start[162]
port 1062 nsew signal input
rlabel metal3 s 279600 30912 280000 30968 6 x_start[163]
port 1063 nsew signal input
rlabel metal3 s 279600 31024 280000 31080 6 x_start[164]
port 1064 nsew signal input
rlabel metal3 s 279600 31136 280000 31192 6 x_start[165]
port 1065 nsew signal input
rlabel metal3 s 279600 31248 280000 31304 6 x_start[166]
port 1066 nsew signal input
rlabel metal3 s 279600 31360 280000 31416 6 x_start[167]
port 1067 nsew signal input
rlabel metal3 s 279600 31472 280000 31528 6 x_start[168]
port 1068 nsew signal input
rlabel metal3 s 279600 31584 280000 31640 6 x_start[169]
port 1069 nsew signal input
rlabel metal3 s 279600 14448 280000 14504 6 x_start[16]
port 1070 nsew signal input
rlabel metal3 s 279600 31696 280000 31752 6 x_start[170]
port 1071 nsew signal input
rlabel metal3 s 279600 31808 280000 31864 6 x_start[171]
port 1072 nsew signal input
rlabel metal3 s 279600 31920 280000 31976 6 x_start[172]
port 1073 nsew signal input
rlabel metal3 s 279600 32032 280000 32088 6 x_start[173]
port 1074 nsew signal input
rlabel metal3 s 279600 32144 280000 32200 6 x_start[174]
port 1075 nsew signal input
rlabel metal3 s 279600 32256 280000 32312 6 x_start[175]
port 1076 nsew signal input
rlabel metal3 s 279600 32368 280000 32424 6 x_start[176]
port 1077 nsew signal input
rlabel metal3 s 279600 32480 280000 32536 6 x_start[177]
port 1078 nsew signal input
rlabel metal3 s 279600 32592 280000 32648 6 x_start[178]
port 1079 nsew signal input
rlabel metal3 s 279600 32704 280000 32760 6 x_start[179]
port 1080 nsew signal input
rlabel metal3 s 279600 14560 280000 14616 6 x_start[17]
port 1081 nsew signal input
rlabel metal3 s 279600 32816 280000 32872 6 x_start[180]
port 1082 nsew signal input
rlabel metal3 s 279600 32928 280000 32984 6 x_start[181]
port 1083 nsew signal input
rlabel metal3 s 279600 33040 280000 33096 6 x_start[182]
port 1084 nsew signal input
rlabel metal3 s 279600 33152 280000 33208 6 x_start[183]
port 1085 nsew signal input
rlabel metal3 s 279600 33264 280000 33320 6 x_start[184]
port 1086 nsew signal input
rlabel metal3 s 279600 33376 280000 33432 6 x_start[185]
port 1087 nsew signal input
rlabel metal3 s 279600 33488 280000 33544 6 x_start[186]
port 1088 nsew signal input
rlabel metal3 s 279600 33600 280000 33656 6 x_start[187]
port 1089 nsew signal input
rlabel metal3 s 279600 33712 280000 33768 6 x_start[188]
port 1090 nsew signal input
rlabel metal3 s 279600 33824 280000 33880 6 x_start[189]
port 1091 nsew signal input
rlabel metal3 s 279600 14672 280000 14728 6 x_start[18]
port 1092 nsew signal input
rlabel metal3 s 279600 33936 280000 33992 6 x_start[190]
port 1093 nsew signal input
rlabel metal3 s 279600 34048 280000 34104 6 x_start[191]
port 1094 nsew signal input
rlabel metal3 s 279600 34160 280000 34216 6 x_start[192]
port 1095 nsew signal input
rlabel metal3 s 279600 34272 280000 34328 6 x_start[193]
port 1096 nsew signal input
rlabel metal3 s 279600 34384 280000 34440 6 x_start[194]
port 1097 nsew signal input
rlabel metal3 s 279600 34496 280000 34552 6 x_start[195]
port 1098 nsew signal input
rlabel metal3 s 279600 34608 280000 34664 6 x_start[196]
port 1099 nsew signal input
rlabel metal3 s 279600 34720 280000 34776 6 x_start[197]
port 1100 nsew signal input
rlabel metal3 s 279600 34832 280000 34888 6 x_start[198]
port 1101 nsew signal input
rlabel metal3 s 279600 34944 280000 35000 6 x_start[199]
port 1102 nsew signal input
rlabel metal3 s 279600 14784 280000 14840 6 x_start[19]
port 1103 nsew signal input
rlabel metal3 s 279600 12768 280000 12824 6 x_start[1]
port 1104 nsew signal input
rlabel metal3 s 279600 35056 280000 35112 6 x_start[200]
port 1105 nsew signal input
rlabel metal3 s 279600 35168 280000 35224 6 x_start[201]
port 1106 nsew signal input
rlabel metal3 s 279600 35280 280000 35336 6 x_start[202]
port 1107 nsew signal input
rlabel metal3 s 279600 35392 280000 35448 6 x_start[203]
port 1108 nsew signal input
rlabel metal3 s 279600 35504 280000 35560 6 x_start[204]
port 1109 nsew signal input
rlabel metal3 s 279600 35616 280000 35672 6 x_start[205]
port 1110 nsew signal input
rlabel metal3 s 279600 35728 280000 35784 6 x_start[206]
port 1111 nsew signal input
rlabel metal3 s 279600 35840 280000 35896 6 x_start[207]
port 1112 nsew signal input
rlabel metal3 s 279600 35952 280000 36008 6 x_start[208]
port 1113 nsew signal input
rlabel metal3 s 279600 36064 280000 36120 6 x_start[209]
port 1114 nsew signal input
rlabel metal3 s 279600 14896 280000 14952 6 x_start[20]
port 1115 nsew signal input
rlabel metal3 s 279600 36176 280000 36232 6 x_start[210]
port 1116 nsew signal input
rlabel metal3 s 279600 36288 280000 36344 6 x_start[211]
port 1117 nsew signal input
rlabel metal3 s 279600 36400 280000 36456 6 x_start[212]
port 1118 nsew signal input
rlabel metal3 s 279600 36512 280000 36568 6 x_start[213]
port 1119 nsew signal input
rlabel metal3 s 279600 36624 280000 36680 6 x_start[214]
port 1120 nsew signal input
rlabel metal3 s 279600 36736 280000 36792 6 x_start[215]
port 1121 nsew signal input
rlabel metal3 s 279600 36848 280000 36904 6 x_start[216]
port 1122 nsew signal input
rlabel metal3 s 279600 36960 280000 37016 6 x_start[217]
port 1123 nsew signal input
rlabel metal3 s 279600 37072 280000 37128 6 x_start[218]
port 1124 nsew signal input
rlabel metal3 s 279600 37184 280000 37240 6 x_start[219]
port 1125 nsew signal input
rlabel metal3 s 279600 15008 280000 15064 6 x_start[21]
port 1126 nsew signal input
rlabel metal3 s 279600 37296 280000 37352 6 x_start[220]
port 1127 nsew signal input
rlabel metal3 s 279600 37408 280000 37464 6 x_start[221]
port 1128 nsew signal input
rlabel metal3 s 279600 37520 280000 37576 6 x_start[222]
port 1129 nsew signal input
rlabel metal3 s 279600 37632 280000 37688 6 x_start[223]
port 1130 nsew signal input
rlabel metal3 s 279600 37744 280000 37800 6 x_start[224]
port 1131 nsew signal input
rlabel metal3 s 279600 37856 280000 37912 6 x_start[225]
port 1132 nsew signal input
rlabel metal3 s 279600 37968 280000 38024 6 x_start[226]
port 1133 nsew signal input
rlabel metal3 s 279600 38080 280000 38136 6 x_start[227]
port 1134 nsew signal input
rlabel metal3 s 279600 38192 280000 38248 6 x_start[228]
port 1135 nsew signal input
rlabel metal3 s 279600 38304 280000 38360 6 x_start[229]
port 1136 nsew signal input
rlabel metal3 s 279600 15120 280000 15176 6 x_start[22]
port 1137 nsew signal input
rlabel metal3 s 279600 38416 280000 38472 6 x_start[230]
port 1138 nsew signal input
rlabel metal3 s 279600 38528 280000 38584 6 x_start[231]
port 1139 nsew signal input
rlabel metal3 s 279600 38640 280000 38696 6 x_start[232]
port 1140 nsew signal input
rlabel metal3 s 279600 38752 280000 38808 6 x_start[233]
port 1141 nsew signal input
rlabel metal3 s 279600 38864 280000 38920 6 x_start[234]
port 1142 nsew signal input
rlabel metal3 s 279600 38976 280000 39032 6 x_start[235]
port 1143 nsew signal input
rlabel metal3 s 279600 39088 280000 39144 6 x_start[236]
port 1144 nsew signal input
rlabel metal3 s 279600 39200 280000 39256 6 x_start[237]
port 1145 nsew signal input
rlabel metal3 s 279600 39312 280000 39368 6 x_start[238]
port 1146 nsew signal input
rlabel metal3 s 279600 39424 280000 39480 6 x_start[239]
port 1147 nsew signal input
rlabel metal3 s 279600 15232 280000 15288 6 x_start[23]
port 1148 nsew signal input
rlabel metal3 s 279600 39536 280000 39592 6 x_start[240]
port 1149 nsew signal input
rlabel metal3 s 279600 39648 280000 39704 6 x_start[241]
port 1150 nsew signal input
rlabel metal3 s 279600 39760 280000 39816 6 x_start[242]
port 1151 nsew signal input
rlabel metal3 s 279600 39872 280000 39928 6 x_start[243]
port 1152 nsew signal input
rlabel metal3 s 279600 39984 280000 40040 6 x_start[244]
port 1153 nsew signal input
rlabel metal3 s 279600 40096 280000 40152 6 x_start[245]
port 1154 nsew signal input
rlabel metal3 s 279600 40208 280000 40264 6 x_start[246]
port 1155 nsew signal input
rlabel metal3 s 279600 40320 280000 40376 6 x_start[247]
port 1156 nsew signal input
rlabel metal3 s 279600 40432 280000 40488 6 x_start[248]
port 1157 nsew signal input
rlabel metal3 s 279600 40544 280000 40600 6 x_start[249]
port 1158 nsew signal input
rlabel metal3 s 279600 15344 280000 15400 6 x_start[24]
port 1159 nsew signal input
rlabel metal3 s 279600 40656 280000 40712 6 x_start[250]
port 1160 nsew signal input
rlabel metal3 s 279600 40768 280000 40824 6 x_start[251]
port 1161 nsew signal input
rlabel metal3 s 279600 40880 280000 40936 6 x_start[252]
port 1162 nsew signal input
rlabel metal3 s 279600 40992 280000 41048 6 x_start[253]
port 1163 nsew signal input
rlabel metal3 s 279600 41104 280000 41160 6 x_start[254]
port 1164 nsew signal input
rlabel metal3 s 279600 41216 280000 41272 6 x_start[255]
port 1165 nsew signal input
rlabel metal3 s 279600 41328 280000 41384 6 x_start[256]
port 1166 nsew signal input
rlabel metal3 s 279600 41440 280000 41496 6 x_start[257]
port 1167 nsew signal input
rlabel metal3 s 279600 41552 280000 41608 6 x_start[258]
port 1168 nsew signal input
rlabel metal3 s 279600 41664 280000 41720 6 x_start[259]
port 1169 nsew signal input
rlabel metal3 s 279600 15456 280000 15512 6 x_start[25]
port 1170 nsew signal input
rlabel metal3 s 279600 41776 280000 41832 6 x_start[260]
port 1171 nsew signal input
rlabel metal3 s 279600 41888 280000 41944 6 x_start[261]
port 1172 nsew signal input
rlabel metal3 s 279600 42000 280000 42056 6 x_start[262]
port 1173 nsew signal input
rlabel metal3 s 279600 42112 280000 42168 6 x_start[263]
port 1174 nsew signal input
rlabel metal3 s 279600 42224 280000 42280 6 x_start[264]
port 1175 nsew signal input
rlabel metal3 s 279600 42336 280000 42392 6 x_start[265]
port 1176 nsew signal input
rlabel metal3 s 279600 42448 280000 42504 6 x_start[266]
port 1177 nsew signal input
rlabel metal3 s 279600 42560 280000 42616 6 x_start[267]
port 1178 nsew signal input
rlabel metal3 s 279600 42672 280000 42728 6 x_start[268]
port 1179 nsew signal input
rlabel metal3 s 279600 42784 280000 42840 6 x_start[269]
port 1180 nsew signal input
rlabel metal3 s 279600 15568 280000 15624 6 x_start[26]
port 1181 nsew signal input
rlabel metal3 s 279600 42896 280000 42952 6 x_start[270]
port 1182 nsew signal input
rlabel metal3 s 279600 43008 280000 43064 6 x_start[271]
port 1183 nsew signal input
rlabel metal3 s 279600 43120 280000 43176 6 x_start[272]
port 1184 nsew signal input
rlabel metal3 s 279600 43232 280000 43288 6 x_start[273]
port 1185 nsew signal input
rlabel metal3 s 279600 43344 280000 43400 6 x_start[274]
port 1186 nsew signal input
rlabel metal3 s 279600 43456 280000 43512 6 x_start[275]
port 1187 nsew signal input
rlabel metal3 s 279600 43568 280000 43624 6 x_start[276]
port 1188 nsew signal input
rlabel metal3 s 279600 43680 280000 43736 6 x_start[277]
port 1189 nsew signal input
rlabel metal3 s 279600 43792 280000 43848 6 x_start[278]
port 1190 nsew signal input
rlabel metal3 s 279600 43904 280000 43960 6 x_start[279]
port 1191 nsew signal input
rlabel metal3 s 279600 15680 280000 15736 6 x_start[27]
port 1192 nsew signal input
rlabel metal3 s 279600 44016 280000 44072 6 x_start[280]
port 1193 nsew signal input
rlabel metal3 s 279600 44128 280000 44184 6 x_start[281]
port 1194 nsew signal input
rlabel metal3 s 279600 44240 280000 44296 6 x_start[282]
port 1195 nsew signal input
rlabel metal3 s 279600 44352 280000 44408 6 x_start[283]
port 1196 nsew signal input
rlabel metal3 s 279600 44464 280000 44520 6 x_start[284]
port 1197 nsew signal input
rlabel metal3 s 279600 44576 280000 44632 6 x_start[285]
port 1198 nsew signal input
rlabel metal3 s 279600 44688 280000 44744 6 x_start[286]
port 1199 nsew signal input
rlabel metal3 s 279600 44800 280000 44856 6 x_start[287]
port 1200 nsew signal input
rlabel metal3 s 279600 44912 280000 44968 6 x_start[288]
port 1201 nsew signal input
rlabel metal3 s 279600 45024 280000 45080 6 x_start[289]
port 1202 nsew signal input
rlabel metal3 s 279600 15792 280000 15848 6 x_start[28]
port 1203 nsew signal input
rlabel metal3 s 279600 45136 280000 45192 6 x_start[290]
port 1204 nsew signal input
rlabel metal3 s 279600 45248 280000 45304 6 x_start[291]
port 1205 nsew signal input
rlabel metal3 s 279600 45360 280000 45416 6 x_start[292]
port 1206 nsew signal input
rlabel metal3 s 279600 45472 280000 45528 6 x_start[293]
port 1207 nsew signal input
rlabel metal3 s 279600 45584 280000 45640 6 x_start[294]
port 1208 nsew signal input
rlabel metal3 s 279600 45696 280000 45752 6 x_start[295]
port 1209 nsew signal input
rlabel metal3 s 279600 45808 280000 45864 6 x_start[296]
port 1210 nsew signal input
rlabel metal3 s 279600 45920 280000 45976 6 x_start[297]
port 1211 nsew signal input
rlabel metal3 s 279600 46032 280000 46088 6 x_start[298]
port 1212 nsew signal input
rlabel metal3 s 279600 46144 280000 46200 6 x_start[299]
port 1213 nsew signal input
rlabel metal3 s 279600 15904 280000 15960 6 x_start[29]
port 1214 nsew signal input
rlabel metal3 s 279600 12880 280000 12936 6 x_start[2]
port 1215 nsew signal input
rlabel metal3 s 279600 46256 280000 46312 6 x_start[300]
port 1216 nsew signal input
rlabel metal3 s 279600 46368 280000 46424 6 x_start[301]
port 1217 nsew signal input
rlabel metal3 s 279600 46480 280000 46536 6 x_start[302]
port 1218 nsew signal input
rlabel metal3 s 279600 46592 280000 46648 6 x_start[303]
port 1219 nsew signal input
rlabel metal3 s 279600 46704 280000 46760 6 x_start[304]
port 1220 nsew signal input
rlabel metal3 s 279600 46816 280000 46872 6 x_start[305]
port 1221 nsew signal input
rlabel metal3 s 279600 46928 280000 46984 6 x_start[306]
port 1222 nsew signal input
rlabel metal3 s 279600 47040 280000 47096 6 x_start[307]
port 1223 nsew signal input
rlabel metal3 s 279600 47152 280000 47208 6 x_start[308]
port 1224 nsew signal input
rlabel metal3 s 279600 47264 280000 47320 6 x_start[309]
port 1225 nsew signal input
rlabel metal3 s 279600 16016 280000 16072 6 x_start[30]
port 1226 nsew signal input
rlabel metal3 s 279600 47376 280000 47432 6 x_start[310]
port 1227 nsew signal input
rlabel metal3 s 279600 47488 280000 47544 6 x_start[311]
port 1228 nsew signal input
rlabel metal3 s 279600 47600 280000 47656 6 x_start[312]
port 1229 nsew signal input
rlabel metal3 s 279600 47712 280000 47768 6 x_start[313]
port 1230 nsew signal input
rlabel metal3 s 279600 47824 280000 47880 6 x_start[314]
port 1231 nsew signal input
rlabel metal3 s 279600 47936 280000 47992 6 x_start[315]
port 1232 nsew signal input
rlabel metal3 s 279600 48048 280000 48104 6 x_start[316]
port 1233 nsew signal input
rlabel metal3 s 279600 48160 280000 48216 6 x_start[317]
port 1234 nsew signal input
rlabel metal3 s 279600 48272 280000 48328 6 x_start[318]
port 1235 nsew signal input
rlabel metal3 s 279600 48384 280000 48440 6 x_start[319]
port 1236 nsew signal input
rlabel metal3 s 279600 16128 280000 16184 6 x_start[31]
port 1237 nsew signal input
rlabel metal3 s 279600 48496 280000 48552 6 x_start[320]
port 1238 nsew signal input
rlabel metal3 s 279600 48608 280000 48664 6 x_start[321]
port 1239 nsew signal input
rlabel metal3 s 279600 48720 280000 48776 6 x_start[322]
port 1240 nsew signal input
rlabel metal3 s 279600 48832 280000 48888 6 x_start[323]
port 1241 nsew signal input
rlabel metal3 s 279600 48944 280000 49000 6 x_start[324]
port 1242 nsew signal input
rlabel metal3 s 279600 49056 280000 49112 6 x_start[325]
port 1243 nsew signal input
rlabel metal3 s 279600 49168 280000 49224 6 x_start[326]
port 1244 nsew signal input
rlabel metal3 s 279600 49280 280000 49336 6 x_start[327]
port 1245 nsew signal input
rlabel metal3 s 279600 49392 280000 49448 6 x_start[328]
port 1246 nsew signal input
rlabel metal3 s 279600 49504 280000 49560 6 x_start[329]
port 1247 nsew signal input
rlabel metal3 s 279600 16240 280000 16296 6 x_start[32]
port 1248 nsew signal input
rlabel metal3 s 279600 49616 280000 49672 6 x_start[330]
port 1249 nsew signal input
rlabel metal3 s 279600 49728 280000 49784 6 x_start[331]
port 1250 nsew signal input
rlabel metal3 s 279600 49840 280000 49896 6 x_start[332]
port 1251 nsew signal input
rlabel metal3 s 279600 49952 280000 50008 6 x_start[333]
port 1252 nsew signal input
rlabel metal3 s 279600 50064 280000 50120 6 x_start[334]
port 1253 nsew signal input
rlabel metal3 s 279600 50176 280000 50232 6 x_start[335]
port 1254 nsew signal input
rlabel metal3 s 279600 50288 280000 50344 6 x_start[336]
port 1255 nsew signal input
rlabel metal3 s 279600 50400 280000 50456 6 x_start[337]
port 1256 nsew signal input
rlabel metal3 s 279600 50512 280000 50568 6 x_start[338]
port 1257 nsew signal input
rlabel metal3 s 279600 50624 280000 50680 6 x_start[339]
port 1258 nsew signal input
rlabel metal3 s 279600 16352 280000 16408 6 x_start[33]
port 1259 nsew signal input
rlabel metal3 s 279600 50736 280000 50792 6 x_start[340]
port 1260 nsew signal input
rlabel metal3 s 279600 50848 280000 50904 6 x_start[341]
port 1261 nsew signal input
rlabel metal3 s 279600 50960 280000 51016 6 x_start[342]
port 1262 nsew signal input
rlabel metal3 s 279600 51072 280000 51128 6 x_start[343]
port 1263 nsew signal input
rlabel metal3 s 279600 51184 280000 51240 6 x_start[344]
port 1264 nsew signal input
rlabel metal3 s 279600 51296 280000 51352 6 x_start[345]
port 1265 nsew signal input
rlabel metal3 s 279600 51408 280000 51464 6 x_start[346]
port 1266 nsew signal input
rlabel metal3 s 279600 51520 280000 51576 6 x_start[347]
port 1267 nsew signal input
rlabel metal3 s 279600 51632 280000 51688 6 x_start[348]
port 1268 nsew signal input
rlabel metal3 s 279600 51744 280000 51800 6 x_start[349]
port 1269 nsew signal input
rlabel metal3 s 279600 16464 280000 16520 6 x_start[34]
port 1270 nsew signal input
rlabel metal3 s 279600 51856 280000 51912 6 x_start[350]
port 1271 nsew signal input
rlabel metal3 s 279600 51968 280000 52024 6 x_start[351]
port 1272 nsew signal input
rlabel metal3 s 279600 52080 280000 52136 6 x_start[352]
port 1273 nsew signal input
rlabel metal3 s 279600 52192 280000 52248 6 x_start[353]
port 1274 nsew signal input
rlabel metal3 s 279600 52304 280000 52360 6 x_start[354]
port 1275 nsew signal input
rlabel metal3 s 279600 52416 280000 52472 6 x_start[355]
port 1276 nsew signal input
rlabel metal3 s 279600 52528 280000 52584 6 x_start[356]
port 1277 nsew signal input
rlabel metal3 s 279600 52640 280000 52696 6 x_start[357]
port 1278 nsew signal input
rlabel metal3 s 279600 52752 280000 52808 6 x_start[358]
port 1279 nsew signal input
rlabel metal3 s 279600 52864 280000 52920 6 x_start[359]
port 1280 nsew signal input
rlabel metal3 s 279600 16576 280000 16632 6 x_start[35]
port 1281 nsew signal input
rlabel metal3 s 279600 52976 280000 53032 6 x_start[360]
port 1282 nsew signal input
rlabel metal3 s 279600 53088 280000 53144 6 x_start[361]
port 1283 nsew signal input
rlabel metal3 s 279600 53200 280000 53256 6 x_start[362]
port 1284 nsew signal input
rlabel metal3 s 279600 53312 280000 53368 6 x_start[363]
port 1285 nsew signal input
rlabel metal3 s 279600 53424 280000 53480 6 x_start[364]
port 1286 nsew signal input
rlabel metal3 s 279600 53536 280000 53592 6 x_start[365]
port 1287 nsew signal input
rlabel metal3 s 279600 53648 280000 53704 6 x_start[366]
port 1288 nsew signal input
rlabel metal3 s 279600 53760 280000 53816 6 x_start[367]
port 1289 nsew signal input
rlabel metal3 s 279600 53872 280000 53928 6 x_start[368]
port 1290 nsew signal input
rlabel metal3 s 279600 53984 280000 54040 6 x_start[369]
port 1291 nsew signal input
rlabel metal3 s 279600 16688 280000 16744 6 x_start[36]
port 1292 nsew signal input
rlabel metal3 s 279600 54096 280000 54152 6 x_start[370]
port 1293 nsew signal input
rlabel metal3 s 279600 54208 280000 54264 6 x_start[371]
port 1294 nsew signal input
rlabel metal3 s 279600 54320 280000 54376 6 x_start[372]
port 1295 nsew signal input
rlabel metal3 s 279600 54432 280000 54488 6 x_start[373]
port 1296 nsew signal input
rlabel metal3 s 279600 54544 280000 54600 6 x_start[374]
port 1297 nsew signal input
rlabel metal3 s 279600 54656 280000 54712 6 x_start[375]
port 1298 nsew signal input
rlabel metal3 s 279600 54768 280000 54824 6 x_start[376]
port 1299 nsew signal input
rlabel metal3 s 279600 54880 280000 54936 6 x_start[377]
port 1300 nsew signal input
rlabel metal3 s 279600 54992 280000 55048 6 x_start[378]
port 1301 nsew signal input
rlabel metal3 s 279600 55104 280000 55160 6 x_start[379]
port 1302 nsew signal input
rlabel metal3 s 279600 16800 280000 16856 6 x_start[37]
port 1303 nsew signal input
rlabel metal3 s 279600 55216 280000 55272 6 x_start[380]
port 1304 nsew signal input
rlabel metal3 s 279600 55328 280000 55384 6 x_start[381]
port 1305 nsew signal input
rlabel metal3 s 279600 55440 280000 55496 6 x_start[382]
port 1306 nsew signal input
rlabel metal3 s 279600 55552 280000 55608 6 x_start[383]
port 1307 nsew signal input
rlabel metal3 s 279600 55664 280000 55720 6 x_start[384]
port 1308 nsew signal input
rlabel metal3 s 279600 55776 280000 55832 6 x_start[385]
port 1309 nsew signal input
rlabel metal3 s 279600 55888 280000 55944 6 x_start[386]
port 1310 nsew signal input
rlabel metal3 s 279600 56000 280000 56056 6 x_start[387]
port 1311 nsew signal input
rlabel metal3 s 279600 56112 280000 56168 6 x_start[388]
port 1312 nsew signal input
rlabel metal3 s 279600 56224 280000 56280 6 x_start[389]
port 1313 nsew signal input
rlabel metal3 s 279600 16912 280000 16968 6 x_start[38]
port 1314 nsew signal input
rlabel metal3 s 279600 56336 280000 56392 6 x_start[390]
port 1315 nsew signal input
rlabel metal3 s 279600 56448 280000 56504 6 x_start[391]
port 1316 nsew signal input
rlabel metal3 s 279600 56560 280000 56616 6 x_start[392]
port 1317 nsew signal input
rlabel metal3 s 279600 56672 280000 56728 6 x_start[393]
port 1318 nsew signal input
rlabel metal3 s 279600 56784 280000 56840 6 x_start[394]
port 1319 nsew signal input
rlabel metal3 s 279600 56896 280000 56952 6 x_start[395]
port 1320 nsew signal input
rlabel metal3 s 279600 57008 280000 57064 6 x_start[396]
port 1321 nsew signal input
rlabel metal3 s 279600 57120 280000 57176 6 x_start[397]
port 1322 nsew signal input
rlabel metal3 s 279600 57232 280000 57288 6 x_start[398]
port 1323 nsew signal input
rlabel metal3 s 279600 57344 280000 57400 6 x_start[399]
port 1324 nsew signal input
rlabel metal3 s 279600 17024 280000 17080 6 x_start[39]
port 1325 nsew signal input
rlabel metal3 s 279600 12992 280000 13048 6 x_start[3]
port 1326 nsew signal input
rlabel metal3 s 279600 57456 280000 57512 6 x_start[400]
port 1327 nsew signal input
rlabel metal3 s 279600 57568 280000 57624 6 x_start[401]
port 1328 nsew signal input
rlabel metal3 s 279600 57680 280000 57736 6 x_start[402]
port 1329 nsew signal input
rlabel metal3 s 279600 57792 280000 57848 6 x_start[403]
port 1330 nsew signal input
rlabel metal3 s 279600 57904 280000 57960 6 x_start[404]
port 1331 nsew signal input
rlabel metal3 s 279600 58016 280000 58072 6 x_start[405]
port 1332 nsew signal input
rlabel metal3 s 279600 58128 280000 58184 6 x_start[406]
port 1333 nsew signal input
rlabel metal3 s 279600 58240 280000 58296 6 x_start[407]
port 1334 nsew signal input
rlabel metal3 s 279600 58352 280000 58408 6 x_start[408]
port 1335 nsew signal input
rlabel metal3 s 279600 58464 280000 58520 6 x_start[409]
port 1336 nsew signal input
rlabel metal3 s 279600 17136 280000 17192 6 x_start[40]
port 1337 nsew signal input
rlabel metal3 s 279600 58576 280000 58632 6 x_start[410]
port 1338 nsew signal input
rlabel metal3 s 279600 58688 280000 58744 6 x_start[411]
port 1339 nsew signal input
rlabel metal3 s 279600 58800 280000 58856 6 x_start[412]
port 1340 nsew signal input
rlabel metal3 s 279600 58912 280000 58968 6 x_start[413]
port 1341 nsew signal input
rlabel metal3 s 279600 59024 280000 59080 6 x_start[414]
port 1342 nsew signal input
rlabel metal3 s 279600 59136 280000 59192 6 x_start[415]
port 1343 nsew signal input
rlabel metal3 s 279600 59248 280000 59304 6 x_start[416]
port 1344 nsew signal input
rlabel metal3 s 279600 59360 280000 59416 6 x_start[417]
port 1345 nsew signal input
rlabel metal3 s 279600 59472 280000 59528 6 x_start[418]
port 1346 nsew signal input
rlabel metal3 s 279600 59584 280000 59640 6 x_start[419]
port 1347 nsew signal input
rlabel metal3 s 279600 17248 280000 17304 6 x_start[41]
port 1348 nsew signal input
rlabel metal3 s 279600 59696 280000 59752 6 x_start[420]
port 1349 nsew signal input
rlabel metal3 s 279600 59808 280000 59864 6 x_start[421]
port 1350 nsew signal input
rlabel metal3 s 279600 59920 280000 59976 6 x_start[422]
port 1351 nsew signal input
rlabel metal3 s 279600 60032 280000 60088 6 x_start[423]
port 1352 nsew signal input
rlabel metal3 s 279600 60144 280000 60200 6 x_start[424]
port 1353 nsew signal input
rlabel metal3 s 279600 60256 280000 60312 6 x_start[425]
port 1354 nsew signal input
rlabel metal3 s 279600 60368 280000 60424 6 x_start[426]
port 1355 nsew signal input
rlabel metal3 s 279600 60480 280000 60536 6 x_start[427]
port 1356 nsew signal input
rlabel metal3 s 279600 60592 280000 60648 6 x_start[428]
port 1357 nsew signal input
rlabel metal3 s 279600 60704 280000 60760 6 x_start[429]
port 1358 nsew signal input
rlabel metal3 s 279600 17360 280000 17416 6 x_start[42]
port 1359 nsew signal input
rlabel metal3 s 279600 60816 280000 60872 6 x_start[430]
port 1360 nsew signal input
rlabel metal3 s 279600 60928 280000 60984 6 x_start[431]
port 1361 nsew signal input
rlabel metal3 s 279600 61040 280000 61096 6 x_start[432]
port 1362 nsew signal input
rlabel metal3 s 279600 61152 280000 61208 6 x_start[433]
port 1363 nsew signal input
rlabel metal3 s 279600 61264 280000 61320 6 x_start[434]
port 1364 nsew signal input
rlabel metal3 s 279600 61376 280000 61432 6 x_start[435]
port 1365 nsew signal input
rlabel metal3 s 279600 61488 280000 61544 6 x_start[436]
port 1366 nsew signal input
rlabel metal3 s 279600 61600 280000 61656 6 x_start[437]
port 1367 nsew signal input
rlabel metal3 s 279600 61712 280000 61768 6 x_start[438]
port 1368 nsew signal input
rlabel metal3 s 279600 61824 280000 61880 6 x_start[439]
port 1369 nsew signal input
rlabel metal3 s 279600 17472 280000 17528 6 x_start[43]
port 1370 nsew signal input
rlabel metal3 s 279600 61936 280000 61992 6 x_start[440]
port 1371 nsew signal input
rlabel metal3 s 279600 62048 280000 62104 6 x_start[441]
port 1372 nsew signal input
rlabel metal3 s 279600 62160 280000 62216 6 x_start[442]
port 1373 nsew signal input
rlabel metal3 s 279600 62272 280000 62328 6 x_start[443]
port 1374 nsew signal input
rlabel metal3 s 279600 62384 280000 62440 6 x_start[444]
port 1375 nsew signal input
rlabel metal3 s 279600 62496 280000 62552 6 x_start[445]
port 1376 nsew signal input
rlabel metal3 s 279600 62608 280000 62664 6 x_start[446]
port 1377 nsew signal input
rlabel metal3 s 279600 62720 280000 62776 6 x_start[447]
port 1378 nsew signal input
rlabel metal3 s 279600 62832 280000 62888 6 x_start[448]
port 1379 nsew signal input
rlabel metal3 s 279600 62944 280000 63000 6 x_start[449]
port 1380 nsew signal input
rlabel metal3 s 279600 17584 280000 17640 6 x_start[44]
port 1381 nsew signal input
rlabel metal3 s 279600 63056 280000 63112 6 x_start[450]
port 1382 nsew signal input
rlabel metal3 s 279600 63168 280000 63224 6 x_start[451]
port 1383 nsew signal input
rlabel metal3 s 279600 63280 280000 63336 6 x_start[452]
port 1384 nsew signal input
rlabel metal3 s 279600 63392 280000 63448 6 x_start[453]
port 1385 nsew signal input
rlabel metal3 s 279600 63504 280000 63560 6 x_start[454]
port 1386 nsew signal input
rlabel metal3 s 279600 63616 280000 63672 6 x_start[455]
port 1387 nsew signal input
rlabel metal3 s 279600 63728 280000 63784 6 x_start[456]
port 1388 nsew signal input
rlabel metal3 s 279600 63840 280000 63896 6 x_start[457]
port 1389 nsew signal input
rlabel metal3 s 279600 63952 280000 64008 6 x_start[458]
port 1390 nsew signal input
rlabel metal3 s 279600 64064 280000 64120 6 x_start[459]
port 1391 nsew signal input
rlabel metal3 s 279600 17696 280000 17752 6 x_start[45]
port 1392 nsew signal input
rlabel metal3 s 279600 64176 280000 64232 6 x_start[460]
port 1393 nsew signal input
rlabel metal3 s 279600 64288 280000 64344 6 x_start[461]
port 1394 nsew signal input
rlabel metal3 s 279600 64400 280000 64456 6 x_start[462]
port 1395 nsew signal input
rlabel metal3 s 279600 64512 280000 64568 6 x_start[463]
port 1396 nsew signal input
rlabel metal3 s 279600 64624 280000 64680 6 x_start[464]
port 1397 nsew signal input
rlabel metal3 s 279600 64736 280000 64792 6 x_start[465]
port 1398 nsew signal input
rlabel metal3 s 279600 64848 280000 64904 6 x_start[466]
port 1399 nsew signal input
rlabel metal3 s 279600 64960 280000 65016 6 x_start[467]
port 1400 nsew signal input
rlabel metal3 s 279600 65072 280000 65128 6 x_start[468]
port 1401 nsew signal input
rlabel metal3 s 279600 65184 280000 65240 6 x_start[469]
port 1402 nsew signal input
rlabel metal3 s 279600 17808 280000 17864 6 x_start[46]
port 1403 nsew signal input
rlabel metal3 s 279600 65296 280000 65352 6 x_start[470]
port 1404 nsew signal input
rlabel metal3 s 279600 65408 280000 65464 6 x_start[471]
port 1405 nsew signal input
rlabel metal3 s 279600 65520 280000 65576 6 x_start[472]
port 1406 nsew signal input
rlabel metal3 s 279600 65632 280000 65688 6 x_start[473]
port 1407 nsew signal input
rlabel metal3 s 279600 65744 280000 65800 6 x_start[474]
port 1408 nsew signal input
rlabel metal3 s 279600 65856 280000 65912 6 x_start[475]
port 1409 nsew signal input
rlabel metal3 s 279600 65968 280000 66024 6 x_start[476]
port 1410 nsew signal input
rlabel metal3 s 279600 66080 280000 66136 6 x_start[477]
port 1411 nsew signal input
rlabel metal3 s 279600 66192 280000 66248 6 x_start[478]
port 1412 nsew signal input
rlabel metal3 s 279600 66304 280000 66360 6 x_start[479]
port 1413 nsew signal input
rlabel metal3 s 279600 17920 280000 17976 6 x_start[47]
port 1414 nsew signal input
rlabel metal3 s 279600 66416 280000 66472 6 x_start[480]
port 1415 nsew signal input
rlabel metal3 s 279600 66528 280000 66584 6 x_start[481]
port 1416 nsew signal input
rlabel metal3 s 279600 66640 280000 66696 6 x_start[482]
port 1417 nsew signal input
rlabel metal3 s 279600 66752 280000 66808 6 x_start[483]
port 1418 nsew signal input
rlabel metal3 s 279600 66864 280000 66920 6 x_start[484]
port 1419 nsew signal input
rlabel metal3 s 279600 66976 280000 67032 6 x_start[485]
port 1420 nsew signal input
rlabel metal3 s 279600 67088 280000 67144 6 x_start[486]
port 1421 nsew signal input
rlabel metal3 s 279600 67200 280000 67256 6 x_start[487]
port 1422 nsew signal input
rlabel metal3 s 279600 67312 280000 67368 6 x_start[488]
port 1423 nsew signal input
rlabel metal3 s 279600 67424 280000 67480 6 x_start[489]
port 1424 nsew signal input
rlabel metal3 s 279600 18032 280000 18088 6 x_start[48]
port 1425 nsew signal input
rlabel metal3 s 279600 67536 280000 67592 6 x_start[490]
port 1426 nsew signal input
rlabel metal3 s 279600 67648 280000 67704 6 x_start[491]
port 1427 nsew signal input
rlabel metal3 s 279600 67760 280000 67816 6 x_start[492]
port 1428 nsew signal input
rlabel metal3 s 279600 67872 280000 67928 6 x_start[493]
port 1429 nsew signal input
rlabel metal3 s 279600 67984 280000 68040 6 x_start[494]
port 1430 nsew signal input
rlabel metal3 s 279600 68096 280000 68152 6 x_start[495]
port 1431 nsew signal input
rlabel metal3 s 279600 68208 280000 68264 6 x_start[496]
port 1432 nsew signal input
rlabel metal3 s 279600 68320 280000 68376 6 x_start[497]
port 1433 nsew signal input
rlabel metal3 s 279600 68432 280000 68488 6 x_start[498]
port 1434 nsew signal input
rlabel metal3 s 279600 68544 280000 68600 6 x_start[499]
port 1435 nsew signal input
rlabel metal3 s 279600 18144 280000 18200 6 x_start[49]
port 1436 nsew signal input
rlabel metal3 s 279600 13104 280000 13160 6 x_start[4]
port 1437 nsew signal input
rlabel metal3 s 279600 68656 280000 68712 6 x_start[500]
port 1438 nsew signal input
rlabel metal3 s 279600 68768 280000 68824 6 x_start[501]
port 1439 nsew signal input
rlabel metal3 s 279600 68880 280000 68936 6 x_start[502]
port 1440 nsew signal input
rlabel metal3 s 279600 68992 280000 69048 6 x_start[503]
port 1441 nsew signal input
rlabel metal3 s 279600 69104 280000 69160 6 x_start[504]
port 1442 nsew signal input
rlabel metal3 s 279600 69216 280000 69272 6 x_start[505]
port 1443 nsew signal input
rlabel metal3 s 279600 69328 280000 69384 6 x_start[506]
port 1444 nsew signal input
rlabel metal3 s 279600 69440 280000 69496 6 x_start[507]
port 1445 nsew signal input
rlabel metal3 s 279600 69552 280000 69608 6 x_start[508]
port 1446 nsew signal input
rlabel metal3 s 279600 69664 280000 69720 6 x_start[509]
port 1447 nsew signal input
rlabel metal3 s 279600 18256 280000 18312 6 x_start[50]
port 1448 nsew signal input
rlabel metal3 s 279600 69776 280000 69832 6 x_start[510]
port 1449 nsew signal input
rlabel metal3 s 279600 69888 280000 69944 6 x_start[511]
port 1450 nsew signal input
rlabel metal3 s 279600 18368 280000 18424 6 x_start[51]
port 1451 nsew signal input
rlabel metal3 s 279600 18480 280000 18536 6 x_start[52]
port 1452 nsew signal input
rlabel metal3 s 279600 18592 280000 18648 6 x_start[53]
port 1453 nsew signal input
rlabel metal3 s 279600 18704 280000 18760 6 x_start[54]
port 1454 nsew signal input
rlabel metal3 s 279600 18816 280000 18872 6 x_start[55]
port 1455 nsew signal input
rlabel metal3 s 279600 18928 280000 18984 6 x_start[56]
port 1456 nsew signal input
rlabel metal3 s 279600 19040 280000 19096 6 x_start[57]
port 1457 nsew signal input
rlabel metal3 s 279600 19152 280000 19208 6 x_start[58]
port 1458 nsew signal input
rlabel metal3 s 279600 19264 280000 19320 6 x_start[59]
port 1459 nsew signal input
rlabel metal3 s 279600 13216 280000 13272 6 x_start[5]
port 1460 nsew signal input
rlabel metal3 s 279600 19376 280000 19432 6 x_start[60]
port 1461 nsew signal input
rlabel metal3 s 279600 19488 280000 19544 6 x_start[61]
port 1462 nsew signal input
rlabel metal3 s 279600 19600 280000 19656 6 x_start[62]
port 1463 nsew signal input
rlabel metal3 s 279600 19712 280000 19768 6 x_start[63]
port 1464 nsew signal input
rlabel metal3 s 279600 19824 280000 19880 6 x_start[64]
port 1465 nsew signal input
rlabel metal3 s 279600 19936 280000 19992 6 x_start[65]
port 1466 nsew signal input
rlabel metal3 s 279600 20048 280000 20104 6 x_start[66]
port 1467 nsew signal input
rlabel metal3 s 279600 20160 280000 20216 6 x_start[67]
port 1468 nsew signal input
rlabel metal3 s 279600 20272 280000 20328 6 x_start[68]
port 1469 nsew signal input
rlabel metal3 s 279600 20384 280000 20440 6 x_start[69]
port 1470 nsew signal input
rlabel metal3 s 279600 13328 280000 13384 6 x_start[6]
port 1471 nsew signal input
rlabel metal3 s 279600 20496 280000 20552 6 x_start[70]
port 1472 nsew signal input
rlabel metal3 s 279600 20608 280000 20664 6 x_start[71]
port 1473 nsew signal input
rlabel metal3 s 279600 20720 280000 20776 6 x_start[72]
port 1474 nsew signal input
rlabel metal3 s 279600 20832 280000 20888 6 x_start[73]
port 1475 nsew signal input
rlabel metal3 s 279600 20944 280000 21000 6 x_start[74]
port 1476 nsew signal input
rlabel metal3 s 279600 21056 280000 21112 6 x_start[75]
port 1477 nsew signal input
rlabel metal3 s 279600 21168 280000 21224 6 x_start[76]
port 1478 nsew signal input
rlabel metal3 s 279600 21280 280000 21336 6 x_start[77]
port 1479 nsew signal input
rlabel metal3 s 279600 21392 280000 21448 6 x_start[78]
port 1480 nsew signal input
rlabel metal3 s 279600 21504 280000 21560 6 x_start[79]
port 1481 nsew signal input
rlabel metal3 s 279600 13440 280000 13496 6 x_start[7]
port 1482 nsew signal input
rlabel metal3 s 279600 21616 280000 21672 6 x_start[80]
port 1483 nsew signal input
rlabel metal3 s 279600 21728 280000 21784 6 x_start[81]
port 1484 nsew signal input
rlabel metal3 s 279600 21840 280000 21896 6 x_start[82]
port 1485 nsew signal input
rlabel metal3 s 279600 21952 280000 22008 6 x_start[83]
port 1486 nsew signal input
rlabel metal3 s 279600 22064 280000 22120 6 x_start[84]
port 1487 nsew signal input
rlabel metal3 s 279600 22176 280000 22232 6 x_start[85]
port 1488 nsew signal input
rlabel metal3 s 279600 22288 280000 22344 6 x_start[86]
port 1489 nsew signal input
rlabel metal3 s 279600 22400 280000 22456 6 x_start[87]
port 1490 nsew signal input
rlabel metal3 s 279600 22512 280000 22568 6 x_start[88]
port 1491 nsew signal input
rlabel metal3 s 279600 22624 280000 22680 6 x_start[89]
port 1492 nsew signal input
rlabel metal3 s 279600 13552 280000 13608 6 x_start[8]
port 1493 nsew signal input
rlabel metal3 s 279600 22736 280000 22792 6 x_start[90]
port 1494 nsew signal input
rlabel metal3 s 279600 22848 280000 22904 6 x_start[91]
port 1495 nsew signal input
rlabel metal3 s 279600 22960 280000 23016 6 x_start[92]
port 1496 nsew signal input
rlabel metal3 s 279600 23072 280000 23128 6 x_start[93]
port 1497 nsew signal input
rlabel metal3 s 279600 23184 280000 23240 6 x_start[94]
port 1498 nsew signal input
rlabel metal3 s 279600 23296 280000 23352 6 x_start[95]
port 1499 nsew signal input
rlabel metal3 s 279600 23408 280000 23464 6 x_start[96]
port 1500 nsew signal input
rlabel metal3 s 279600 23520 280000 23576 6 x_start[97]
port 1501 nsew signal input
rlabel metal3 s 279600 23632 280000 23688 6 x_start[98]
port 1502 nsew signal input
rlabel metal3 s 279600 23744 280000 23800 6 x_start[99]
port 1503 nsew signal input
rlabel metal3 s 279600 13664 280000 13720 6 x_start[9]
port 1504 nsew signal input
rlabel metal2 s 104608 0 104664 400 6 y[0]
port 1505 nsew signal input
rlabel metal2 s 138208 0 138264 400 6 y[100]
port 1506 nsew signal input
rlabel metal2 s 138544 0 138600 400 6 y[101]
port 1507 nsew signal input
rlabel metal2 s 138880 0 138936 400 6 y[102]
port 1508 nsew signal input
rlabel metal2 s 139216 0 139272 400 6 y[103]
port 1509 nsew signal input
rlabel metal2 s 139552 0 139608 400 6 y[104]
port 1510 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 y[105]
port 1511 nsew signal input
rlabel metal2 s 140224 0 140280 400 6 y[106]
port 1512 nsew signal input
rlabel metal2 s 140560 0 140616 400 6 y[107]
port 1513 nsew signal input
rlabel metal2 s 140896 0 140952 400 6 y[108]
port 1514 nsew signal input
rlabel metal2 s 141232 0 141288 400 6 y[109]
port 1515 nsew signal input
rlabel metal2 s 107968 0 108024 400 6 y[10]
port 1516 nsew signal input
rlabel metal2 s 141568 0 141624 400 6 y[110]
port 1517 nsew signal input
rlabel metal2 s 141904 0 141960 400 6 y[111]
port 1518 nsew signal input
rlabel metal2 s 142240 0 142296 400 6 y[112]
port 1519 nsew signal input
rlabel metal2 s 142576 0 142632 400 6 y[113]
port 1520 nsew signal input
rlabel metal2 s 142912 0 142968 400 6 y[114]
port 1521 nsew signal input
rlabel metal2 s 143248 0 143304 400 6 y[115]
port 1522 nsew signal input
rlabel metal2 s 143584 0 143640 400 6 y[116]
port 1523 nsew signal input
rlabel metal2 s 143920 0 143976 400 6 y[117]
port 1524 nsew signal input
rlabel metal2 s 144256 0 144312 400 6 y[118]
port 1525 nsew signal input
rlabel metal2 s 144592 0 144648 400 6 y[119]
port 1526 nsew signal input
rlabel metal2 s 108304 0 108360 400 6 y[11]
port 1527 nsew signal input
rlabel metal2 s 144928 0 144984 400 6 y[120]
port 1528 nsew signal input
rlabel metal2 s 145264 0 145320 400 6 y[121]
port 1529 nsew signal input
rlabel metal2 s 145600 0 145656 400 6 y[122]
port 1530 nsew signal input
rlabel metal2 s 145936 0 145992 400 6 y[123]
port 1531 nsew signal input
rlabel metal2 s 146272 0 146328 400 6 y[124]
port 1532 nsew signal input
rlabel metal2 s 146608 0 146664 400 6 y[125]
port 1533 nsew signal input
rlabel metal2 s 146944 0 147000 400 6 y[126]
port 1534 nsew signal input
rlabel metal2 s 147280 0 147336 400 6 y[127]
port 1535 nsew signal input
rlabel metal2 s 147616 0 147672 400 6 y[128]
port 1536 nsew signal input
rlabel metal2 s 147952 0 148008 400 6 y[129]
port 1537 nsew signal input
rlabel metal2 s 108640 0 108696 400 6 y[12]
port 1538 nsew signal input
rlabel metal2 s 148288 0 148344 400 6 y[130]
port 1539 nsew signal input
rlabel metal2 s 148624 0 148680 400 6 y[131]
port 1540 nsew signal input
rlabel metal2 s 148960 0 149016 400 6 y[132]
port 1541 nsew signal input
rlabel metal2 s 149296 0 149352 400 6 y[133]
port 1542 nsew signal input
rlabel metal2 s 149632 0 149688 400 6 y[134]
port 1543 nsew signal input
rlabel metal2 s 149968 0 150024 400 6 y[135]
port 1544 nsew signal input
rlabel metal2 s 150304 0 150360 400 6 y[136]
port 1545 nsew signal input
rlabel metal2 s 150640 0 150696 400 6 y[137]
port 1546 nsew signal input
rlabel metal2 s 150976 0 151032 400 6 y[138]
port 1547 nsew signal input
rlabel metal2 s 151312 0 151368 400 6 y[139]
port 1548 nsew signal input
rlabel metal2 s 108976 0 109032 400 6 y[13]
port 1549 nsew signal input
rlabel metal2 s 151648 0 151704 400 6 y[140]
port 1550 nsew signal input
rlabel metal2 s 151984 0 152040 400 6 y[141]
port 1551 nsew signal input
rlabel metal2 s 152320 0 152376 400 6 y[142]
port 1552 nsew signal input
rlabel metal2 s 152656 0 152712 400 6 y[143]
port 1553 nsew signal input
rlabel metal2 s 152992 0 153048 400 6 y[144]
port 1554 nsew signal input
rlabel metal2 s 153328 0 153384 400 6 y[145]
port 1555 nsew signal input
rlabel metal2 s 153664 0 153720 400 6 y[146]
port 1556 nsew signal input
rlabel metal2 s 154000 0 154056 400 6 y[147]
port 1557 nsew signal input
rlabel metal2 s 154336 0 154392 400 6 y[148]
port 1558 nsew signal input
rlabel metal2 s 154672 0 154728 400 6 y[149]
port 1559 nsew signal input
rlabel metal2 s 109312 0 109368 400 6 y[14]
port 1560 nsew signal input
rlabel metal2 s 155008 0 155064 400 6 y[150]
port 1561 nsew signal input
rlabel metal2 s 155344 0 155400 400 6 y[151]
port 1562 nsew signal input
rlabel metal2 s 155680 0 155736 400 6 y[152]
port 1563 nsew signal input
rlabel metal2 s 156016 0 156072 400 6 y[153]
port 1564 nsew signal input
rlabel metal2 s 156352 0 156408 400 6 y[154]
port 1565 nsew signal input
rlabel metal2 s 156688 0 156744 400 6 y[155]
port 1566 nsew signal input
rlabel metal2 s 157024 0 157080 400 6 y[156]
port 1567 nsew signal input
rlabel metal2 s 157360 0 157416 400 6 y[157]
port 1568 nsew signal input
rlabel metal2 s 157696 0 157752 400 6 y[158]
port 1569 nsew signal input
rlabel metal2 s 158032 0 158088 400 6 y[159]
port 1570 nsew signal input
rlabel metal2 s 109648 0 109704 400 6 y[15]
port 1571 nsew signal input
rlabel metal2 s 158368 0 158424 400 6 y[160]
port 1572 nsew signal input
rlabel metal2 s 158704 0 158760 400 6 y[161]
port 1573 nsew signal input
rlabel metal2 s 159040 0 159096 400 6 y[162]
port 1574 nsew signal input
rlabel metal2 s 159376 0 159432 400 6 y[163]
port 1575 nsew signal input
rlabel metal2 s 159712 0 159768 400 6 y[164]
port 1576 nsew signal input
rlabel metal2 s 160048 0 160104 400 6 y[165]
port 1577 nsew signal input
rlabel metal2 s 160384 0 160440 400 6 y[166]
port 1578 nsew signal input
rlabel metal2 s 160720 0 160776 400 6 y[167]
port 1579 nsew signal input
rlabel metal2 s 161056 0 161112 400 6 y[168]
port 1580 nsew signal input
rlabel metal2 s 161392 0 161448 400 6 y[169]
port 1581 nsew signal input
rlabel metal2 s 109984 0 110040 400 6 y[16]
port 1582 nsew signal input
rlabel metal2 s 161728 0 161784 400 6 y[170]
port 1583 nsew signal input
rlabel metal2 s 162064 0 162120 400 6 y[171]
port 1584 nsew signal input
rlabel metal2 s 162400 0 162456 400 6 y[172]
port 1585 nsew signal input
rlabel metal2 s 162736 0 162792 400 6 y[173]
port 1586 nsew signal input
rlabel metal2 s 163072 0 163128 400 6 y[174]
port 1587 nsew signal input
rlabel metal2 s 163408 0 163464 400 6 y[175]
port 1588 nsew signal input
rlabel metal2 s 163744 0 163800 400 6 y[176]
port 1589 nsew signal input
rlabel metal2 s 164080 0 164136 400 6 y[177]
port 1590 nsew signal input
rlabel metal2 s 164416 0 164472 400 6 y[178]
port 1591 nsew signal input
rlabel metal2 s 164752 0 164808 400 6 y[179]
port 1592 nsew signal input
rlabel metal2 s 110320 0 110376 400 6 y[17]
port 1593 nsew signal input
rlabel metal2 s 165088 0 165144 400 6 y[180]
port 1594 nsew signal input
rlabel metal2 s 165424 0 165480 400 6 y[181]
port 1595 nsew signal input
rlabel metal2 s 165760 0 165816 400 6 y[182]
port 1596 nsew signal input
rlabel metal2 s 166096 0 166152 400 6 y[183]
port 1597 nsew signal input
rlabel metal2 s 166432 0 166488 400 6 y[184]
port 1598 nsew signal input
rlabel metal2 s 166768 0 166824 400 6 y[185]
port 1599 nsew signal input
rlabel metal2 s 167104 0 167160 400 6 y[186]
port 1600 nsew signal input
rlabel metal2 s 167440 0 167496 400 6 y[187]
port 1601 nsew signal input
rlabel metal2 s 167776 0 167832 400 6 y[188]
port 1602 nsew signal input
rlabel metal2 s 168112 0 168168 400 6 y[189]
port 1603 nsew signal input
rlabel metal2 s 110656 0 110712 400 6 y[18]
port 1604 nsew signal input
rlabel metal2 s 168448 0 168504 400 6 y[190]
port 1605 nsew signal input
rlabel metal2 s 168784 0 168840 400 6 y[191]
port 1606 nsew signal input
rlabel metal2 s 169120 0 169176 400 6 y[192]
port 1607 nsew signal input
rlabel metal2 s 169456 0 169512 400 6 y[193]
port 1608 nsew signal input
rlabel metal2 s 169792 0 169848 400 6 y[194]
port 1609 nsew signal input
rlabel metal2 s 170128 0 170184 400 6 y[195]
port 1610 nsew signal input
rlabel metal2 s 170464 0 170520 400 6 y[196]
port 1611 nsew signal input
rlabel metal2 s 170800 0 170856 400 6 y[197]
port 1612 nsew signal input
rlabel metal2 s 171136 0 171192 400 6 y[198]
port 1613 nsew signal input
rlabel metal2 s 171472 0 171528 400 6 y[199]
port 1614 nsew signal input
rlabel metal2 s 110992 0 111048 400 6 y[19]
port 1615 nsew signal input
rlabel metal2 s 104944 0 105000 400 6 y[1]
port 1616 nsew signal input
rlabel metal2 s 171808 0 171864 400 6 y[200]
port 1617 nsew signal input
rlabel metal2 s 172144 0 172200 400 6 y[201]
port 1618 nsew signal input
rlabel metal2 s 172480 0 172536 400 6 y[202]
port 1619 nsew signal input
rlabel metal2 s 172816 0 172872 400 6 y[203]
port 1620 nsew signal input
rlabel metal2 s 173152 0 173208 400 6 y[204]
port 1621 nsew signal input
rlabel metal2 s 173488 0 173544 400 6 y[205]
port 1622 nsew signal input
rlabel metal2 s 173824 0 173880 400 6 y[206]
port 1623 nsew signal input
rlabel metal2 s 174160 0 174216 400 6 y[207]
port 1624 nsew signal input
rlabel metal2 s 174496 0 174552 400 6 y[208]
port 1625 nsew signal input
rlabel metal2 s 174832 0 174888 400 6 y[209]
port 1626 nsew signal input
rlabel metal2 s 111328 0 111384 400 6 y[20]
port 1627 nsew signal input
rlabel metal2 s 175168 0 175224 400 6 y[210]
port 1628 nsew signal input
rlabel metal2 s 175504 0 175560 400 6 y[211]
port 1629 nsew signal input
rlabel metal2 s 175840 0 175896 400 6 y[212]
port 1630 nsew signal input
rlabel metal2 s 176176 0 176232 400 6 y[213]
port 1631 nsew signal input
rlabel metal2 s 176512 0 176568 400 6 y[214]
port 1632 nsew signal input
rlabel metal2 s 176848 0 176904 400 6 y[215]
port 1633 nsew signal input
rlabel metal2 s 177184 0 177240 400 6 y[216]
port 1634 nsew signal input
rlabel metal2 s 177520 0 177576 400 6 y[217]
port 1635 nsew signal input
rlabel metal2 s 177856 0 177912 400 6 y[218]
port 1636 nsew signal input
rlabel metal2 s 178192 0 178248 400 6 y[219]
port 1637 nsew signal input
rlabel metal2 s 111664 0 111720 400 6 y[21]
port 1638 nsew signal input
rlabel metal2 s 178528 0 178584 400 6 y[220]
port 1639 nsew signal input
rlabel metal2 s 178864 0 178920 400 6 y[221]
port 1640 nsew signal input
rlabel metal2 s 179200 0 179256 400 6 y[222]
port 1641 nsew signal input
rlabel metal2 s 179536 0 179592 400 6 y[223]
port 1642 nsew signal input
rlabel metal2 s 179872 0 179928 400 6 y[224]
port 1643 nsew signal input
rlabel metal2 s 180208 0 180264 400 6 y[225]
port 1644 nsew signal input
rlabel metal2 s 180544 0 180600 400 6 y[226]
port 1645 nsew signal input
rlabel metal2 s 180880 0 180936 400 6 y[227]
port 1646 nsew signal input
rlabel metal2 s 181216 0 181272 400 6 y[228]
port 1647 nsew signal input
rlabel metal2 s 181552 0 181608 400 6 y[229]
port 1648 nsew signal input
rlabel metal2 s 112000 0 112056 400 6 y[22]
port 1649 nsew signal input
rlabel metal2 s 181888 0 181944 400 6 y[230]
port 1650 nsew signal input
rlabel metal2 s 182224 0 182280 400 6 y[231]
port 1651 nsew signal input
rlabel metal2 s 182560 0 182616 400 6 y[232]
port 1652 nsew signal input
rlabel metal2 s 182896 0 182952 400 6 y[233]
port 1653 nsew signal input
rlabel metal2 s 183232 0 183288 400 6 y[234]
port 1654 nsew signal input
rlabel metal2 s 183568 0 183624 400 6 y[235]
port 1655 nsew signal input
rlabel metal2 s 183904 0 183960 400 6 y[236]
port 1656 nsew signal input
rlabel metal2 s 184240 0 184296 400 6 y[237]
port 1657 nsew signal input
rlabel metal2 s 184576 0 184632 400 6 y[238]
port 1658 nsew signal input
rlabel metal2 s 184912 0 184968 400 6 y[239]
port 1659 nsew signal input
rlabel metal2 s 112336 0 112392 400 6 y[23]
port 1660 nsew signal input
rlabel metal2 s 185248 0 185304 400 6 y[240]
port 1661 nsew signal input
rlabel metal2 s 185584 0 185640 400 6 y[241]
port 1662 nsew signal input
rlabel metal2 s 185920 0 185976 400 6 y[242]
port 1663 nsew signal input
rlabel metal2 s 186256 0 186312 400 6 y[243]
port 1664 nsew signal input
rlabel metal2 s 186592 0 186648 400 6 y[244]
port 1665 nsew signal input
rlabel metal2 s 186928 0 186984 400 6 y[245]
port 1666 nsew signal input
rlabel metal2 s 187264 0 187320 400 6 y[246]
port 1667 nsew signal input
rlabel metal2 s 187600 0 187656 400 6 y[247]
port 1668 nsew signal input
rlabel metal2 s 187936 0 187992 400 6 y[248]
port 1669 nsew signal input
rlabel metal2 s 188272 0 188328 400 6 y[249]
port 1670 nsew signal input
rlabel metal2 s 112672 0 112728 400 6 y[24]
port 1671 nsew signal input
rlabel metal2 s 188608 0 188664 400 6 y[250]
port 1672 nsew signal input
rlabel metal2 s 188944 0 189000 400 6 y[251]
port 1673 nsew signal input
rlabel metal2 s 189280 0 189336 400 6 y[252]
port 1674 nsew signal input
rlabel metal2 s 189616 0 189672 400 6 y[253]
port 1675 nsew signal input
rlabel metal2 s 189952 0 190008 400 6 y[254]
port 1676 nsew signal input
rlabel metal2 s 190288 0 190344 400 6 y[255]
port 1677 nsew signal input
rlabel metal2 s 190624 0 190680 400 6 y[256]
port 1678 nsew signal input
rlabel metal2 s 190960 0 191016 400 6 y[257]
port 1679 nsew signal input
rlabel metal2 s 191296 0 191352 400 6 y[258]
port 1680 nsew signal input
rlabel metal2 s 191632 0 191688 400 6 y[259]
port 1681 nsew signal input
rlabel metal2 s 113008 0 113064 400 6 y[25]
port 1682 nsew signal input
rlabel metal2 s 191968 0 192024 400 6 y[260]
port 1683 nsew signal input
rlabel metal2 s 192304 0 192360 400 6 y[261]
port 1684 nsew signal input
rlabel metal2 s 192640 0 192696 400 6 y[262]
port 1685 nsew signal input
rlabel metal2 s 192976 0 193032 400 6 y[263]
port 1686 nsew signal input
rlabel metal2 s 193312 0 193368 400 6 y[264]
port 1687 nsew signal input
rlabel metal2 s 193648 0 193704 400 6 y[265]
port 1688 nsew signal input
rlabel metal2 s 193984 0 194040 400 6 y[266]
port 1689 nsew signal input
rlabel metal2 s 194320 0 194376 400 6 y[267]
port 1690 nsew signal input
rlabel metal2 s 194656 0 194712 400 6 y[268]
port 1691 nsew signal input
rlabel metal2 s 194992 0 195048 400 6 y[269]
port 1692 nsew signal input
rlabel metal2 s 113344 0 113400 400 6 y[26]
port 1693 nsew signal input
rlabel metal2 s 195328 0 195384 400 6 y[270]
port 1694 nsew signal input
rlabel metal2 s 195664 0 195720 400 6 y[271]
port 1695 nsew signal input
rlabel metal2 s 196000 0 196056 400 6 y[272]
port 1696 nsew signal input
rlabel metal2 s 196336 0 196392 400 6 y[273]
port 1697 nsew signal input
rlabel metal2 s 196672 0 196728 400 6 y[274]
port 1698 nsew signal input
rlabel metal2 s 197008 0 197064 400 6 y[275]
port 1699 nsew signal input
rlabel metal2 s 197344 0 197400 400 6 y[276]
port 1700 nsew signal input
rlabel metal2 s 197680 0 197736 400 6 y[277]
port 1701 nsew signal input
rlabel metal2 s 198016 0 198072 400 6 y[278]
port 1702 nsew signal input
rlabel metal2 s 198352 0 198408 400 6 y[279]
port 1703 nsew signal input
rlabel metal2 s 113680 0 113736 400 6 y[27]
port 1704 nsew signal input
rlabel metal2 s 198688 0 198744 400 6 y[280]
port 1705 nsew signal input
rlabel metal2 s 199024 0 199080 400 6 y[281]
port 1706 nsew signal input
rlabel metal2 s 199360 0 199416 400 6 y[282]
port 1707 nsew signal input
rlabel metal2 s 199696 0 199752 400 6 y[283]
port 1708 nsew signal input
rlabel metal2 s 200032 0 200088 400 6 y[284]
port 1709 nsew signal input
rlabel metal2 s 200368 0 200424 400 6 y[285]
port 1710 nsew signal input
rlabel metal2 s 200704 0 200760 400 6 y[286]
port 1711 nsew signal input
rlabel metal2 s 201040 0 201096 400 6 y[287]
port 1712 nsew signal input
rlabel metal2 s 201376 0 201432 400 6 y[288]
port 1713 nsew signal input
rlabel metal2 s 201712 0 201768 400 6 y[289]
port 1714 nsew signal input
rlabel metal2 s 114016 0 114072 400 6 y[28]
port 1715 nsew signal input
rlabel metal2 s 202048 0 202104 400 6 y[290]
port 1716 nsew signal input
rlabel metal2 s 202384 0 202440 400 6 y[291]
port 1717 nsew signal input
rlabel metal2 s 202720 0 202776 400 6 y[292]
port 1718 nsew signal input
rlabel metal2 s 203056 0 203112 400 6 y[293]
port 1719 nsew signal input
rlabel metal2 s 203392 0 203448 400 6 y[294]
port 1720 nsew signal input
rlabel metal2 s 203728 0 203784 400 6 y[295]
port 1721 nsew signal input
rlabel metal2 s 204064 0 204120 400 6 y[296]
port 1722 nsew signal input
rlabel metal2 s 204400 0 204456 400 6 y[297]
port 1723 nsew signal input
rlabel metal2 s 204736 0 204792 400 6 y[298]
port 1724 nsew signal input
rlabel metal2 s 205072 0 205128 400 6 y[299]
port 1725 nsew signal input
rlabel metal2 s 114352 0 114408 400 6 y[29]
port 1726 nsew signal input
rlabel metal2 s 105280 0 105336 400 6 y[2]
port 1727 nsew signal input
rlabel metal2 s 205408 0 205464 400 6 y[300]
port 1728 nsew signal input
rlabel metal2 s 205744 0 205800 400 6 y[301]
port 1729 nsew signal input
rlabel metal2 s 206080 0 206136 400 6 y[302]
port 1730 nsew signal input
rlabel metal2 s 206416 0 206472 400 6 y[303]
port 1731 nsew signal input
rlabel metal2 s 206752 0 206808 400 6 y[304]
port 1732 nsew signal input
rlabel metal2 s 207088 0 207144 400 6 y[305]
port 1733 nsew signal input
rlabel metal2 s 207424 0 207480 400 6 y[306]
port 1734 nsew signal input
rlabel metal2 s 207760 0 207816 400 6 y[307]
port 1735 nsew signal input
rlabel metal2 s 208096 0 208152 400 6 y[308]
port 1736 nsew signal input
rlabel metal2 s 208432 0 208488 400 6 y[309]
port 1737 nsew signal input
rlabel metal2 s 114688 0 114744 400 6 y[30]
port 1738 nsew signal input
rlabel metal2 s 208768 0 208824 400 6 y[310]
port 1739 nsew signal input
rlabel metal2 s 209104 0 209160 400 6 y[311]
port 1740 nsew signal input
rlabel metal2 s 209440 0 209496 400 6 y[312]
port 1741 nsew signal input
rlabel metal2 s 209776 0 209832 400 6 y[313]
port 1742 nsew signal input
rlabel metal2 s 210112 0 210168 400 6 y[314]
port 1743 nsew signal input
rlabel metal2 s 210448 0 210504 400 6 y[315]
port 1744 nsew signal input
rlabel metal2 s 210784 0 210840 400 6 y[316]
port 1745 nsew signal input
rlabel metal2 s 211120 0 211176 400 6 y[317]
port 1746 nsew signal input
rlabel metal2 s 211456 0 211512 400 6 y[318]
port 1747 nsew signal input
rlabel metal2 s 211792 0 211848 400 6 y[319]
port 1748 nsew signal input
rlabel metal2 s 115024 0 115080 400 6 y[31]
port 1749 nsew signal input
rlabel metal2 s 212128 0 212184 400 6 y[320]
port 1750 nsew signal input
rlabel metal2 s 212464 0 212520 400 6 y[321]
port 1751 nsew signal input
rlabel metal2 s 212800 0 212856 400 6 y[322]
port 1752 nsew signal input
rlabel metal2 s 213136 0 213192 400 6 y[323]
port 1753 nsew signal input
rlabel metal2 s 213472 0 213528 400 6 y[324]
port 1754 nsew signal input
rlabel metal2 s 213808 0 213864 400 6 y[325]
port 1755 nsew signal input
rlabel metal2 s 214144 0 214200 400 6 y[326]
port 1756 nsew signal input
rlabel metal2 s 214480 0 214536 400 6 y[327]
port 1757 nsew signal input
rlabel metal2 s 214816 0 214872 400 6 y[328]
port 1758 nsew signal input
rlabel metal2 s 215152 0 215208 400 6 y[329]
port 1759 nsew signal input
rlabel metal2 s 115360 0 115416 400 6 y[32]
port 1760 nsew signal input
rlabel metal2 s 215488 0 215544 400 6 y[330]
port 1761 nsew signal input
rlabel metal2 s 215824 0 215880 400 6 y[331]
port 1762 nsew signal input
rlabel metal2 s 216160 0 216216 400 6 y[332]
port 1763 nsew signal input
rlabel metal2 s 216496 0 216552 400 6 y[333]
port 1764 nsew signal input
rlabel metal2 s 216832 0 216888 400 6 y[334]
port 1765 nsew signal input
rlabel metal2 s 217168 0 217224 400 6 y[335]
port 1766 nsew signal input
rlabel metal2 s 217504 0 217560 400 6 y[336]
port 1767 nsew signal input
rlabel metal2 s 217840 0 217896 400 6 y[337]
port 1768 nsew signal input
rlabel metal2 s 218176 0 218232 400 6 y[338]
port 1769 nsew signal input
rlabel metal2 s 218512 0 218568 400 6 y[339]
port 1770 nsew signal input
rlabel metal2 s 115696 0 115752 400 6 y[33]
port 1771 nsew signal input
rlabel metal2 s 218848 0 218904 400 6 y[340]
port 1772 nsew signal input
rlabel metal2 s 219184 0 219240 400 6 y[341]
port 1773 nsew signal input
rlabel metal2 s 219520 0 219576 400 6 y[342]
port 1774 nsew signal input
rlabel metal2 s 219856 0 219912 400 6 y[343]
port 1775 nsew signal input
rlabel metal2 s 220192 0 220248 400 6 y[344]
port 1776 nsew signal input
rlabel metal2 s 220528 0 220584 400 6 y[345]
port 1777 nsew signal input
rlabel metal2 s 220864 0 220920 400 6 y[346]
port 1778 nsew signal input
rlabel metal2 s 221200 0 221256 400 6 y[347]
port 1779 nsew signal input
rlabel metal2 s 221536 0 221592 400 6 y[348]
port 1780 nsew signal input
rlabel metal2 s 221872 0 221928 400 6 y[349]
port 1781 nsew signal input
rlabel metal2 s 116032 0 116088 400 6 y[34]
port 1782 nsew signal input
rlabel metal2 s 222208 0 222264 400 6 y[350]
port 1783 nsew signal input
rlabel metal2 s 222544 0 222600 400 6 y[351]
port 1784 nsew signal input
rlabel metal2 s 222880 0 222936 400 6 y[352]
port 1785 nsew signal input
rlabel metal2 s 223216 0 223272 400 6 y[353]
port 1786 nsew signal input
rlabel metal2 s 223552 0 223608 400 6 y[354]
port 1787 nsew signal input
rlabel metal2 s 223888 0 223944 400 6 y[355]
port 1788 nsew signal input
rlabel metal2 s 224224 0 224280 400 6 y[356]
port 1789 nsew signal input
rlabel metal2 s 224560 0 224616 400 6 y[357]
port 1790 nsew signal input
rlabel metal2 s 224896 0 224952 400 6 y[358]
port 1791 nsew signal input
rlabel metal2 s 225232 0 225288 400 6 y[359]
port 1792 nsew signal input
rlabel metal2 s 116368 0 116424 400 6 y[35]
port 1793 nsew signal input
rlabel metal2 s 225568 0 225624 400 6 y[360]
port 1794 nsew signal input
rlabel metal2 s 225904 0 225960 400 6 y[361]
port 1795 nsew signal input
rlabel metal2 s 226240 0 226296 400 6 y[362]
port 1796 nsew signal input
rlabel metal2 s 226576 0 226632 400 6 y[363]
port 1797 nsew signal input
rlabel metal2 s 226912 0 226968 400 6 y[364]
port 1798 nsew signal input
rlabel metal2 s 227248 0 227304 400 6 y[365]
port 1799 nsew signal input
rlabel metal2 s 227584 0 227640 400 6 y[366]
port 1800 nsew signal input
rlabel metal2 s 227920 0 227976 400 6 y[367]
port 1801 nsew signal input
rlabel metal2 s 228256 0 228312 400 6 y[368]
port 1802 nsew signal input
rlabel metal2 s 228592 0 228648 400 6 y[369]
port 1803 nsew signal input
rlabel metal2 s 116704 0 116760 400 6 y[36]
port 1804 nsew signal input
rlabel metal2 s 228928 0 228984 400 6 y[370]
port 1805 nsew signal input
rlabel metal2 s 229264 0 229320 400 6 y[371]
port 1806 nsew signal input
rlabel metal2 s 229600 0 229656 400 6 y[372]
port 1807 nsew signal input
rlabel metal2 s 229936 0 229992 400 6 y[373]
port 1808 nsew signal input
rlabel metal2 s 230272 0 230328 400 6 y[374]
port 1809 nsew signal input
rlabel metal2 s 230608 0 230664 400 6 y[375]
port 1810 nsew signal input
rlabel metal2 s 230944 0 231000 400 6 y[376]
port 1811 nsew signal input
rlabel metal2 s 231280 0 231336 400 6 y[377]
port 1812 nsew signal input
rlabel metal2 s 231616 0 231672 400 6 y[378]
port 1813 nsew signal input
rlabel metal2 s 231952 0 232008 400 6 y[379]
port 1814 nsew signal input
rlabel metal2 s 117040 0 117096 400 6 y[37]
port 1815 nsew signal input
rlabel metal2 s 232288 0 232344 400 6 y[380]
port 1816 nsew signal input
rlabel metal2 s 232624 0 232680 400 6 y[381]
port 1817 nsew signal input
rlabel metal2 s 232960 0 233016 400 6 y[382]
port 1818 nsew signal input
rlabel metal2 s 233296 0 233352 400 6 y[383]
port 1819 nsew signal input
rlabel metal2 s 233632 0 233688 400 6 y[384]
port 1820 nsew signal input
rlabel metal2 s 233968 0 234024 400 6 y[385]
port 1821 nsew signal input
rlabel metal2 s 234304 0 234360 400 6 y[386]
port 1822 nsew signal input
rlabel metal2 s 234640 0 234696 400 6 y[387]
port 1823 nsew signal input
rlabel metal2 s 234976 0 235032 400 6 y[388]
port 1824 nsew signal input
rlabel metal2 s 235312 0 235368 400 6 y[389]
port 1825 nsew signal input
rlabel metal2 s 117376 0 117432 400 6 y[38]
port 1826 nsew signal input
rlabel metal2 s 235648 0 235704 400 6 y[390]
port 1827 nsew signal input
rlabel metal2 s 235984 0 236040 400 6 y[391]
port 1828 nsew signal input
rlabel metal2 s 236320 0 236376 400 6 y[392]
port 1829 nsew signal input
rlabel metal2 s 236656 0 236712 400 6 y[393]
port 1830 nsew signal input
rlabel metal2 s 236992 0 237048 400 6 y[394]
port 1831 nsew signal input
rlabel metal2 s 237328 0 237384 400 6 y[395]
port 1832 nsew signal input
rlabel metal2 s 237664 0 237720 400 6 y[396]
port 1833 nsew signal input
rlabel metal2 s 238000 0 238056 400 6 y[397]
port 1834 nsew signal input
rlabel metal2 s 238336 0 238392 400 6 y[398]
port 1835 nsew signal input
rlabel metal2 s 238672 0 238728 400 6 y[399]
port 1836 nsew signal input
rlabel metal2 s 117712 0 117768 400 6 y[39]
port 1837 nsew signal input
rlabel metal2 s 105616 0 105672 400 6 y[3]
port 1838 nsew signal input
rlabel metal2 s 239008 0 239064 400 6 y[400]
port 1839 nsew signal input
rlabel metal2 s 239344 0 239400 400 6 y[401]
port 1840 nsew signal input
rlabel metal2 s 239680 0 239736 400 6 y[402]
port 1841 nsew signal input
rlabel metal2 s 240016 0 240072 400 6 y[403]
port 1842 nsew signal input
rlabel metal2 s 240352 0 240408 400 6 y[404]
port 1843 nsew signal input
rlabel metal2 s 240688 0 240744 400 6 y[405]
port 1844 nsew signal input
rlabel metal2 s 241024 0 241080 400 6 y[406]
port 1845 nsew signal input
rlabel metal2 s 241360 0 241416 400 6 y[407]
port 1846 nsew signal input
rlabel metal2 s 241696 0 241752 400 6 y[408]
port 1847 nsew signal input
rlabel metal2 s 242032 0 242088 400 6 y[409]
port 1848 nsew signal input
rlabel metal2 s 118048 0 118104 400 6 y[40]
port 1849 nsew signal input
rlabel metal2 s 242368 0 242424 400 6 y[410]
port 1850 nsew signal input
rlabel metal2 s 242704 0 242760 400 6 y[411]
port 1851 nsew signal input
rlabel metal2 s 243040 0 243096 400 6 y[412]
port 1852 nsew signal input
rlabel metal2 s 243376 0 243432 400 6 y[413]
port 1853 nsew signal input
rlabel metal2 s 243712 0 243768 400 6 y[414]
port 1854 nsew signal input
rlabel metal2 s 244048 0 244104 400 6 y[415]
port 1855 nsew signal input
rlabel metal2 s 244384 0 244440 400 6 y[416]
port 1856 nsew signal input
rlabel metal2 s 244720 0 244776 400 6 y[417]
port 1857 nsew signal input
rlabel metal2 s 245056 0 245112 400 6 y[418]
port 1858 nsew signal input
rlabel metal2 s 245392 0 245448 400 6 y[419]
port 1859 nsew signal input
rlabel metal2 s 118384 0 118440 400 6 y[41]
port 1860 nsew signal input
rlabel metal2 s 245728 0 245784 400 6 y[420]
port 1861 nsew signal input
rlabel metal2 s 246064 0 246120 400 6 y[421]
port 1862 nsew signal input
rlabel metal2 s 246400 0 246456 400 6 y[422]
port 1863 nsew signal input
rlabel metal2 s 246736 0 246792 400 6 y[423]
port 1864 nsew signal input
rlabel metal2 s 247072 0 247128 400 6 y[424]
port 1865 nsew signal input
rlabel metal2 s 247408 0 247464 400 6 y[425]
port 1866 nsew signal input
rlabel metal2 s 247744 0 247800 400 6 y[426]
port 1867 nsew signal input
rlabel metal2 s 248080 0 248136 400 6 y[427]
port 1868 nsew signal input
rlabel metal2 s 248416 0 248472 400 6 y[428]
port 1869 nsew signal input
rlabel metal2 s 248752 0 248808 400 6 y[429]
port 1870 nsew signal input
rlabel metal2 s 118720 0 118776 400 6 y[42]
port 1871 nsew signal input
rlabel metal2 s 249088 0 249144 400 6 y[430]
port 1872 nsew signal input
rlabel metal2 s 249424 0 249480 400 6 y[431]
port 1873 nsew signal input
rlabel metal2 s 249760 0 249816 400 6 y[432]
port 1874 nsew signal input
rlabel metal2 s 250096 0 250152 400 6 y[433]
port 1875 nsew signal input
rlabel metal2 s 250432 0 250488 400 6 y[434]
port 1876 nsew signal input
rlabel metal2 s 250768 0 250824 400 6 y[435]
port 1877 nsew signal input
rlabel metal2 s 251104 0 251160 400 6 y[436]
port 1878 nsew signal input
rlabel metal2 s 251440 0 251496 400 6 y[437]
port 1879 nsew signal input
rlabel metal2 s 251776 0 251832 400 6 y[438]
port 1880 nsew signal input
rlabel metal2 s 252112 0 252168 400 6 y[439]
port 1881 nsew signal input
rlabel metal2 s 119056 0 119112 400 6 y[43]
port 1882 nsew signal input
rlabel metal2 s 252448 0 252504 400 6 y[440]
port 1883 nsew signal input
rlabel metal2 s 252784 0 252840 400 6 y[441]
port 1884 nsew signal input
rlabel metal2 s 253120 0 253176 400 6 y[442]
port 1885 nsew signal input
rlabel metal2 s 253456 0 253512 400 6 y[443]
port 1886 nsew signal input
rlabel metal2 s 253792 0 253848 400 6 y[444]
port 1887 nsew signal input
rlabel metal2 s 254128 0 254184 400 6 y[445]
port 1888 nsew signal input
rlabel metal2 s 254464 0 254520 400 6 y[446]
port 1889 nsew signal input
rlabel metal2 s 254800 0 254856 400 6 y[447]
port 1890 nsew signal input
rlabel metal2 s 255136 0 255192 400 6 y[448]
port 1891 nsew signal input
rlabel metal2 s 255472 0 255528 400 6 y[449]
port 1892 nsew signal input
rlabel metal2 s 119392 0 119448 400 6 y[44]
port 1893 nsew signal input
rlabel metal2 s 255808 0 255864 400 6 y[450]
port 1894 nsew signal input
rlabel metal2 s 256144 0 256200 400 6 y[451]
port 1895 nsew signal input
rlabel metal2 s 256480 0 256536 400 6 y[452]
port 1896 nsew signal input
rlabel metal2 s 256816 0 256872 400 6 y[453]
port 1897 nsew signal input
rlabel metal2 s 257152 0 257208 400 6 y[454]
port 1898 nsew signal input
rlabel metal2 s 257488 0 257544 400 6 y[455]
port 1899 nsew signal input
rlabel metal2 s 257824 0 257880 400 6 y[456]
port 1900 nsew signal input
rlabel metal2 s 258160 0 258216 400 6 y[457]
port 1901 nsew signal input
rlabel metal2 s 258496 0 258552 400 6 y[458]
port 1902 nsew signal input
rlabel metal2 s 258832 0 258888 400 6 y[459]
port 1903 nsew signal input
rlabel metal2 s 119728 0 119784 400 6 y[45]
port 1904 nsew signal input
rlabel metal2 s 259168 0 259224 400 6 y[460]
port 1905 nsew signal input
rlabel metal2 s 259504 0 259560 400 6 y[461]
port 1906 nsew signal input
rlabel metal2 s 259840 0 259896 400 6 y[462]
port 1907 nsew signal input
rlabel metal2 s 260176 0 260232 400 6 y[463]
port 1908 nsew signal input
rlabel metal2 s 260512 0 260568 400 6 y[464]
port 1909 nsew signal input
rlabel metal2 s 260848 0 260904 400 6 y[465]
port 1910 nsew signal input
rlabel metal2 s 261184 0 261240 400 6 y[466]
port 1911 nsew signal input
rlabel metal2 s 261520 0 261576 400 6 y[467]
port 1912 nsew signal input
rlabel metal2 s 261856 0 261912 400 6 y[468]
port 1913 nsew signal input
rlabel metal2 s 262192 0 262248 400 6 y[469]
port 1914 nsew signal input
rlabel metal2 s 120064 0 120120 400 6 y[46]
port 1915 nsew signal input
rlabel metal2 s 262528 0 262584 400 6 y[470]
port 1916 nsew signal input
rlabel metal2 s 262864 0 262920 400 6 y[471]
port 1917 nsew signal input
rlabel metal2 s 263200 0 263256 400 6 y[472]
port 1918 nsew signal input
rlabel metal2 s 263536 0 263592 400 6 y[473]
port 1919 nsew signal input
rlabel metal2 s 263872 0 263928 400 6 y[474]
port 1920 nsew signal input
rlabel metal2 s 264208 0 264264 400 6 y[475]
port 1921 nsew signal input
rlabel metal2 s 264544 0 264600 400 6 y[476]
port 1922 nsew signal input
rlabel metal2 s 264880 0 264936 400 6 y[477]
port 1923 nsew signal input
rlabel metal2 s 265216 0 265272 400 6 y[478]
port 1924 nsew signal input
rlabel metal2 s 265552 0 265608 400 6 y[479]
port 1925 nsew signal input
rlabel metal2 s 120400 0 120456 400 6 y[47]
port 1926 nsew signal input
rlabel metal2 s 265888 0 265944 400 6 y[480]
port 1927 nsew signal input
rlabel metal2 s 266224 0 266280 400 6 y[481]
port 1928 nsew signal input
rlabel metal2 s 266560 0 266616 400 6 y[482]
port 1929 nsew signal input
rlabel metal2 s 266896 0 266952 400 6 y[483]
port 1930 nsew signal input
rlabel metal2 s 267232 0 267288 400 6 y[484]
port 1931 nsew signal input
rlabel metal2 s 267568 0 267624 400 6 y[485]
port 1932 nsew signal input
rlabel metal2 s 267904 0 267960 400 6 y[486]
port 1933 nsew signal input
rlabel metal2 s 268240 0 268296 400 6 y[487]
port 1934 nsew signal input
rlabel metal2 s 268576 0 268632 400 6 y[488]
port 1935 nsew signal input
rlabel metal2 s 268912 0 268968 400 6 y[489]
port 1936 nsew signal input
rlabel metal2 s 120736 0 120792 400 6 y[48]
port 1937 nsew signal input
rlabel metal2 s 269248 0 269304 400 6 y[490]
port 1938 nsew signal input
rlabel metal2 s 269584 0 269640 400 6 y[491]
port 1939 nsew signal input
rlabel metal2 s 269920 0 269976 400 6 y[492]
port 1940 nsew signal input
rlabel metal2 s 270256 0 270312 400 6 y[493]
port 1941 nsew signal input
rlabel metal2 s 270592 0 270648 400 6 y[494]
port 1942 nsew signal input
rlabel metal2 s 270928 0 270984 400 6 y[495]
port 1943 nsew signal input
rlabel metal2 s 271264 0 271320 400 6 y[496]
port 1944 nsew signal input
rlabel metal2 s 271600 0 271656 400 6 y[497]
port 1945 nsew signal input
rlabel metal2 s 271936 0 271992 400 6 y[498]
port 1946 nsew signal input
rlabel metal2 s 272272 0 272328 400 6 y[499]
port 1947 nsew signal input
rlabel metal2 s 121072 0 121128 400 6 y[49]
port 1948 nsew signal input
rlabel metal2 s 105952 0 106008 400 6 y[4]
port 1949 nsew signal input
rlabel metal2 s 272608 0 272664 400 6 y[500]
port 1950 nsew signal input
rlabel metal2 s 272944 0 273000 400 6 y[501]
port 1951 nsew signal input
rlabel metal2 s 273280 0 273336 400 6 y[502]
port 1952 nsew signal input
rlabel metal2 s 273616 0 273672 400 6 y[503]
port 1953 nsew signal input
rlabel metal2 s 273952 0 274008 400 6 y[504]
port 1954 nsew signal input
rlabel metal2 s 274288 0 274344 400 6 y[505]
port 1955 nsew signal input
rlabel metal2 s 274624 0 274680 400 6 y[506]
port 1956 nsew signal input
rlabel metal2 s 274960 0 275016 400 6 y[507]
port 1957 nsew signal input
rlabel metal2 s 275296 0 275352 400 6 y[508]
port 1958 nsew signal input
rlabel metal2 s 275632 0 275688 400 6 y[509]
port 1959 nsew signal input
rlabel metal2 s 121408 0 121464 400 6 y[50]
port 1960 nsew signal input
rlabel metal2 s 275968 0 276024 400 6 y[510]
port 1961 nsew signal input
rlabel metal2 s 276304 0 276360 400 6 y[511]
port 1962 nsew signal input
rlabel metal2 s 121744 0 121800 400 6 y[51]
port 1963 nsew signal input
rlabel metal2 s 122080 0 122136 400 6 y[52]
port 1964 nsew signal input
rlabel metal2 s 122416 0 122472 400 6 y[53]
port 1965 nsew signal input
rlabel metal2 s 122752 0 122808 400 6 y[54]
port 1966 nsew signal input
rlabel metal2 s 123088 0 123144 400 6 y[55]
port 1967 nsew signal input
rlabel metal2 s 123424 0 123480 400 6 y[56]
port 1968 nsew signal input
rlabel metal2 s 123760 0 123816 400 6 y[57]
port 1969 nsew signal input
rlabel metal2 s 124096 0 124152 400 6 y[58]
port 1970 nsew signal input
rlabel metal2 s 124432 0 124488 400 6 y[59]
port 1971 nsew signal input
rlabel metal2 s 106288 0 106344 400 6 y[5]
port 1972 nsew signal input
rlabel metal2 s 124768 0 124824 400 6 y[60]
port 1973 nsew signal input
rlabel metal2 s 125104 0 125160 400 6 y[61]
port 1974 nsew signal input
rlabel metal2 s 125440 0 125496 400 6 y[62]
port 1975 nsew signal input
rlabel metal2 s 125776 0 125832 400 6 y[63]
port 1976 nsew signal input
rlabel metal2 s 126112 0 126168 400 6 y[64]
port 1977 nsew signal input
rlabel metal2 s 126448 0 126504 400 6 y[65]
port 1978 nsew signal input
rlabel metal2 s 126784 0 126840 400 6 y[66]
port 1979 nsew signal input
rlabel metal2 s 127120 0 127176 400 6 y[67]
port 1980 nsew signal input
rlabel metal2 s 127456 0 127512 400 6 y[68]
port 1981 nsew signal input
rlabel metal2 s 127792 0 127848 400 6 y[69]
port 1982 nsew signal input
rlabel metal2 s 106624 0 106680 400 6 y[6]
port 1983 nsew signal input
rlabel metal2 s 128128 0 128184 400 6 y[70]
port 1984 nsew signal input
rlabel metal2 s 128464 0 128520 400 6 y[71]
port 1985 nsew signal input
rlabel metal2 s 128800 0 128856 400 6 y[72]
port 1986 nsew signal input
rlabel metal2 s 129136 0 129192 400 6 y[73]
port 1987 nsew signal input
rlabel metal2 s 129472 0 129528 400 6 y[74]
port 1988 nsew signal input
rlabel metal2 s 129808 0 129864 400 6 y[75]
port 1989 nsew signal input
rlabel metal2 s 130144 0 130200 400 6 y[76]
port 1990 nsew signal input
rlabel metal2 s 130480 0 130536 400 6 y[77]
port 1991 nsew signal input
rlabel metal2 s 130816 0 130872 400 6 y[78]
port 1992 nsew signal input
rlabel metal2 s 131152 0 131208 400 6 y[79]
port 1993 nsew signal input
rlabel metal2 s 106960 0 107016 400 6 y[7]
port 1994 nsew signal input
rlabel metal2 s 131488 0 131544 400 6 y[80]
port 1995 nsew signal input
rlabel metal2 s 131824 0 131880 400 6 y[81]
port 1996 nsew signal input
rlabel metal2 s 132160 0 132216 400 6 y[82]
port 1997 nsew signal input
rlabel metal2 s 132496 0 132552 400 6 y[83]
port 1998 nsew signal input
rlabel metal2 s 132832 0 132888 400 6 y[84]
port 1999 nsew signal input
rlabel metal2 s 133168 0 133224 400 6 y[85]
port 2000 nsew signal input
rlabel metal2 s 133504 0 133560 400 6 y[86]
port 2001 nsew signal input
rlabel metal2 s 133840 0 133896 400 6 y[87]
port 2002 nsew signal input
rlabel metal2 s 134176 0 134232 400 6 y[88]
port 2003 nsew signal input
rlabel metal2 s 134512 0 134568 400 6 y[89]
port 2004 nsew signal input
rlabel metal2 s 107296 0 107352 400 6 y[8]
port 2005 nsew signal input
rlabel metal2 s 134848 0 134904 400 6 y[90]
port 2006 nsew signal input
rlabel metal2 s 135184 0 135240 400 6 y[91]
port 2007 nsew signal input
rlabel metal2 s 135520 0 135576 400 6 y[92]
port 2008 nsew signal input
rlabel metal2 s 135856 0 135912 400 6 y[93]
port 2009 nsew signal input
rlabel metal2 s 136192 0 136248 400 6 y[94]
port 2010 nsew signal input
rlabel metal2 s 136528 0 136584 400 6 y[95]
port 2011 nsew signal input
rlabel metal2 s 136864 0 136920 400 6 y[96]
port 2012 nsew signal input
rlabel metal2 s 137200 0 137256 400 6 y[97]
port 2013 nsew signal input
rlabel metal2 s 137536 0 137592 400 6 y[98]
port 2014 nsew signal input
rlabel metal2 s 137872 0 137928 400 6 y[99]
port 2015 nsew signal input
rlabel metal2 s 107632 0 107688 400 6 y[9]
port 2016 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8024524
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/tjrpu/runs/23_11_20_09_11/results/signoff/tjrpu.magic.gds
string GDS_START 220450
<< end >>

