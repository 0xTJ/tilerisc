magic
tech gf180mcuD
magscale 1 5
timestamp 1700946866
<< obsm1 >>
rect 672 1471 54320 58561
<< metal2 >>
rect 3920 59600 3976 60000
rect 4368 59600 4424 60000
rect 4816 59600 4872 60000
rect 5264 59600 5320 60000
rect 5712 59600 5768 60000
rect 6160 59600 6216 60000
rect 6608 59600 6664 60000
rect 7056 59600 7112 60000
rect 7504 59600 7560 60000
rect 7952 59600 8008 60000
rect 8400 59600 8456 60000
rect 8848 59600 8904 60000
rect 9296 59600 9352 60000
rect 9744 59600 9800 60000
rect 10192 59600 10248 60000
rect 10640 59600 10696 60000
rect 11088 59600 11144 60000
rect 11536 59600 11592 60000
rect 11984 59600 12040 60000
rect 12432 59600 12488 60000
rect 12880 59600 12936 60000
rect 13328 59600 13384 60000
rect 13776 59600 13832 60000
rect 14224 59600 14280 60000
rect 14672 59600 14728 60000
rect 15120 59600 15176 60000
rect 15568 59600 15624 60000
rect 16016 59600 16072 60000
rect 16464 59600 16520 60000
rect 16912 59600 16968 60000
rect 17360 59600 17416 60000
rect 17808 59600 17864 60000
rect 18256 59600 18312 60000
rect 18704 59600 18760 60000
rect 19152 59600 19208 60000
rect 19600 59600 19656 60000
rect 20048 59600 20104 60000
rect 20496 59600 20552 60000
rect 20944 59600 21000 60000
rect 21392 59600 21448 60000
rect 21840 59600 21896 60000
rect 22288 59600 22344 60000
rect 22736 59600 22792 60000
rect 23184 59600 23240 60000
rect 23632 59600 23688 60000
rect 24080 59600 24136 60000
rect 24528 59600 24584 60000
rect 24976 59600 25032 60000
rect 25424 59600 25480 60000
rect 25872 59600 25928 60000
rect 26320 59600 26376 60000
rect 26768 59600 26824 60000
rect 27216 59600 27272 60000
rect 27664 59600 27720 60000
rect 28112 59600 28168 60000
rect 28560 59600 28616 60000
rect 29008 59600 29064 60000
rect 29456 59600 29512 60000
rect 29904 59600 29960 60000
rect 30352 59600 30408 60000
rect 30800 59600 30856 60000
rect 31248 59600 31304 60000
rect 31696 59600 31752 60000
rect 32144 59600 32200 60000
rect 32592 59600 32648 60000
rect 33040 59600 33096 60000
rect 33488 59600 33544 60000
rect 33936 59600 33992 60000
rect 34384 59600 34440 60000
rect 34832 59600 34888 60000
rect 35280 59600 35336 60000
rect 35728 59600 35784 60000
rect 36176 59600 36232 60000
rect 36624 59600 36680 60000
rect 37072 59600 37128 60000
rect 37520 59600 37576 60000
rect 37968 59600 38024 60000
rect 38416 59600 38472 60000
rect 38864 59600 38920 60000
rect 39312 59600 39368 60000
rect 39760 59600 39816 60000
rect 40208 59600 40264 60000
rect 40656 59600 40712 60000
rect 41104 59600 41160 60000
rect 41552 59600 41608 60000
rect 42000 59600 42056 60000
rect 42448 59600 42504 60000
rect 42896 59600 42952 60000
rect 43344 59600 43400 60000
rect 43792 59600 43848 60000
rect 44240 59600 44296 60000
rect 44688 59600 44744 60000
rect 45136 59600 45192 60000
rect 45584 59600 45640 60000
rect 46032 59600 46088 60000
rect 46480 59600 46536 60000
rect 46928 59600 46984 60000
rect 47376 59600 47432 60000
rect 47824 59600 47880 60000
rect 48272 59600 48328 60000
rect 48720 59600 48776 60000
rect 49168 59600 49224 60000
rect 49616 59600 49672 60000
rect 50064 59600 50120 60000
rect 50512 59600 50568 60000
rect 50960 59600 51016 60000
rect 560 0 616 400
rect 1120 0 1176 400
rect 1680 0 1736 400
rect 2240 0 2296 400
rect 2800 0 2856 400
rect 3360 0 3416 400
rect 3920 0 3976 400
rect 4480 0 4536 400
rect 5040 0 5096 400
rect 5600 0 5656 400
rect 6160 0 6216 400
rect 6720 0 6776 400
rect 7280 0 7336 400
rect 7840 0 7896 400
rect 8400 0 8456 400
rect 8960 0 9016 400
rect 9520 0 9576 400
rect 10080 0 10136 400
rect 10640 0 10696 400
rect 11200 0 11256 400
rect 11760 0 11816 400
rect 12320 0 12376 400
rect 12880 0 12936 400
rect 13440 0 13496 400
rect 14000 0 14056 400
rect 14560 0 14616 400
rect 15120 0 15176 400
rect 15680 0 15736 400
rect 16240 0 16296 400
rect 16800 0 16856 400
rect 17360 0 17416 400
rect 17920 0 17976 400
rect 18480 0 18536 400
rect 19040 0 19096 400
rect 19600 0 19656 400
rect 20160 0 20216 400
rect 20720 0 20776 400
rect 21280 0 21336 400
rect 21840 0 21896 400
rect 22400 0 22456 400
rect 22960 0 23016 400
rect 23520 0 23576 400
rect 24080 0 24136 400
rect 24640 0 24696 400
rect 25200 0 25256 400
rect 25760 0 25816 400
rect 26320 0 26376 400
rect 26880 0 26936 400
rect 27440 0 27496 400
rect 28000 0 28056 400
rect 28560 0 28616 400
rect 29120 0 29176 400
rect 29680 0 29736 400
rect 30240 0 30296 400
rect 30800 0 30856 400
rect 31360 0 31416 400
rect 31920 0 31976 400
rect 32480 0 32536 400
rect 33040 0 33096 400
rect 33600 0 33656 400
rect 34160 0 34216 400
rect 34720 0 34776 400
rect 35280 0 35336 400
rect 35840 0 35896 400
rect 36400 0 36456 400
rect 36960 0 37016 400
rect 37520 0 37576 400
rect 38080 0 38136 400
rect 38640 0 38696 400
rect 39200 0 39256 400
rect 39760 0 39816 400
rect 40320 0 40376 400
rect 40880 0 40936 400
rect 41440 0 41496 400
rect 42000 0 42056 400
rect 42560 0 42616 400
rect 43120 0 43176 400
rect 43680 0 43736 400
rect 44240 0 44296 400
rect 44800 0 44856 400
rect 45360 0 45416 400
rect 45920 0 45976 400
rect 46480 0 46536 400
rect 47040 0 47096 400
rect 47600 0 47656 400
rect 48160 0 48216 400
rect 48720 0 48776 400
rect 49280 0 49336 400
rect 49840 0 49896 400
rect 50400 0 50456 400
rect 50960 0 51016 400
rect 51520 0 51576 400
rect 52080 0 52136 400
rect 52640 0 52696 400
rect 53200 0 53256 400
rect 53760 0 53816 400
rect 54320 0 54376 400
<< obsm2 >>
rect 574 59570 3890 59682
rect 4006 59570 4338 59682
rect 4454 59570 4786 59682
rect 4902 59570 5234 59682
rect 5350 59570 5682 59682
rect 5798 59570 6130 59682
rect 6246 59570 6578 59682
rect 6694 59570 7026 59682
rect 7142 59570 7474 59682
rect 7590 59570 7922 59682
rect 8038 59570 8370 59682
rect 8486 59570 8818 59682
rect 8934 59570 9266 59682
rect 9382 59570 9714 59682
rect 9830 59570 10162 59682
rect 10278 59570 10610 59682
rect 10726 59570 11058 59682
rect 11174 59570 11506 59682
rect 11622 59570 11954 59682
rect 12070 59570 12402 59682
rect 12518 59570 12850 59682
rect 12966 59570 13298 59682
rect 13414 59570 13746 59682
rect 13862 59570 14194 59682
rect 14310 59570 14642 59682
rect 14758 59570 15090 59682
rect 15206 59570 15538 59682
rect 15654 59570 15986 59682
rect 16102 59570 16434 59682
rect 16550 59570 16882 59682
rect 16998 59570 17330 59682
rect 17446 59570 17778 59682
rect 17894 59570 18226 59682
rect 18342 59570 18674 59682
rect 18790 59570 19122 59682
rect 19238 59570 19570 59682
rect 19686 59570 20018 59682
rect 20134 59570 20466 59682
rect 20582 59570 20914 59682
rect 21030 59570 21362 59682
rect 21478 59570 21810 59682
rect 21926 59570 22258 59682
rect 22374 59570 22706 59682
rect 22822 59570 23154 59682
rect 23270 59570 23602 59682
rect 23718 59570 24050 59682
rect 24166 59570 24498 59682
rect 24614 59570 24946 59682
rect 25062 59570 25394 59682
rect 25510 59570 25842 59682
rect 25958 59570 26290 59682
rect 26406 59570 26738 59682
rect 26854 59570 27186 59682
rect 27302 59570 27634 59682
rect 27750 59570 28082 59682
rect 28198 59570 28530 59682
rect 28646 59570 28978 59682
rect 29094 59570 29426 59682
rect 29542 59570 29874 59682
rect 29990 59570 30322 59682
rect 30438 59570 30770 59682
rect 30886 59570 31218 59682
rect 31334 59570 31666 59682
rect 31782 59570 32114 59682
rect 32230 59570 32562 59682
rect 32678 59570 33010 59682
rect 33126 59570 33458 59682
rect 33574 59570 33906 59682
rect 34022 59570 34354 59682
rect 34470 59570 34802 59682
rect 34918 59570 35250 59682
rect 35366 59570 35698 59682
rect 35814 59570 36146 59682
rect 36262 59570 36594 59682
rect 36710 59570 37042 59682
rect 37158 59570 37490 59682
rect 37606 59570 37938 59682
rect 38054 59570 38386 59682
rect 38502 59570 38834 59682
rect 38950 59570 39282 59682
rect 39398 59570 39730 59682
rect 39846 59570 40178 59682
rect 40294 59570 40626 59682
rect 40742 59570 41074 59682
rect 41190 59570 41522 59682
rect 41638 59570 41970 59682
rect 42086 59570 42418 59682
rect 42534 59570 42866 59682
rect 42982 59570 43314 59682
rect 43430 59570 43762 59682
rect 43878 59570 44210 59682
rect 44326 59570 44658 59682
rect 44774 59570 45106 59682
rect 45222 59570 45554 59682
rect 45670 59570 46002 59682
rect 46118 59570 46450 59682
rect 46566 59570 46898 59682
rect 47014 59570 47346 59682
rect 47462 59570 47794 59682
rect 47910 59570 48242 59682
rect 48358 59570 48690 59682
rect 48806 59570 49138 59682
rect 49254 59570 49586 59682
rect 49702 59570 50034 59682
rect 50150 59570 50482 59682
rect 50598 59570 50930 59682
rect 51046 59570 54418 59682
rect 574 430 54418 59570
rect 646 350 1090 430
rect 1206 350 1650 430
rect 1766 350 2210 430
rect 2326 350 2770 430
rect 2886 350 3330 430
rect 3446 350 3890 430
rect 4006 350 4450 430
rect 4566 350 5010 430
rect 5126 350 5570 430
rect 5686 350 6130 430
rect 6246 350 6690 430
rect 6806 350 7250 430
rect 7366 350 7810 430
rect 7926 350 8370 430
rect 8486 350 8930 430
rect 9046 350 9490 430
rect 9606 350 10050 430
rect 10166 350 10610 430
rect 10726 350 11170 430
rect 11286 350 11730 430
rect 11846 350 12290 430
rect 12406 350 12850 430
rect 12966 350 13410 430
rect 13526 350 13970 430
rect 14086 350 14530 430
rect 14646 350 15090 430
rect 15206 350 15650 430
rect 15766 350 16210 430
rect 16326 350 16770 430
rect 16886 350 17330 430
rect 17446 350 17890 430
rect 18006 350 18450 430
rect 18566 350 19010 430
rect 19126 350 19570 430
rect 19686 350 20130 430
rect 20246 350 20690 430
rect 20806 350 21250 430
rect 21366 350 21810 430
rect 21926 350 22370 430
rect 22486 350 22930 430
rect 23046 350 23490 430
rect 23606 350 24050 430
rect 24166 350 24610 430
rect 24726 350 25170 430
rect 25286 350 25730 430
rect 25846 350 26290 430
rect 26406 350 26850 430
rect 26966 350 27410 430
rect 27526 350 27970 430
rect 28086 350 28530 430
rect 28646 350 29090 430
rect 29206 350 29650 430
rect 29766 350 30210 430
rect 30326 350 30770 430
rect 30886 350 31330 430
rect 31446 350 31890 430
rect 32006 350 32450 430
rect 32566 350 33010 430
rect 33126 350 33570 430
rect 33686 350 34130 430
rect 34246 350 34690 430
rect 34806 350 35250 430
rect 35366 350 35810 430
rect 35926 350 36370 430
rect 36486 350 36930 430
rect 37046 350 37490 430
rect 37606 350 38050 430
rect 38166 350 38610 430
rect 38726 350 39170 430
rect 39286 350 39730 430
rect 39846 350 40290 430
rect 40406 350 40850 430
rect 40966 350 41410 430
rect 41526 350 41970 430
rect 42086 350 42530 430
rect 42646 350 43090 430
rect 43206 350 43650 430
rect 43766 350 44210 430
rect 44326 350 44770 430
rect 44886 350 45330 430
rect 45446 350 45890 430
rect 46006 350 46450 430
rect 46566 350 47010 430
rect 47126 350 47570 430
rect 47686 350 48130 430
rect 48246 350 48690 430
rect 48806 350 49250 430
rect 49366 350 49810 430
rect 49926 350 50370 430
rect 50486 350 50930 430
rect 51046 350 51490 430
rect 51606 350 52050 430
rect 52166 350 52610 430
rect 52726 350 53170 430
rect 53286 350 53730 430
rect 53846 350 54290 430
rect 54406 350 54418 430
<< obsm3 >>
rect 569 686 54423 58898
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
<< obsm4 >>
rect 4662 58468 54194 58847
rect 4662 1508 9874 58468
rect 10094 1508 17554 58468
rect 17774 1508 25234 58468
rect 25454 1508 32914 58468
rect 33134 1508 40594 58468
rect 40814 1508 48274 58468
rect 48494 1508 54194 58468
rect 4662 681 54194 1508
<< labels >>
rlabel metal2 s 560 0 616 400 6 clk
port 1 nsew signal input
rlabel metal2 s 1120 0 1176 400 6 inst[0]
port 2 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 inst[10]
port 3 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 inst[11]
port 4 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 inst[12]
port 5 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 inst[13]
port 6 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 inst[14]
port 7 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 inst[15]
port 8 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 inst[16]
port 9 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 inst[17]
port 10 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 inst[18]
port 11 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 inst[19]
port 12 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 inst[1]
port 13 nsew signal input
rlabel metal2 s 12320 0 12376 400 6 inst[20]
port 14 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 inst[21]
port 15 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 inst[22]
port 16 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 inst[23]
port 17 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 inst[24]
port 18 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 inst[25]
port 19 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 inst[26]
port 20 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 inst[27]
port 21 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 inst[28]
port 22 nsew signal input
rlabel metal2 s 17360 0 17416 400 6 inst[29]
port 23 nsew signal input
rlabel metal2 s 2240 0 2296 400 6 inst[2]
port 24 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 inst[30]
port 25 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 inst[31]
port 26 nsew signal input
rlabel metal2 s 2800 0 2856 400 6 inst[3]
port 27 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 inst[4]
port 28 nsew signal input
rlabel metal2 s 3920 0 3976 400 6 inst[5]
port 29 nsew signal input
rlabel metal2 s 4480 0 4536 400 6 inst[6]
port 30 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 inst[7]
port 31 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 inst[8]
port 32 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 inst[9]
port 33 nsew signal input
rlabel metal2 s 50960 59600 51016 60000 6 mem_addr[0]
port 34 nsew signal output
rlabel metal2 s 46480 59600 46536 60000 6 mem_addr[10]
port 35 nsew signal output
rlabel metal2 s 46032 59600 46088 60000 6 mem_addr[11]
port 36 nsew signal output
rlabel metal2 s 45584 59600 45640 60000 6 mem_addr[12]
port 37 nsew signal output
rlabel metal2 s 45136 59600 45192 60000 6 mem_addr[13]
port 38 nsew signal output
rlabel metal2 s 44688 59600 44744 60000 6 mem_addr[14]
port 39 nsew signal output
rlabel metal2 s 44240 59600 44296 60000 6 mem_addr[15]
port 40 nsew signal output
rlabel metal2 s 43792 59600 43848 60000 6 mem_addr[16]
port 41 nsew signal output
rlabel metal2 s 43344 59600 43400 60000 6 mem_addr[17]
port 42 nsew signal output
rlabel metal2 s 42896 59600 42952 60000 6 mem_addr[18]
port 43 nsew signal output
rlabel metal2 s 42448 59600 42504 60000 6 mem_addr[19]
port 44 nsew signal output
rlabel metal2 s 50512 59600 50568 60000 6 mem_addr[1]
port 45 nsew signal output
rlabel metal2 s 42000 59600 42056 60000 6 mem_addr[20]
port 46 nsew signal output
rlabel metal2 s 41552 59600 41608 60000 6 mem_addr[21]
port 47 nsew signal output
rlabel metal2 s 41104 59600 41160 60000 6 mem_addr[22]
port 48 nsew signal output
rlabel metal2 s 40656 59600 40712 60000 6 mem_addr[23]
port 49 nsew signal output
rlabel metal2 s 40208 59600 40264 60000 6 mem_addr[24]
port 50 nsew signal output
rlabel metal2 s 39760 59600 39816 60000 6 mem_addr[25]
port 51 nsew signal output
rlabel metal2 s 39312 59600 39368 60000 6 mem_addr[26]
port 52 nsew signal output
rlabel metal2 s 38864 59600 38920 60000 6 mem_addr[27]
port 53 nsew signal output
rlabel metal2 s 38416 59600 38472 60000 6 mem_addr[28]
port 54 nsew signal output
rlabel metal2 s 37968 59600 38024 60000 6 mem_addr[29]
port 55 nsew signal output
rlabel metal2 s 50064 59600 50120 60000 6 mem_addr[2]
port 56 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 mem_addr[30]
port 57 nsew signal output
rlabel metal2 s 37072 59600 37128 60000 6 mem_addr[31]
port 58 nsew signal output
rlabel metal2 s 49616 59600 49672 60000 6 mem_addr[3]
port 59 nsew signal output
rlabel metal2 s 49168 59600 49224 60000 6 mem_addr[4]
port 60 nsew signal output
rlabel metal2 s 48720 59600 48776 60000 6 mem_addr[5]
port 61 nsew signal output
rlabel metal2 s 48272 59600 48328 60000 6 mem_addr[6]
port 62 nsew signal output
rlabel metal2 s 47824 59600 47880 60000 6 mem_addr[7]
port 63 nsew signal output
rlabel metal2 s 47376 59600 47432 60000 6 mem_addr[8]
port 64 nsew signal output
rlabel metal2 s 46928 59600 46984 60000 6 mem_addr[9]
port 65 nsew signal output
rlabel metal2 s 34384 59600 34440 60000 6 mem_ld_dat[0]
port 66 nsew signal input
rlabel metal2 s 29904 59600 29960 60000 6 mem_ld_dat[10]
port 67 nsew signal input
rlabel metal2 s 29456 59600 29512 60000 6 mem_ld_dat[11]
port 68 nsew signal input
rlabel metal2 s 29008 59600 29064 60000 6 mem_ld_dat[12]
port 69 nsew signal input
rlabel metal2 s 28560 59600 28616 60000 6 mem_ld_dat[13]
port 70 nsew signal input
rlabel metal2 s 28112 59600 28168 60000 6 mem_ld_dat[14]
port 71 nsew signal input
rlabel metal2 s 27664 59600 27720 60000 6 mem_ld_dat[15]
port 72 nsew signal input
rlabel metal2 s 27216 59600 27272 60000 6 mem_ld_dat[16]
port 73 nsew signal input
rlabel metal2 s 26768 59600 26824 60000 6 mem_ld_dat[17]
port 74 nsew signal input
rlabel metal2 s 26320 59600 26376 60000 6 mem_ld_dat[18]
port 75 nsew signal input
rlabel metal2 s 25872 59600 25928 60000 6 mem_ld_dat[19]
port 76 nsew signal input
rlabel metal2 s 33936 59600 33992 60000 6 mem_ld_dat[1]
port 77 nsew signal input
rlabel metal2 s 25424 59600 25480 60000 6 mem_ld_dat[20]
port 78 nsew signal input
rlabel metal2 s 24976 59600 25032 60000 6 mem_ld_dat[21]
port 79 nsew signal input
rlabel metal2 s 24528 59600 24584 60000 6 mem_ld_dat[22]
port 80 nsew signal input
rlabel metal2 s 24080 59600 24136 60000 6 mem_ld_dat[23]
port 81 nsew signal input
rlabel metal2 s 23632 59600 23688 60000 6 mem_ld_dat[24]
port 82 nsew signal input
rlabel metal2 s 23184 59600 23240 60000 6 mem_ld_dat[25]
port 83 nsew signal input
rlabel metal2 s 22736 59600 22792 60000 6 mem_ld_dat[26]
port 84 nsew signal input
rlabel metal2 s 22288 59600 22344 60000 6 mem_ld_dat[27]
port 85 nsew signal input
rlabel metal2 s 21840 59600 21896 60000 6 mem_ld_dat[28]
port 86 nsew signal input
rlabel metal2 s 21392 59600 21448 60000 6 mem_ld_dat[29]
port 87 nsew signal input
rlabel metal2 s 33488 59600 33544 60000 6 mem_ld_dat[2]
port 88 nsew signal input
rlabel metal2 s 20944 59600 21000 60000 6 mem_ld_dat[30]
port 89 nsew signal input
rlabel metal2 s 20496 59600 20552 60000 6 mem_ld_dat[31]
port 90 nsew signal input
rlabel metal2 s 33040 59600 33096 60000 6 mem_ld_dat[3]
port 91 nsew signal input
rlabel metal2 s 32592 59600 32648 60000 6 mem_ld_dat[4]
port 92 nsew signal input
rlabel metal2 s 32144 59600 32200 60000 6 mem_ld_dat[5]
port 93 nsew signal input
rlabel metal2 s 31696 59600 31752 60000 6 mem_ld_dat[6]
port 94 nsew signal input
rlabel metal2 s 31248 59600 31304 60000 6 mem_ld_dat[7]
port 95 nsew signal input
rlabel metal2 s 30800 59600 30856 60000 6 mem_ld_dat[8]
port 96 nsew signal input
rlabel metal2 s 30352 59600 30408 60000 6 mem_ld_dat[9]
port 97 nsew signal input
rlabel metal2 s 36624 59600 36680 60000 6 mem_ld_en
port 98 nsew signal output
rlabel metal2 s 36176 59600 36232 60000 6 mem_ld_mask[0]
port 99 nsew signal output
rlabel metal2 s 35728 59600 35784 60000 6 mem_ld_mask[1]
port 100 nsew signal output
rlabel metal2 s 35280 59600 35336 60000 6 mem_ld_mask[2]
port 101 nsew signal output
rlabel metal2 s 34832 59600 34888 60000 6 mem_ld_mask[3]
port 102 nsew signal output
rlabel metal2 s 17808 59600 17864 60000 6 mem_st_dat[0]
port 103 nsew signal output
rlabel metal2 s 13328 59600 13384 60000 6 mem_st_dat[10]
port 104 nsew signal output
rlabel metal2 s 12880 59600 12936 60000 6 mem_st_dat[11]
port 105 nsew signal output
rlabel metal2 s 12432 59600 12488 60000 6 mem_st_dat[12]
port 106 nsew signal output
rlabel metal2 s 11984 59600 12040 60000 6 mem_st_dat[13]
port 107 nsew signal output
rlabel metal2 s 11536 59600 11592 60000 6 mem_st_dat[14]
port 108 nsew signal output
rlabel metal2 s 11088 59600 11144 60000 6 mem_st_dat[15]
port 109 nsew signal output
rlabel metal2 s 10640 59600 10696 60000 6 mem_st_dat[16]
port 110 nsew signal output
rlabel metal2 s 10192 59600 10248 60000 6 mem_st_dat[17]
port 111 nsew signal output
rlabel metal2 s 9744 59600 9800 60000 6 mem_st_dat[18]
port 112 nsew signal output
rlabel metal2 s 9296 59600 9352 60000 6 mem_st_dat[19]
port 113 nsew signal output
rlabel metal2 s 17360 59600 17416 60000 6 mem_st_dat[1]
port 114 nsew signal output
rlabel metal2 s 8848 59600 8904 60000 6 mem_st_dat[20]
port 115 nsew signal output
rlabel metal2 s 8400 59600 8456 60000 6 mem_st_dat[21]
port 116 nsew signal output
rlabel metal2 s 7952 59600 8008 60000 6 mem_st_dat[22]
port 117 nsew signal output
rlabel metal2 s 7504 59600 7560 60000 6 mem_st_dat[23]
port 118 nsew signal output
rlabel metal2 s 7056 59600 7112 60000 6 mem_st_dat[24]
port 119 nsew signal output
rlabel metal2 s 6608 59600 6664 60000 6 mem_st_dat[25]
port 120 nsew signal output
rlabel metal2 s 6160 59600 6216 60000 6 mem_st_dat[26]
port 121 nsew signal output
rlabel metal2 s 5712 59600 5768 60000 6 mem_st_dat[27]
port 122 nsew signal output
rlabel metal2 s 5264 59600 5320 60000 6 mem_st_dat[28]
port 123 nsew signal output
rlabel metal2 s 4816 59600 4872 60000 6 mem_st_dat[29]
port 124 nsew signal output
rlabel metal2 s 16912 59600 16968 60000 6 mem_st_dat[2]
port 125 nsew signal output
rlabel metal2 s 4368 59600 4424 60000 6 mem_st_dat[30]
port 126 nsew signal output
rlabel metal2 s 3920 59600 3976 60000 6 mem_st_dat[31]
port 127 nsew signal output
rlabel metal2 s 16464 59600 16520 60000 6 mem_st_dat[3]
port 128 nsew signal output
rlabel metal2 s 16016 59600 16072 60000 6 mem_st_dat[4]
port 129 nsew signal output
rlabel metal2 s 15568 59600 15624 60000 6 mem_st_dat[5]
port 130 nsew signal output
rlabel metal2 s 15120 59600 15176 60000 6 mem_st_dat[6]
port 131 nsew signal output
rlabel metal2 s 14672 59600 14728 60000 6 mem_st_dat[7]
port 132 nsew signal output
rlabel metal2 s 14224 59600 14280 60000 6 mem_st_dat[8]
port 133 nsew signal output
rlabel metal2 s 13776 59600 13832 60000 6 mem_st_dat[9]
port 134 nsew signal output
rlabel metal2 s 20048 59600 20104 60000 6 mem_st_en
port 135 nsew signal output
rlabel metal2 s 19600 59600 19656 60000 6 mem_st_mask[0]
port 136 nsew signal output
rlabel metal2 s 19152 59600 19208 60000 6 mem_st_mask[1]
port 137 nsew signal output
rlabel metal2 s 18704 59600 18760 60000 6 mem_st_mask[2]
port 138 nsew signal output
rlabel metal2 s 18256 59600 18312 60000 6 mem_st_mask[3]
port 139 nsew signal output
rlabel metal2 s 19040 0 19096 400 6 pc[0]
port 140 nsew signal input
rlabel metal2 s 24640 0 24696 400 6 pc[10]
port 141 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 pc[11]
port 142 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 pc[12]
port 143 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 pc[13]
port 144 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 pc[14]
port 145 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 pc[15]
port 146 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 pc[16]
port 147 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 pc[17]
port 148 nsew signal input
rlabel metal2 s 29120 0 29176 400 6 pc[18]
port 149 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 pc[19]
port 150 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 pc[1]
port 151 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 pc[20]
port 152 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 pc[21]
port 153 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 pc[22]
port 154 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 pc[23]
port 155 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 pc[24]
port 156 nsew signal input
rlabel metal2 s 33040 0 33096 400 6 pc[25]
port 157 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 pc[26]
port 158 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 pc[27]
port 159 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 pc[28]
port 160 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 pc[29]
port 161 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 pc[2]
port 162 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 pc[30]
port 163 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 pc[31]
port 164 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 pc[3]
port 165 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 pc[4]
port 166 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 pc[5]
port 167 nsew signal input
rlabel metal2 s 22400 0 22456 400 6 pc[6]
port 168 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 pc[7]
port 169 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 pc[8]
port 170 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 pc[9]
port 171 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 pc_next[0]
port 172 nsew signal output
rlabel metal2 s 42560 0 42616 400 6 pc_next[10]
port 173 nsew signal output
rlabel metal2 s 43120 0 43176 400 6 pc_next[11]
port 174 nsew signal output
rlabel metal2 s 43680 0 43736 400 6 pc_next[12]
port 175 nsew signal output
rlabel metal2 s 44240 0 44296 400 6 pc_next[13]
port 176 nsew signal output
rlabel metal2 s 44800 0 44856 400 6 pc_next[14]
port 177 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 pc_next[15]
port 178 nsew signal output
rlabel metal2 s 45920 0 45976 400 6 pc_next[16]
port 179 nsew signal output
rlabel metal2 s 46480 0 46536 400 6 pc_next[17]
port 180 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 pc_next[18]
port 181 nsew signal output
rlabel metal2 s 47600 0 47656 400 6 pc_next[19]
port 182 nsew signal output
rlabel metal2 s 37520 0 37576 400 6 pc_next[1]
port 183 nsew signal output
rlabel metal2 s 48160 0 48216 400 6 pc_next[20]
port 184 nsew signal output
rlabel metal2 s 48720 0 48776 400 6 pc_next[21]
port 185 nsew signal output
rlabel metal2 s 49280 0 49336 400 6 pc_next[22]
port 186 nsew signal output
rlabel metal2 s 49840 0 49896 400 6 pc_next[23]
port 187 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 pc_next[24]
port 188 nsew signal output
rlabel metal2 s 50960 0 51016 400 6 pc_next[25]
port 189 nsew signal output
rlabel metal2 s 51520 0 51576 400 6 pc_next[26]
port 190 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 pc_next[27]
port 191 nsew signal output
rlabel metal2 s 52640 0 52696 400 6 pc_next[28]
port 192 nsew signal output
rlabel metal2 s 53200 0 53256 400 6 pc_next[29]
port 193 nsew signal output
rlabel metal2 s 38080 0 38136 400 6 pc_next[2]
port 194 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 pc_next[30]
port 195 nsew signal output
rlabel metal2 s 54320 0 54376 400 6 pc_next[31]
port 196 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 pc_next[3]
port 197 nsew signal output
rlabel metal2 s 39200 0 39256 400 6 pc_next[4]
port 198 nsew signal output
rlabel metal2 s 39760 0 39816 400 6 pc_next[5]
port 199 nsew signal output
rlabel metal2 s 40320 0 40376 400 6 pc_next[6]
port 200 nsew signal output
rlabel metal2 s 40880 0 40936 400 6 pc_next[7]
port 201 nsew signal output
rlabel metal2 s 41440 0 41496 400 6 pc_next[8]
port 202 nsew signal output
rlabel metal2 s 42000 0 42056 400 6 pc_next[9]
port 203 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 204 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 205 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 205 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 55000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11518434
string GDS_FILE /home/thomas/Documents/Projects/tilerisc/openlane/rv_core/runs/23_11_25_16_09/results/signoff/tinyrv.magic.gds
string GDS_START 534584
<< end >>

