VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180_ram_64x8_wrapper
  CLASS BLOCK ;
  FOREIGN gf180_ram_64x8_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 444.860 BY 243.880 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.720 239.880 265.280 243.880 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.220 239.880 273.780 243.880 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.720 239.880 282.280 243.880 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.720 239.880 155.280 243.880 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.720 239.880 160.280 243.880 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.720 239.880 164.280 243.880 ;
    END
  END A[5]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.220 239.880 184.780 243.880 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.220 239.880 296.780 243.880 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 239.880 427.280 243.880 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.720 239.880 375.280 243.880 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 368.720 239.880 369.280 243.880 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.720 239.880 317.280 243.880 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.720 239.880 129.280 243.880 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.220 239.880 77.780 243.880 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.720 239.880 71.280 243.880 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.720 239.880 19.280 243.880 ;
    END
  END D[7]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.840 239.880 233.400 243.880 ;
    END
  END GWEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 419.220 239.880 419.780 243.880 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.220 239.880 378.780 243.880 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.220 239.880 365.780 243.880 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.720 239.880 325.280 243.880 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.220 239.880 121.780 243.880 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.220 239.880 80.780 243.880 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.220 239.880 67.780 243.880 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.720 239.880 27.280 243.880 ;
    END
  END Q[7]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 5.220 15.680 8.220 227.360 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 428.630 15.680 431.630 227.360 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 9.220 15.680 12.220 227.360 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 432.630 15.680 435.630 227.360 ;
    END
  END VSS
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.220 239.880 423.780 243.880 ;
    END
  END WEN[0]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.720 239.880 373.280 243.880 ;
    END
  END WEN[1]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 239.880 371.280 243.880 ;
    END
  END WEN[2]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.720 239.880 319.280 243.880 ;
    END
  END WEN[3]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.220 239.880 125.780 243.880 ;
    END
  END WEN[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.970 239.880 75.530 243.880 ;
    END
  END WEN[5]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.720 239.880 73.280 243.880 ;
    END
  END WEN[6]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.220 239.880 22.780 243.880 ;
    END
  END WEN[7]
  OBS
      LAYER Metal1 ;
        RECT 5.000 5.000 436.860 237.880 ;
      LAYER Metal2 ;
        RECT 5.000 239.580 18.420 240.520 ;
        RECT 19.580 239.580 21.920 240.520 ;
        RECT 23.080 239.580 26.420 240.520 ;
        RECT 27.580 239.580 66.920 240.520 ;
        RECT 68.080 239.580 70.420 240.520 ;
        RECT 71.580 239.580 72.420 240.520 ;
        RECT 73.580 239.580 74.670 240.520 ;
        RECT 75.830 239.580 76.920 240.520 ;
        RECT 78.080 239.580 79.920 240.520 ;
        RECT 81.080 239.580 120.920 240.520 ;
        RECT 122.080 239.580 124.920 240.520 ;
        RECT 126.080 239.580 128.420 240.520 ;
        RECT 129.580 239.580 154.420 240.520 ;
        RECT 155.580 239.580 159.420 240.520 ;
        RECT 160.580 239.580 163.420 240.520 ;
        RECT 164.580 239.580 183.920 240.520 ;
        RECT 185.080 239.580 232.540 240.520 ;
        RECT 233.700 239.580 264.420 240.520 ;
        RECT 265.580 239.580 272.920 240.520 ;
        RECT 274.080 239.580 281.420 240.520 ;
        RECT 282.580 239.580 295.920 240.520 ;
        RECT 297.080 239.580 316.420 240.520 ;
        RECT 317.580 239.580 318.420 240.520 ;
        RECT 319.580 239.580 324.420 240.520 ;
        RECT 325.580 239.580 364.920 240.520 ;
        RECT 366.080 239.580 368.420 240.520 ;
        RECT 369.580 239.580 370.420 240.520 ;
        RECT 371.580 239.580 372.420 240.520 ;
        RECT 373.580 239.580 374.420 240.520 ;
        RECT 375.580 239.580 377.920 240.520 ;
        RECT 379.080 239.580 418.920 240.520 ;
        RECT 420.080 239.580 422.920 240.520 ;
        RECT 424.080 239.580 426.420 240.520 ;
        RECT 427.580 239.580 436.860 240.520 ;
        RECT 5.000 5.000 436.860 239.580 ;
      LAYER Metal3 ;
        RECT 5.000 5.000 436.860 237.880 ;
  END
END gf180_ram_64x8_wrapper
END LIBRARY

