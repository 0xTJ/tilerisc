* NGSPICE file created from interp_tri.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

.subckt interp_tri clk vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[2] wbs_adr_i[3]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ x_end[0] x_end[1] x_end[2] x_end[3] x_end[4] x_end[5] x_end[6] x_end[7] x_start[0]
+ x_start[1] x_start[2] x_start[3] x_start[4] x_start[5] x_start[6] x_start[7] y[0]
+ y[1] y[2] y[3] y[4] y[5] y[6] y[7]
X_2106_ _1290_ _1291_ _1292_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2037_ _1162_ _1168_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output37_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer7 _0178_ net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1996__A2 _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ _0007_ clknet_1_0__leaf_clk net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2655_ net21 _0500_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1606_ _0731_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_14_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2586_ _0334_ _0448_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1537_ _0672_ _0609_ _0613_ _0728_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1468_ _0651_ _0656_ _0659_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1399_ _0590_ _0591_ t_reg\[1\] _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_37_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1902__A2 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2526__C _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2440_ _0308_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_11_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2371_ _0260_ _0222_ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__A1 _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2707_ net19 _0531_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2638_ _0494_ _0495_ _0491_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2569_ _0443_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input36_I y[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1940_ _1042_ _1128_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1871_ _0971_ _0974_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2423_ _0157_ _1136_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2354_ _0897_ _0246_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2285_ _0151_ _0155_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2294__A1 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _1200_ _1257_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1923_ _1028_ _1108_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1785_ _0968_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1854_ _0924_ _0965_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2406_ _0252_ _0291_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2337_ _0174_ _0228_ _0229_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2268_ _0156_ _0162_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2199_ c\[0\]\[0\] _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2733__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2276__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__A1 _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0674_ _0761_ _0762_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2122_ _1196_ _1259_ _1308_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2053_ _1224_ _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xrebuffer17 _0802_ net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_16_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1837_ _0673_ _1024_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1768_ _0919_ _0940_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _1088_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _0811_ _0825_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput53 net53 x_start[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput42 net42 x_end[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2671_ net10 _0510_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ _0023_ clknet_1_0__leaf_clk t_reg\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1622_ delta_t\[9\] _0754_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1553_ _0744_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1484_ _0621_ _0675_ _0676_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2191__A3 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2105_ _1243_ _1245_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2036_ _1174_ _1175_ _1223_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2403__A1 _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer8 _0599_ net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2723_ _0006_ clknet_1_1__leaf_clk net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2654_ _1181_ _0498_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1536_ _0728_ _0672_ _0608_ _0613_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1605_ _0726_ _0796_ net84 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2585_ _0296_ _0448_ _0455_ _0453_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1398_ _0570_ _0572_ _0575_ _0577_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_38_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1467_ _0645_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2019_ _1147_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_19_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1666__A2 _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2615__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2091__A2 _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2370_ _0099_ _0080_ _1130_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _0544_ _0545_ _0540_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2499_ _0363_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2637_ net16 _0489_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1519_ _0637_ _0662_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2568_ _0443_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input29_I y[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1870_ _0971_ _0974_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ _0208_ _0245_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2422_ _0261_ _0312_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2284_ _0879_ _0983_ _0177_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_19_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2055__A2 _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1999_ _1144_ _1147_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_30_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1922_ _1029_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1853_ _0968_ _0975_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1784_ _0970_ _0971_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_24_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _1113_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2336_ _0122_ _1047_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2267_ _0158_ _0161_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2198_ _0079_ _0081_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2276__A2 _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2121_ _1197_ _1258_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer18 _0735_ net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__1702__A1 a\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2052_ _1226_ _1239_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_32_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _1093_ _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1836_ _1026_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1767_ _0877_ _0916_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1698_ _0887_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2319_ _0171_ _0210_ _0211_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input11_I wbs_dat_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput43 net43 x_end[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_33_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1781__I _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2723__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2670_ b\[1\]\[3\] _0513_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1552_ _0681_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1621_ _0584_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2104_ _1243_ _1245_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input3_I wbs_adr_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ _0634_ _0635_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2035_ _1155_ _0934_ _1172_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1819_ _0838_ _0839_ _0807_ _0552_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer9 _0797_ net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2633__A2 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2722_ _0005_ clknet_1_1__leaf_clk net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_14_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2653_ _0505_ _0506_ _0502_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2584_ net19 _0443_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1604_ _0760_ _0763_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1535_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1397_ _0559_ _0561_ _0564_ _0566_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
X_1466_ _0658_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2018_ _1205_ _1186_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2379__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2705_ net18 _0536_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2636_ _0927_ _0486_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2498_ _0285_ _1285_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1449_ _0610_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2567_ net4 _0442_ _0414_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_4_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2542__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1518_ _0663_ _0669_ _0710_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_2_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1575__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2352_ _0209_ _0212_ _0244_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2283_ c\[0\]\[6\] _0693_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2421_ _0185_ _0262_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _1150_ _1180_ _1186_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2619_ _0479_ _0480_ _0476_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ _1032_ _1107_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1852_ _0967_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1783_ _0972_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1548__A2 a\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2404_ _0295_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2266_ _0159_ _0160_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2335_ c\[0\]\[5\] _0969_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2197_ _0077_ _0082_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2120_ _1267_ _1289_ _1306_ _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_21_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer19 net98 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2051_ _1232_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1835_ _0948_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_32_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1904_ _1071_ _0610_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1697_ _0888_ _0614_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1766_ _0871_ _0955_ _0956_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2318_ _0173_ _0198_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2249_ _0764_ _0137_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput44 net44 x_end[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__1923__A2 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1551_ delta_t\[8\] _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1620_ _0554_ _0775_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1482_ _0634_ _0635_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2103_ _1220_ _1242_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2034_ _1157_ _1178_ _1221_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1818_ _1008_ _0910_ _0908_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ _0919_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1602__A1 _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1669__A1 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1841__A1 _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2721_ _0004_ clknet_1_1__leaf_clk net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2652_ net20 _0500_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1465_ _0657_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1603_ _0760_ _0763_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1534_ a\[0\]\[4\] _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2583_ _1082_ _0444_ _0454_ _0453_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2017_ _1150_ _1180_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_fanout54_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1396_ delta_t\[2\] _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0270_ _0541_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2635_ _0492_ _0493_ _0491_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2497_ _0382_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2566_ net3 _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2736__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1517_ _0692_ _0709_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1448_ b\[0\]\[1\] _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1379_ net36 _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_33_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2297__A1 c\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2049__A1 a\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0267_ _0273_ _0261_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2351_ _0215_ _0234_ _0243_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2282_ _0158_ _0161_ _0175_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ _1182_ _1185_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2212__A1 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2212__B2 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ net14 _0474_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2549_ _0596_ _0424_ _0430_ _0429_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input34_I y[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2690__A1 _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1851_ _0978_ _1039_ _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1920_ _1109_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2442__A1 _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ _0293_ _0294_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1782_ _0928_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2334_ _0225_ _0226_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2265_ c\[0\]\[4\] _0652_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2196_ _0087_ _0090_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2559__C _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ _1236_ _1237_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_32_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1834_ _0897_ _1024_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ _1091_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ _0874_ _0942_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1696_ a\[0\]\[6\] _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2317_ _0173_ _0198_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2248_ _0115_ _0141_ _0142_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2179_ delta_t\[0\] _1354_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_35_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput45 net45 x_end[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2645__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1620__A2 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1384__A1 _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1550_ _0588_ _0600_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_1481_ _0673_ _0615_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2102_ _1269_ _1274_ _1288_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2033_ _1160_ _1177_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1748_ _0921_ _0930_ _0939_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1611__A2 a\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1817_ _0554_ _0556_ _0906_ _0907_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_40_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1679_ _0794_ _0717_ _0768_ _0870_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_8_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2618__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1669__A2 _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _0003_ clknet_1_1__leaf_clk net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2651_ _1183_ _0498_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1602_ _0794_ _0659_ _0768_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2582_ net18 _0445_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1464_ _0639_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1533_ _0670_ _0691_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1395_ _0587_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2016_ _1202_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1832__A2 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2703_ _0542_ _0543_ _0540_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2565_ _0437_ _0440_ _0441_ _0436_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2634_ net11 _0489_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1516_ _0694_ _0708_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1378_ a\[1\]\[7\] b\[1\]\[7\] _0562_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2496_ _1290_ _0383_ _0384_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1447_ _0638_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1741__A1 b\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2049__A2 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2350_ _0235_ _0238_ _0242_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_2281_ _0174_ _0160_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1996_ _1183_ _1184_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ a\[1\]\[6\] _0465_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2548_ net17 _0425_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2479_ _0351_ _0361_ _0368_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_input27_I wbs_stb_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2726__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1850_ _0963_ _0976_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2442__A2 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1781_ _0695_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2402_ _0249_ _0250_ _0292_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2333_ _0220_ _0224_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ c\[0\]\[0\] _0922_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2195_ _0088_ _0089_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2681__A2 _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2197__A1 _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _1079_ _1167_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2121__A1 _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2424__A2 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2188__A1 _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ _0986_ _0633_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1833_ _0951_ _1023_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ _0874_ _0942_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2316_ _0176_ _0178_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1695_ _0803_ _0885_ _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2103__A1 _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2247_ _0118_ _0138_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2178_ t_reg\[0\] _1312_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput46 net46 x_start[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2590__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ _0672_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2581__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2032_ _1150_ _1218_ _1219_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2636__A2 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ _1281_ _1284_ _1287_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_17_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ _0931_ _0938_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1816_ _0905_ _0908_ _1005_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1678_ _0798_ _0828_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2572__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2627__A2 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1366__A2 _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2650_ _0503_ _0504_ _0502_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1601_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1532_ _0663_ _0669_ _0710_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2581_ _0897_ _0444_ _0452_ _0453_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_38_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1394_ _0586_ _0583_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_input1_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1463_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2015_ _1124_ _1189_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2779_ _0064_ net61 b\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2536__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2583__C _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1511__A2 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__I b\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2702_ net17 _0536_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2495_ _0357_ _0358_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2564_ _0573_ _0440_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1515_ _0697_ _0700_ _0707_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2527__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2633_ _0651_ _0486_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1377_ net33 _0569_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_4_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1446_ _0615_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1741__A2 _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout70 net71 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_24_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _0159_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2616_ _0477_ _0478_ _0476_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1995_ _1047_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2478_ _0363_ _0367_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1429_ delta_t\[7\] _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2547_ _0589_ _0424_ _0427_ _0429_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_38_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1780_ _0793_ _0934_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1402__A1 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2401_ _0249_ _0250_ _0292_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2332_ _0220_ _0224_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _0157_ _0658_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2194_ _0083_ _0086_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1978_ _1165_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2518__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2360__A2 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ _0954_ _0957_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1901_ _1000_ _1089_ _1090_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1763_ _0877_ _0953_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1694_ _0804_ _0805_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2315_ _0199_ _0202_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_27_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2246_ _0118_ _0138_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2177_ _1353_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_11_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2073__I _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput47 net47 x_start[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2100_ _1078_ _1230_ _1286_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2031_ _1154_ _1179_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1815_ _0905_ _0908_ _1005_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1746_ _0936_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1677_ _0792_ _0867_ _0868_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2229_ _0122_ _0658_ _0973_ _1356_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2739__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2012__A1 _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2315__A2 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1826__A1 b\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2003__A1 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1462_ _0654_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1600_ b\[0\]\[4\] _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2580_ _0409_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1531_ _0711_ _0712_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1393_ _0585_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2014_ _1126_ _1201_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2778_ _0063_ net64 b\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1729_ _0837_ _0842_ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_36_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2701_ _0260_ _0541_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _0487_ _0490_ _0491_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2494_ _0357_ _0358_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2563_ _0412_ _0439_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1445_ b\[0\]\[2\] _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2527__A2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1514_ _0701_ _0704_ _0706_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1376_ a\[1\]\[4\] b\[1\]\[4\] _0562_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1425__I a\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout71 net72 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout60 net72 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2445__A1 _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1994_ b\[0\]\[6\] _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ net13 _0474_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ _0313_ _0366_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1428_ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2546_ _0428_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_41_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1359_ a\[0\]\[0\] _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_21_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2675__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2695__B _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _1029_ _0252_ _0291_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_21_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1402__A2 _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2262_ c\[0\]\[5\] _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2331_ _0186_ _0223_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2193_ _0616_ _0636_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _0999_ _0775_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2529_ _0413_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input32_I y[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1880__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2648__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1831_ _0960_ _0978_ _1021_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_37_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__I _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1900_ _1001_ _1003_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1762_ _0878_ _0952_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1693_ _0804_ _0805_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2314_ _0865_ _0203_ _0206_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2245_ _0716_ _0139_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2176_ _1349_ _0822_ _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_35_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput48 net48 x_start[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput37 net37 wbs_ack_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_34_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ _1154_ _1179_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ _0933_ _0935_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1814_ _0906_ _0907_ _0619_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _0791_ _0857_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2228_ _0122_ _1356_ _0657_ _0973_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2159_ _1335_ _0683_ _1338_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_8_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2003__A2 _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1461_ _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2597__C _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1392_ _0584_ t_reg\[3\] _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
X_1530_ _0715_ _0719_ _0722_ _0663_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_10_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2013_ _1141_ _1188_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2777_ _0062_ net62 b\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1728_ _0836_ _0843_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_13_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1753__A1 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1659_ _0831_ _0851_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2729__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0531_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2631_ _0460_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2562_ _0438_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2401__B _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2493_ _0283_ _1244_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1513_ _0641_ _0705_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1444_ _0617_ _0636_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1375_ _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout61 net63 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout72 net75 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _1181_ _1100_ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2614_ a\[1\]\[5\] _0465_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2545_ net2 _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2684__A2 _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2476_ _0268_ _0355_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1358_ _0551_ net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1427_ _0619_ _0614_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2261_ _0151_ _0155_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2330_ _0221_ _0222_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2192_ _0083_ _0086_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _1163_ _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2354__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2528_ net24 _0406_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2459_ _0346_ _0348_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input25_I wbs_sel_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1830_ _0979_ _0980_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_32_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1761_ _0879_ _0915_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_25_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2584__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2313_ _0170_ _0204_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1692_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2639__A2 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2244_ _0115_ _0118_ _0138_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2175_ _1350_ _1351_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1959_ _1069_ _1097_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_16_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2575__A1 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput38 net38 x_end[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput49 net49 x_start[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_9_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1744_ _0933_ _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1813_ _1000_ _1001_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2557__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1780__A2 _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1675_ _0791_ _0857_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1534__I a\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2227_ c\[0\]\[4\] _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _1197_ _1133_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2158_ _0604_ _0628_ _1337_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2548__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1460_ _0652_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1391_ _0567_ _0578_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2012_ _1115_ _1198_ _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2185__I c\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2776_ _0061_ net61 b\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1727_ _0917_ _0918_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1658_ _0845_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_5_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1753__A2 _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2702__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1589_ _0773_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2492_ _0349_ _0369_ _0380_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1512_ _0646_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2561_ net26 _0406_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2630_ net6 _0489_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1374_ _0559_ _0561_ _0564_ _0566_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_2_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1443_ _0621_ _0634_ _0635_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2759_ _0044_ net58 a\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout62 net63 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout73 net75 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1653__A1 b\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ b\[0\]\[7\] _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2613_ _0473_ _0475_ _0476_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2475_ _0355_ _0364_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2544_ net16 _0425_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1357_ net27 net5 _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1426_ _0618_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2719__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2260_ _0152_ _0153_ _0154_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2191_ _0084_ _0085_ _0655_ _0659_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_28_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0838_ _0839_ _1082_ _0896_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2354__A2 _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2458_ _0322_ _0347_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1409_ _0568_ _0579_ _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2527_ net4 net3 _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input18_I wbs_dat_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2389_ _0236_ _0229_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1691_ _0729_ _0881_ _0882_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ _0869_ _0949_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2312_ _0205_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2243_ _0764_ _0137_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2174_ _1344_ _1347_ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2272__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput39 net39 x_end[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1958_ _1145_ _1146_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1889_ _1008_ _1005_ _1078_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__A1 _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1730__I _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2309__A2 _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1743_ _0695_ _0934_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1812_ _1002_ _0775_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1674_ _0853_ _0856_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_15_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2226_ _0095_ _0119_ _0120_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2493__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2646__I _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2157_ _1333_ _1336_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2088_ _1163_ _1229_ _1233_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1460__I _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ delta_t\[4\] _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2011_ _1119_ _1190_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _0060_ net67 b\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1657_ _0846_ _0849_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1588_ _0774_ _0780_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1726_ _0845_ _0850_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2376__I _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2209_ _0692_ _0103_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1441__A2 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2491_ _0351_ _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2560_ net7 _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1511_ b\[0\]\[0\] _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1442_ _0555_ _0610_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1373_ net34 _0565_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__2696__A1 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2758_ _0043_ net59 a\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2689_ net6 _0531_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_18_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1709_ _0894_ _0900_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout74 net75 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout63 net68 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1653__A2 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0460_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1991_ _1154_ _1179_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_15_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2474_ _0157_ _1285_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1425_ a\[0\]\[2\] _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2543_ _1314_ _0424_ _0426_ _0410_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_18_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A2 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1399__A1 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2190_ _1356_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_35_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1626__A2 _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1974_ _0727_ _0671_ _0840_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2457_ _0324_ _0328_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2388_ _0236_ _0229_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1408_ t_reg\[4\] _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2526_ _1349_ _0407_ _0411_ _0410_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_11_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1463__I _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1690_ net96 net95 _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2311_ _0170_ _0204_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2242_ _0121_ _0136_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2173_ _0744_ _0754_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1957_ _1048_ _1051_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2272__A2 _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2509_ _1289_ _0393_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1888_ _0618_ _1010_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input30_I y[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2791_ _0076_ net68 c\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1811_ _0672_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1673_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2199__I c\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1742_ _0835_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2225_ _0093_ _0101_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2662__I _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2087_ _1272_ _1273_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2156_ _0604_ _0628_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1756__A1 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_32_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2236__A2 c\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2010_ _1119_ _1190_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _0059_ net70 b\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1725_ _0834_ _0844_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1986__A1 a\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1656_ _0847_ _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1587_ _0778_ _0779_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2208_ _0092_ _0102_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2139_ delta_t\[2\] t_reg\[2\] _1312_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_27_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ _0361_ _0368_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1441_ _0557_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1510_ _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1372_ a\[1\]\[5\] b\[1\]\[5\] _0562_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2688_ _0531_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1423__A3 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ _0895_ _0899_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2757_ _0042_ net58 a\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1639_ _0778_ _0779_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout64 net66 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout75 net1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1990_ _1157_ _1178_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_15_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2611_ net12 _0474_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2542_ net11 _0425_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2742__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2473_ _0313_ _0317_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1424_ _0616_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_33_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2357__A1 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1399__A2 _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1973_ _1011_ _1161_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2587__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2525_ net23 _0407_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2456_ _0324_ _0345_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2387_ _0228_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1407_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2310_ _0864_ _0203_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2241_ _0125_ _0135_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2172_ delta_t\[9\] _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1956_ _1049_ _1050_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1887_ _1004_ _1012_ _1011_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2508_ _0394_ _0396_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ _0310_ _0320_ _0329_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_input23_I wbs_dat_i[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1741_ b\[0\]\[4\] _0932_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2790_ _0075_ net69 c\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1810_ _0728_ _0702_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1672_ _0619_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2224_ _0093_ _0101_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2155_ delta_t\[6\] _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2086_ _1261_ _1244_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1939_ _1127_ _1052_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1756__A2 _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2705__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ _0878_ _0879_ _0915_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2773_ _0058_ net69 b\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1655_ b\[0\]\[3\] _0705_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout73_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1586_ b\[0\]\[1\] _0702_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2069_ _1204_ _1256_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2207_ _0093_ _0095_ _0101_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2138_ _0589_ _0595_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1977__A2 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1371_ _0563_ net35 _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1440_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2687_ _0483_ _0405_ _0414_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1707_ _0897_ _0734_ _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2756_ _0041_ net59 a\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1638_ _0773_ _0781_ _0830_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1569_ _0677_ _0690_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout65 net66 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout54 net56 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2063__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ _0462_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2472_ _0261_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2541_ _0415_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1423_ _0555_ _0557_ _0610_ _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_38_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2357__A2 _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2739_ _0022_ clknet_1_0__leaf_clk t_reg\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2284__A1 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _1080_ _1086_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2455_ _1205_ _0327_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2524_ _0679_ _0407_ _0408_ _0410_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_11_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2386_ _0276_ _0241_ _0277_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1406_ delta_t\[4\] _0585_ _0594_ _0597_ _0598_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_14_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2732__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2524__C _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2240_ _0128_ _0134_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2171_ _1348_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_31_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1955_ _1142_ _1102_ _1143_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ _0995_ _1074_ _1075_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2438_ _0322_ _0324_ _0328_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_2507_ _0362_ _0366_ _0395_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input16_I wbs_dat_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2369_ _0260_ _0084_ _0222_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1755__I _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ _0647_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1671_ _0861_ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I wbs_dat_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2085_ _1270_ _1271_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2223_ _0116_ _0117_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2154_ _1334_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1869_ _1056_ _1057_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1938_ _1045_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2772_ _0057_ net63 b\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1723_ net90 _0884_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1654_ b\[0\]\[4\] _0642_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1395__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1371__A1 _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2206_ _0096_ _0098_ _0100_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1585_ b\[0\]\[0\] _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2068_ _1210_ _1212_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_fanout66_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ _1320_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2090__A2 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1370_ a\[1\]\[6\] b\[1\]\[6\] _0562_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2686_ _0529_ _0530_ _0526_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1637_ _0770_ _0782_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1706_ _0727_ _0632_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2755_ _0040_ net57 a\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1499_ _0670_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1568_ _0677_ _0690_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout55 net56 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout66 net68 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2471_ _0354_ _0356_ _0360_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1422_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2540_ _0416_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2738_ _0021_ clknet_1_0__leaf_clk t_reg\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2669_ _0517_ _0518_ _0516_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1583__I _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2293__A2 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__A2 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__A3 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1668__I _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1971_ _1158_ _1159_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2454_ _0342_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2385_ _0239_ _0240_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2523_ _0409_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1547__A1 a\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1405_ _0596_ _0595_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput1 wb_clk_i net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2202__I c\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2170_ _1344_ _1347_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1954_ _1099_ _1101_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1885_ _0998_ _1013_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ _1150_ _1180_ _0327_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2506_ _0312_ _0366_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2368_ _0099_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2299_ _0159_ _0192_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_34_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1998__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _0790_ _0859_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1922__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2222_ _0692_ _0103_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2084_ _1224_ _1240_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2153_ _1330_ _0628_ _1333_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1937_ _1055_ _1104_ _1125_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1856__I b\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ _1017_ _1018_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1799_ _0890_ _0988_ _0989_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2641__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2771_ _0056_ net73 b\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2632__A2 _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1653_ b\[0\]\[5\] _0696_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1722_ _0913_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1584_ _0776_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _0099_ _0639_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2067_ _1248_ _1254_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2136_ delta_t\[2\] _0595_ _1319_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_36_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2311__A1 _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2550__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2369__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1705_ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2754_ _0039_ net58 a\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ net15 _0522_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1567_ _0731_ _0739_ net87 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1636_ _0795_ _0798_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2119_ _1293_ _1296_ _1305_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1498_ _0674_ _0677_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_1_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout67 net68 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout56 net60 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2543__C _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _1220_ _1242_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_2_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2668_ net9 _0510_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2737_ _0020_ clknet_1_0__leaf_clk t_reg\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2599_ _0465_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1619_ _0618_ _0686_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__A3 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2520__A4 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1970_ _1088_ _1095_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2522_ net2 _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _0308_ _0330_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2384_ _0985_ _1016_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1404_ _0589_ _0592_ _0595_ _0596_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_11_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 wb_rst_i net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1953_ _1066_ _1098_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1884_ _0998_ _1013_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ _0268_ _0355_ _0315_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2436_ _0325_ _0326_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2367_ _0227_ _0230_ _0225_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2298_ c\[0\]\[4\] _0647_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1686__A1 b\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0583_ _0605_ _1332_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2221_ _0092_ _0102_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2083_ _1226_ _1239_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2402__A3 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1936_ _1043_ _1053_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1867_ _1019_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1798_ _0893_ _0912_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input21_I wbs_dat_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2419_ _0275_ _0289_ _0309_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1904__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2770_ _0055_ net73 b\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1721_ _0890_ _0893_ _0912_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_13_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1652_ _0834_ _0844_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1583_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2204_ c\[0\]\[3\] _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2135_ _1317_ _1318_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2066_ _1250_ _1253_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1919_ _1028_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_4_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2684_ b\[1\]\[7\] _0512_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2369__A2 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2753_ _0038_ net57 a\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1704_ a\[0\]\[3\] _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1566_ _0740_ _0741_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1497_ _0678_ _0688_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1635_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2118_ _1297_ _1303_ _1304_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_1_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ a\[0\]\[7\] _0703_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout68 net71 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout57 net59 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2735__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1420_ _0611_ net80 _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2667_ b\[1\]\[2\] _0513_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2736_ _0019_ clknet_1_0__leaf_clk t_reg\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1618_ _0740_ _0809_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2598_ _0404_ _0442_ _0439_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1549_ net98 _0612_ _0625_ _0733_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__2450__A1 _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2126__I _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2441__A1 _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ net22 _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2452_ _0310_ _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2383_ _0259_ _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1403_ delta_t\[3\] _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_34_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 wbs_adr_i[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2719_ _0002_ clknet_1_1__leaf_clk net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2423__A1 _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1952_ _1129_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_31_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1883_ _1070_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2435_ c\[0\]\[6\] _1047_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2504_ _0354_ _0391_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2366_ _0234_ _0243_ _0232_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2297_ c\[0\]\[5\] _0653_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2082_ _1220_ _1242_ _1268_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2220_ _0105_ _0113_ _0114_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2151_ _1328_ _1331_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _1121_ _1123_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1866_ _0985_ _1016_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1610__A2 a\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1797_ _0893_ _0912_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2418_ _0259_ _0274_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2349_ _0985_ _1016_ _0241_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA_input14_I wbs_dat_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1651_ _0836_ _0843_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1720_ _0901_ _0904_ _0911_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1582_ _0753_ _0755_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I wbs_dat_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2065_ _1127_ _1252_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2791__CLK net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ _0097_ _0643_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2134_ delta_t\[0\] t_reg\[0\] _0814_ _1315_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_29_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1918_ _1029_ _1032_ _1107_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1849_ _0979_ _0980_ _1020_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2683_ _0527_ _0528_ _0526_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ _0729_ _0802_ net97 _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1703_ _0727_ _0671_ _0632_ _0687_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2752_ _0037_ net57 a\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1496_ _0554_ _0632_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1565_ _0552_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2117_ _1044_ _1042_ _1252_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2048_ _1234_ _1235_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout69 net70 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net59 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ _0514_ _0515_ _0516_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2597_ _0437_ _0463_ _0464_ _0453_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1617_ _0807_ _0737_ _0734_ _0757_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2735_ _0018_ clknet_1_0__leaf_clk t_reg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1548_ _0686_ a\[0\]\[1\] _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1479_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2660__C _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2451_ _0319_ _0329_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2520_ _0404_ _0405_ net25 _0406_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_11_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1402_ _0590_ _0591_ t_reg\[2\] _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2382_ _0267_ _0273_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput4 wbs_adr_i[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _0001_ clknet_1_1__leaf_clk net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2725__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ net19 _0500_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__I c\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__C _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1951_ _1127_ _1139_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ _1071_ _0696_ _0993_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ _0235_ _0255_ _0256_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2434_ c\[0\]\[7\] _1100_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2503_ _0356_ _0360_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2296_ _0184_ _0189_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2081_ _1222_ _1241_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2150_ _0583_ _0605_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1934_ _1059_ _1121_ _1122_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_8_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1865_ _1054_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1796_ _0986_ _0639_ _0887_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2417_ _0305_ _0288_ _0307_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2348_ _0239_ _0240_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2571__A1 _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2279_ _0146_ _0164_ _0172_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2314__A1 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1650_ _0837_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1581_ b\[0\]\[2\] _0646_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2305__A1 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ c\[0\]\[2\] _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2064_ _1135_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2133_ delta_t\[1\] t_reg\[1\] _1312_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1917_ _1035_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1848_ _0979_ _1036_ _1037_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1779_ b\[0\]\[5\] _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2544__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2751_ _0036_ net61 bflip vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2573__C _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2682_ net14 _0522_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1633_ _0806_ _0811_ _0825_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1564_ _0753_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1702_ a\[0\]\[5\] _0609_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1495_ _0556_ _0687_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2116_ _1298_ _1299_ _1302_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_12_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2047_ _0888_ _0776_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout59 net60 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2734_ _0017_ clknet_1_0__leaf_clk t_reg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2665_ _0428_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2596_ a\[1\]\[0\] _0462_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1547_ a\[0\]\[2\] _0631_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1616_ _0808_ _0734_ _0757_ _0737_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_5_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1478_ a\[0\]\[3\] _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2450_ _0301_ _0338_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2381_ _0269_ _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1401_ _0589_ _0592_ _0593_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_11_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 wbs_cyc_i net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_34_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2717_ _0000_ clknet_1_1__leaf_clk net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2648_ _1046_ _0498_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2579_ net17 _0445_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1950_ _1135_ _1138_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_31_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2581__C _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__I b\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2502_ _0356_ _0360_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_24_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1881_ a\[0\]\[7\] _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2364_ _0238_ _0242_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2433_ _0269_ _0272_ _0323_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2295_ _0186_ _0187_ _0188_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_2_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2080_ _1212_ _1255_ _1266_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1933_ _1120_ _1103_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_33_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput30 y[1] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1864_ _1043_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1795_ _0888_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2416_ _0278_ _0306_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2347_ c\[0\]\[7\] _0693_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2278_ _0149_ _0163_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1834__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__A2 _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2738__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1600__I b\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _0701_ _0771_ _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_13_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2201_ _0078_ _0932_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2132_ _1316_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _1046_ _1133_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_14_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1916_ _1038_ _1105_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1847_ _0980_ _1020_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _0932_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2516__I _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2681_ b\[1\]\[6\] _0512_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2750_ _0035_ net55 delta_t\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1701_ net85 _0891_ _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1494_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1632_ _0812_ _0813_ _0824_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1563_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2115_ _1217_ _1247_ _1301_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2046_ _1163_ _1166_ _1233_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__A1 _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2664_ net8 _0510_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2733_ _0016_ clknet_1_0__leaf_clk t_reg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2595_ _0462_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1546_ _0732_ _0736_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1477_ _0617_ _0636_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1615_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _1216_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2435__A1 c\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0174_ _0271_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1400_ _0590_ _0591_ delta_t\[1\] t_reg\[0\] _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xinput6 wbs_dat_i[0] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2647_ _0499_ _0501_ _0502_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2716_ _0027_ net55 delta_t\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1529_ _0720_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2578_ _0449_ _0451_ _0423_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2408__A1 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_31_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1880_ _0986_ _0652_ _0991_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2501_ _0361_ _0368_ _0389_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2363_ _0238_ _0242_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2432_ _0236_ _0271_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2294_ _0080_ _0777_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput31 y[2] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1932_ _1120_ _1103_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1863_ _1045_ _1052_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xinput20 wbs_dat_i[6] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2415_ _0282_ _0288_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1794_ _0984_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2346_ c\[0\]\[6\] _0654_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2277_ _0870_ _0123_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1834__A2 _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1761__A1 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2062_ _1042_ _1249_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2200_ _0094_ _0735_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2131_ _1313_ _1315_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_29_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1846_ _0980_ _1020_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1915_ _1041_ _1055_ _1104_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1777_ _0925_ _0964_ _0966_ _0967_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1504__A1 _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2329_ _0097_ _0922_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input12_I wbs_dat_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__A1 _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_31_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2680_ _0524_ _0525_ _0526_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1631_ _0819_ _0823_ a\[0\]\[0\] _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1700_ net99 _0825_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1493_ _0682_ _0685_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_1_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1562_ delta_t\[9\] _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2114_ _1215_ _1300_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I wbs_adr_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ _1029_ _0673_ _0841_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2728__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1829_ _0985_ _1016_ _1019_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_32_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__I c\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2690__C _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2732_ _0015_ clknet_1_1__leaf_clk net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2663_ b\[1\]\[1\] _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2594_ _0404_ _0442_ _0438_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1707__A1 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ a\[0\]\[1\] _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1545_ _0737_ _0735_ _0689_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_5_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1476_ _0649_ _0668_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_37_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2028_ _1131_ _1138_ _1134_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_20_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 wbs_dat_i[16] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer2_I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2646_ _0460_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2577_ net16 _0450_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2715_ _0026_ net54 delta_t\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1459_ _0642_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1528_ _0715_ _0719_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2431_ _1142_ _0287_ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2500_ _0388_ _0367_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2335__A1 c\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2583__A1 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2362_ _0176_ net82 _0244_ _0253_ net76 _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_2293_ _0130_ _0703_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2638__A2 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1377__A2 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2629_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1368__A2 _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1614__I a\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput32 y[3] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1931_ _1062_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput21 wbs_dat_i[7] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1862_ _1048_ _1051_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1793_ net91 _0981_ _0982_ _0983_ _0879_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_12_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 wbs_dat_i[19] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2414_ _0282_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2345_ _0236_ _0192_ _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2276_ _0713_ _0166_ _0169_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1761__A2 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2061_ _1127_ _1139_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2710__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2130_ _1314_ _0592_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1914_ _1059_ _1062_ _1103_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_29_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1845_ _0960_ _1033_ _1034_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1776_ _0927_ _0925_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2328_ _0130_ _0777_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2701__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1504__A2 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2259_ _0078_ _0928_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1743__A2 _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1630_ _0820_ _0821_ _0822_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_39_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1492_ _0625_ _0630_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1561_ _0573_ t_reg\[8\] _0584_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2113_ _1217_ _1247_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2044_ _1228_ _1231_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ _1017_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1759_ _0866_ _0943_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2731_ _0014_ clknet_1_1__leaf_clk net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2662_ _0512_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2593_ _0458_ _0459_ _0461_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1613_ _0803_ _0804_ _0805_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1544_ _0552_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ _0651_ _0656_ _0666_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_37_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2027_ _1205_ _1213_ _1214_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout55_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2538__I _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2718__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 wbs_dat_i[17] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0549_ _0550_ _0410_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2183__I c\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2645_ net18 _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2576_ _0404_ _0405_ _0419_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1527_ _0666_ _0667_ _0668_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1389_ _0581_ delta_t\[6\] _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1458_ _0650_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1616__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1919__A2 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2041__A1 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2032__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ _0234_ _0243_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2430_ _0284_ _0286_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2292_ _0185_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input35_I y[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2628_ _0419_ _0484_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2559_ _0747_ _0417_ _0435_ _0436_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1837__A1 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1930_ _1117_ _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2005__A1 _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 y[4] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 wbs_dat_i[1] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput22 wbs_dat_i[8] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1861_ _1049_ _1050_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1792_ _0880_ _0883_ _0913_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2413_ _0258_ _0302_ _0303_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2344_ _0191_ _0193_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2275_ _0140_ _0167_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2060_ _1215_ _1217_ _1247_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2474__A1 _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1913_ _1066_ _1098_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_29_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2226__A1 _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1844_ _0954_ _1022_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1775_ _0926_ _0965_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_12_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2258_ _0097_ _0835_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2327_ _0186_ _0218_ _0219_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2189_ _0078_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0743_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_39_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2112_ _1131_ _1251_ _1134_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1491_ _0622_ _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2447__A1 _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2043_ _1080_ _1230_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1827_ b\[0\]\[7\] _0658_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1689_ net86 _0826_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1758_ _0866_ _0943_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2730_ _0013_ clknet_1_1__leaf_clk net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2661_ _0439_ _0484_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_14_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2592_ _0460_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1612_ _0671_ net79 _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1543_ _0553_ _0735_ _0689_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1474_ _0660_ _0664_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _1182_ _1185_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1882__A2 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 wbs_dat_i[18] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2644_ _0488_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2713_ net21 _0535_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1808__I a\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2575_ _0865_ _0448_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1457_ _0641_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1526_ _0667_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1388_ _0568_ _0579_ _0580_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_37_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2009_ _1155_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1453__I _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0199_ _0202_ _0245_ _0251_ _0212_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2291_ c\[0\]\[1\] _0841_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1543__A1 _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2408__B _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2099__A2 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2627_ _0660_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2489_ _0344_ _0370_ _0377_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2558_ _0409_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input28_I wbs_we_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1509_ _0687_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1837__A2 _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1860_ _0695_ _0923_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput34 y[5] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 wbs_dat_i[9] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ _0884_ _0914_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 wbs_dat_i[20] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2274_ _0168_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2412_ _0257_ _0290_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2343_ _0174_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _1160_ _1177_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2562__I _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__A2 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1843_ _0978_ _1021_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1912_ _1099_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1774_ _0927_ _0923_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2326_ _0187_ _0188_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2257_ _0099_ _0647_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2188_ _0077_ _0082_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_18_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2392__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1490_ _0624_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ _1181_ _1244_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2042_ _1165_ _1229_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1826_ b\[0\]\[6\] _0654_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1757_ _0863_ _0945_ _0947_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1688_ _0797_ _0827_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2309_ _0199_ _0202_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_input10_I wbs_dat_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1949__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2677__A2 _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0437_ _0510_ _0511_ _0422_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1611_ _0608_ a\[0\]\[4\] _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2591_ net2 _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1542_ _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_1473_ _0651_ _0664_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2025_ _1186_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input2_I wb_rst_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2789_ _0074_ net74 c\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2741__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1809_ _0999_ _0633_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A1 c\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2643_ _0794_ _0498_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2712_ _0283_ _0541_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2574_ _0443_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1387_ t_reg\[5\] _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1525_ _0716_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1456_ _0640_ _0644_ _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2008_ _1113_ _1195_ _1193_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ _0182_ _0154_ _0183_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_22_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2559__A1 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0485_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2557_ net21 _0416_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2488_ _0340_ _0371_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1508_ _0638_ _0643_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1439_ net78 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1790_ _0884_ _0914_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput13 wbs_dat_i[21] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 y[6] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2411_ _0275_ _0289_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xinput24 wbs_sel_i[0] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ _0952_ _0177_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2713__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2273_ _0140_ _0167_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1988_ _1169_ _1176_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2609_ a\[1\]\[4\] _0466_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2704__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1842_ _0957_ _1030_ _1031_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1911_ b\[0\]\[6\] _1100_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1773_ _0926_ _0929_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_12_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2325_ _0187_ _0188_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2256_ _0131_ _0150_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2187_ _0079_ _0081_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1967__A2 _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2110_ _1183_ _1285_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2041_ _1113_ _1084_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _1015_ _0981_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1756_ _0865_ _0944_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ _0726_ _0796_ _0828_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_2308_ _0145_ _0200_ _0201_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2393__I c\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2239_ _0129_ _0133_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2071__A1 _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1949__A2 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2590_ net21 _0450_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1610_ _0613_ a\[0\]\[5\] _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1541_ net88 _0733_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1472_ _0660_ _0654_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2024_ _1141_ _1188_ _1211_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_20_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1739_ b\[0\]\[5\] _0653_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2788_ _0073_ net70 c\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1808_ a\[0\]\[5\] _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1858__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2283__A1 c\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2711_ _0547_ _0548_ _0540_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2642_ _0485_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2573_ _0808_ _0444_ _0447_ _0436_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1524_ _0664_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1455_ _0645_ _0647_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1386_ _0578_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2007_ _1115_ _1191_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2017__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2265__A1 c\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2008__A1 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2487_ _0337_ _0374_ _0375_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0414_ _0484_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2556_ _0433_ _0434_ _0423_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1507_ _0640_ _0698_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_37_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1369_ bflip _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1438_ _0625_ _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput36 y[7] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 wbs_sel_i[1] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput14 wbs_dat_i[22] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2410_ net81 _0300_ _0297_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2341_ _0232_ _0233_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2272_ _0808_ _0166_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1987_ _1174_ _1175_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input33_I y[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2608_ _0471_ _0472_ _0461_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2539_ _0418_ _0421_ _0423_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2640__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ _0969_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1841_ _0951_ _1023_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1772_ _0961_ _0939_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2324_ _0190_ _0194_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2255_ _0129_ _0133_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2186_ _0080_ _0657_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2689__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ _1011_ _1227_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _0946_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1686_ b\[0\]\[6\] _0693_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ _0987_ _0990_ _1014_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2238_ _0131_ _0132_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2307_ _0143_ _0165_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2169_ _1342_ _1345_ _1346_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1646__A2 _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1540_ delta_t\[8\] _0681_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1471_ _0659_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2023_ _1129_ _1140_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1807_ _0901_ _0996_ _0997_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1738_ _0926_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2787_ _0072_ net69 c\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1669_ _0713_ _0858_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1555__A1 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2710_ net20 _0535_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A2 _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2641_ _0496_ _0497_ _0491_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1454_ _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1523_ _0557_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2572_ net11 _0445_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1385_ _0570_ _0572_ _0575_ _0577_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_42_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ _1193_ _1194_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2265__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ _0483_ _0442_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2486_ _0334_ _0372_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1437_ net77 net83 _0626_ _0627_ _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_10_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1506_ _0644_ _0648_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2555_ net20 _0420_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1368_ net30 _0560_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_18_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2592__I _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput26 wbs_sel_i[2] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 wbs_dat_i[23] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2340_ _0216_ _0217_ _0231_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2271_ _0143_ _0165_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ a\[0\]\[7\] _0646_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2607_ net10 _0463_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2468__A2 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2469_ _0357_ _0358_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2538_ _0422_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input26_I wbs_sel_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2721__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1840_ _0954_ _1022_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_29_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ _0921_ _0930_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2323_ _0184_ _0189_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2254_ _0147_ _0148_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2185_ c\[0\]\[2\] _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2744__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1969_ _1077_ _1087_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1823_ _0995_ _0998_ _1013_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_25_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1685_ _0875_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1754_ _0863_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2237_ _0130_ _0643_ _0705_ _0097_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2306_ _0146_ _0164_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2168_ _0622_ _0745_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2099_ _0864_ _1285_ _0905_ _1230_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_31_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1470_ _0637_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2708__C _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2022_ _1207_ _1209_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2589__A1 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2786_ _0071_ net69 c\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1806_ _0904_ _0911_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1668_ _0860_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1737_ _0927_ _0928_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1599_ _0725_ _0787_ _0788_ _0724_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_36_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2640_ net17 _0489_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1522_ _0617_ _0714_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_10_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2571_ _0553_ _0444_ _0446_ _0436_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1453_ _0633_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1384_ _0576_ net32 _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2005_ _1111_ _1112_ _1192_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1584__I _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2769_ _0054_ net73 b\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ net4 _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _1335_ _0417_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2485_ _0334_ _0372_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1367_ a\[1\]\[1\] b\[1\]\[1\] bflip _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1436_ delta_t\[6\] _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1505_ _0644_ _0648_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2707__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput16 wbs_dat_i[2] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput27 wbs_stb_i net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2270_ _0145_ _0146_ _0164_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1985_ _1172_ _1173_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2606_ a\[1\]\[3\] _0466_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2537_ _0409_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2399_ _0254_ _0257_ _0290_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2468_ _0285_ _1137_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1419_ delta_t\[5\] _0602_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input19_I wbs_dat_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ _0921_ _0930_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2322_ _0213_ _0197_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2184_ _0078_ _0653_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2253_ _0125_ _0135_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__I _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1968_ _1093_ _1094_ _1156_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1899_ _1001_ _1003_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2310__A2 _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1753_ _0865_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1822_ _1004_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1684_ _0846_ _0849_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_13_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2305_ _0171_ _0173_ _0198_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2236_ _0130_ c\[0\]\[2\] _0642_ _0705_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2167_ _0622_ _0745_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2098_ _1133_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1803__A1 a\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ _1144_ _1208_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2734__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1736_ _0777_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2785_ _0070_ net63 c\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1805_ _0904_ _0911_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1598_ _0784_ _0786_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1667_ _0790_ _0859_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_36_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ _0091_ _0104_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ net6 _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1383_ a\[1\]\[3\] b\[1\]\[3\] _0573_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1452_ b\[0\]\[0\] _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1521_ _0557_ _0656_ _0664_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2004_ _1111_ _1112_ _1192_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2699_ _0538_ _0539_ _0540_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2768_ _0053_ net73 b\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1719_ _0909_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _0481_ _0482_ _0476_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1504_ _0695_ _0696_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2553_ _1330_ _0417_ _0432_ _0429_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1366_ net31 _0558_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2484_ _0373_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1435_ _0581_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2652__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1391__A1 _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2643__A1 _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 wbs_dat_i[3] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput28 wbs_we_i net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1382__A1 _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2634__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1984_ _0888_ _0702_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2467_ _0283_ _1184_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2605_ _0469_ _0470_ _0461_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2536_ net6 _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2398_ _0258_ _0275_ _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1418_ _0588_ _0600_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2124__I _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _0181_ _0196_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2252_ _0128_ _0134_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2183_ c\[0\]\[1\] _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1155_ _0932_ _1091_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1898_ _1077_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input31_I y[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2519_ net28 net37 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__1649__A2 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1812__A2 _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1683_ _0847_ _0848_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A1 b\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1821_ _1006_ _1007_ _1009_ _1011_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_1752_ _0866_ _0869_ _0943_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_2304_ _0176_ _0178_ _0197_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_29_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2235_ c\[0\]\[3\] _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2166_ _0744_ _0754_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2097_ _1282_ _1283_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1778__I _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2047__A2 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2020_ _1147_ _1187_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2784_ _0069_ net74 c\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1735_ _0638_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1666_ _0713_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1804_ _0993_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1597_ _0553_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2218_ _0090_ _0106_ _0112_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2149_ _0604_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2201__A2 _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A1 b\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1520_ _0555_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1382_ _0574_ net29 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1451_ _0641_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2003_ _1113_ _1115_ _1191_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_26_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2767_ _0052_ net66 a\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2698_ _0428_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1649_ b\[0\]\[0\] _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1718_ _0619_ _0776_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__I a\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2498__A2 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2724__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2186__A1 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2127__I _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2483_ _0334_ _0337_ _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2621_ net15 _0474_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1503_ _0615_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ net19 _0416_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1365_ a\[1\]\[2\] b\[1\]\[2\] bflip _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1434_ delta_t\[6\] _0581_ _0602_ delta_t\[5\] _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__1391__A2 _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 wbs_dat_i[4] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput29 y[0] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ net9 _0463_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1983_ _1081_ _1170_ _1171_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1373__A2 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2466_ _0314_ _0355_ _0315_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1417_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2570__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2535_ _0412_ _0419_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2397_ _0278_ _0282_ _0288_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_14_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2313__A1 _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2405__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2320_ _0176_ _0178_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2251_ _0798_ _0828_ _0123_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__2552__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ _1356_ _0969_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _0986_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1897_ _1080_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2449_ _0304_ _0331_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input24_I wbs_sel_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ net3 _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0864_ _1010_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_17_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1682_ _0872_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1751_ _0871_ _0874_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1576__A2 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2303_ _0181_ _0196_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2234_ c\[0\]\[1\] _0835_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2525__A1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2165_ _1343_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2096_ _1232_ _1238_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1949_ _1046_ _1137_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2783_ _0068_ net67 b\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1803_ a\[0\]\[7\] _0614_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1734_ _0924_ _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1596_ _0724_ _0788_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1665_ _0791_ _0792_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_13_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout74_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ _0108_ _0109_ _0111_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2079_ _1210_ _1265_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2148_ _1329_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1450_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1400__A1 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1381_ a\[1\]\[0\] b\[1\]\[0\] _0573_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2002_ _1119_ _1190_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2766_ _0051_ net65 a\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2697_ net16 _0536_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1579_ _0704_ _0706_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_6_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1717_ _0905_ _0908_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1648_ _0840_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2110__A2 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ a\[1\]\[7\] _0465_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2571__C _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2482_ _0340_ _0371_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1502_ b\[0\]\[3\] _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1433_ _0582_ _0612_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2551_ _1325_ _0424_ _0431_ _0429_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_37_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1364_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1860__A1 _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2749_ _0034_ net57 delta_t\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_14_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1892__I a\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1679__A1 _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput19 wbs_dat_i[5] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1842__A1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1982_ _1002_ _1084_ _1083_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2603_ a\[1\]\[2\] _0466_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2534_ _0413_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2396_ _1066_ _1098_ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2465_ _0316_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1416_ _0608_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1833__A1 _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2086__A1 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2561__A2 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2077__A1 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2250_ _0121_ _0136_ _0144_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2181_ c\[0\]\[0\] _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2737__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1965_ _1073_ _1152_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_7_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2517_ net4 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1896_ _1081_ _1083_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2448_ _0304_ _0331_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2379_ _0270_ _1136_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I wbs_dat_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2059__A1 _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2298__A1 c\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2470__A1 _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1750_ _0877_ _0916_ _0941_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _0829_ _0852_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2302_ _0195_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2233_ _0096_ _0126_ _0127_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input9_I wbs_dat_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2164_ _0747_ _0745_ _1342_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2095_ _1228_ _1231_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1948_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1879_ _0987_ _1067_ _1068_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_16_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2680__B _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2691__A1 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2782_ _0067_ net65 b\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ _0650_ _0645_ _0922_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_25_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1802_ _0991_ _0992_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_25_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1595_ _0725_ _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1664_ _0853_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout67_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2682__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2147_ _1325_ _0605_ _1328_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2216_ _0110_ _0107_ _0715_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2078_ _1212_ _1255_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2434__A1 c\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2425__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1380_ bflip _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1400__A2 _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2001_ _1124_ _1189_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2765_ _0050_ net66 a\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2696_ _0080_ _0532_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1716_ _0906_ _0907_ _0555_ _0556_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_13_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1578_ _0704_ _0706_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1647_ _0838_ _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2655__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer20 _0826_ net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2550_ net18 _0425_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2481_ _0344_ _0370_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1432_ _0622_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1363_ a\[0\]\[0\] _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1501_ _0650_ _0693_ _0649_ _0665_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__2637__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2679_ _0428_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2748_ _0033_ net55 delta_t\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1981_ _1002_ _1084_ _1083_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_15_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2602_ _0467_ _0468_ _0461_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2533_ delta_t\[0\] _0417_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2395_ _0284_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2464_ _1205_ _0352_ _0353_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1415_ net94 _0607_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_3_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A1 _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2683__B _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1521__B2 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2180_ _1355_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__I _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _1076_ _1151_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1895_ _1002_ _1084_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2516_ _0403_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2447_ _0299_ _0335_ _0336_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2378_ _0122_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_3_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2301_ _0190_ _0194_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1680_ _0831_ _0851_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2232_ _0098_ _0100_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2163_ _1335_ _0683_ _1341_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_28_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _1275_ _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1947_ _0973_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1878_ _0990_ _1014_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2517__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2727__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2781_ _0066_ net65 b\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1732_ _0650_ _0645_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1663_ _0764_ _0854_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1801_ a\[0\]\[6\] _0609_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1594_ _0784_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2077_ _1261_ _1263_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2146_ delta_t\[3\] _0586_ _1327_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2215_ _0086_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1945__A1 _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A2 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ _1126_ _1141_ _1188_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2585__C _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2764_ _0049_ net64 a\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2695_ _0534_ _0537_ _0526_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1646_ t_reg\[9\] _0814_ _0815_ _0818_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1715_ _0823_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1577_ _0768_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xrebuffer10 _0806_ net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer21 _0802_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_2129_ delta_t\[1\] _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1918__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2686__B _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1909__A1 b\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2480_ _0349_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1500_ _0657_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2582__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1431_ _0568_ _0579_ _0623_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1362_ _0554_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2678_ net13 _0522_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2747_ _0032_ net54 delta_t\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1629_ t_reg\[9\] _0584_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2573__A1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ _1162_ _1168_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xrebuffer1 _0215_ net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2463_ _0325_ _0326_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2601_ net8 _0463_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2532_ _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2555__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2394_ _0285_ _1100_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1414_ _0588_ _0600_ _0603_ _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2760__CLK net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1597__A2 _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ _1076_ _1151_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2528__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1894_ _0840_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2446_ _0332_ _0296_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2515_ _0716_ _0139_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2377_ _0268_ net93 _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2300_ _0191_ _0193_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2231_ _0098_ _0100_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2093_ _1276_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2162_ _1338_ _1340_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2623__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1946_ _1132_ _1134_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1877_ _0990_ _1014_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input22_I wbs_dat_i[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1724__A2 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2429_ _0319_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1800_ _0894_ _0900_ _0895_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2780_ _0065_ net64 b\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1731_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1662_ _0767_ _0783_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2214_ _0094_ _0716_ _0717_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1593_ _0692_ _0709_ _0785_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2076_ _1200_ _1257_ _1262_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2145_ _1326_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1929_ _1038_ _1105_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2370__A2 _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2763_ _0048_ net61 a\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2694_ net11 _0536_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1576_ b\[0\]\[4\] _0696_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1645_ _0820_ _0821_ _0822_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1714_ _0819_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 net92 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout72_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2059_ _1220_ _1242_ _1246_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xrebuffer22 _0826_ net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2128_ delta_t\[0\] t_reg\[0\] _1312_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1909__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1430_ t_reg\[6\] _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1361_ a\[0\]\[1\] _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2631__I _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2746_ _0031_ net54 delta_t\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2677_ b\[1\]\[5\] _0512_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1559_ _0746_ _0749_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1628_ _0743_ _0752_ _0756_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2089__A1 _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1827__A1 b\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2004__A1 _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ a\[1\]\[1\] _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer2 _0587_ net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2462_ _0325_ _0326_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2393_ c\[0\]\[6\] _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1413_ _0604_ _0605_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2531_ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ _0012_ clknet_1_1__leaf_clk net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2234__A1 c\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _1096_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2181__I c\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__A2 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1893_ _1082_ _0757_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_11_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2514_ _0402_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2445_ _0296_ _0332_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2376_ _0157_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_3_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2519__A2 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2230_ _0123_ _0124_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2694__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2092_ _1277_ _1278_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2161_ _1335_ _0683_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1945_ _0794_ _0972_ _1133_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1724__A3 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1876_ _0984_ _1064_ _1065_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2685__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2359_ _0209_ _0244_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2428_ _0311_ _0318_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2437__A1 _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I wbs_dat_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ _0841_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ _0767_ _0783_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1592_ _0694_ _0708_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input7_I wbs_dat_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2144_ delta_t\[3\] _0586_ _1323_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2213_ _0715_ _0107_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2075_ _1202_ _1203_ _1256_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1928_ _1041_ _1116_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ _0793_ _0928_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2762_ _0047_ net64 a\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _0808_ _0737_ _0838_ _0839_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2693_ _0535_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1575_ b\[0\]\[3\] _0652_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1644_ _0641_ _0776_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer12 net100 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer23 _0582_ net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2127_ _0814_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2058_ _1243_ _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2274__I _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1360_ _0552_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2676_ _0521_ _0523_ _0516_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0030_ net54 delta_t\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1489_ _0679_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1558_ _0684_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1627_ _0815_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer3 _0631_ net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2530_ _0412_ _0414_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2392_ _0283_ _0655_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2461_ _0320_ _0329_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1412_ _0602_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ _0011_ clknet_1_1__leaf_clk net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2659_ b\[1\]\[0\] _0509_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1809__A2 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1961_ _1066_ _1148_ _1149_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1892_ a\[0\]\[4\] _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2513_ _0376_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2444_ _1197_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2375_ _0261_ _0266_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2207__A2 _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _1339_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2446__A2 _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1361__I a\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2091_ _1071_ _1184_ _1236_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1944_ _1130_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1875_ _1063_ _1015_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2427_ _0313_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ _0207_ _0247_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2289_ _0152_ _0153_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2373__A1 _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2125__A1 _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1591_ _0764_ _0767_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1660_ _0829_ _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2143_ _0583_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2212_ _0085_ _0656_ _0717_ _0084_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_36_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2074_ _1071_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _1055_ _1104_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1858_ _1046_ _1047_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1975__B _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1789_ _0931_ _0938_ _0936_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2346__A1 c\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2740__CLK clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2761_ _0046_ net62 a\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2692_ _0483_ _0405_ _0419_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1643_ _0638_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1712_ _0812_ _0902_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2585__A1 _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1574_ _0697_ _0765_ _0766_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2126_ _1311_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2057_ _1183_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer13 net89 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xrebuffer24 _0811_ net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_13_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1379__A2 _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2567__A1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2319__A1 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2675_ net12 _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1626_ t_reg\[9\] _0814_ _0815_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_14_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0029_ net56 delta_t\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1488_ _0568_ _0579_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1557_ _0744_ _0681_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2109_ _1294_ _1295_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2460_ _0311_ _0318_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer4 net78 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2391_ c\[0\]\[7\] _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2712__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1411_ delta_t\[5\] _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_14_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _0010_ clknet_1_1__leaf_clk net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2658_ _0509_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2589_ _1261_ _0448_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1609_ _0799_ _0800_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1449__I _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1960_ _1069_ _1097_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1891_ _0999_ _0687_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2443_ _0333_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2512_ _1261_ _0378_ _0400_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_11_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2374_ _0185_ _0223_ _0264_ _0265_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_3_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1718__A2 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2090_ _1155_ _1137_ _1234_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1642__I _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1654__A1 b\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1943_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1874_ _1063_ _1015_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2426_ _0314_ _0316_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_39_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2357_ _0673_ _0246_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2288_ _0152_ _0153_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1893__A1 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2373__A2 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2125__A2 _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ _0770_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2073_ _1260_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_28_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2211_ _0088_ _0089_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2142_ _1324_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1926_ _1032_ _1107_ _1114_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1788_ _0878_ _0952_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1857_ _0934_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_12_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2409_ _0257_ _0290_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input20_I wbs_dat_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__A1 c\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2691_ _0084_ _0532_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2760_ _0045_ net56 a\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1642_ _0703_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1711_ _0813_ _0824_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1573_ _0700_ _0707_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2056_ _1136_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer14 _0685_ net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xrebuffer25 _0759_ net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2125_ _0553_ _0789_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1909_ b\[0\]\[7\] _0655_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2264__A1 c\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput50 net50 x_start[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2007__A1 _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2743_ _0028_ net58 delta_t\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2674_ _0509_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1556_ _0629_ _0748_ _0627_ _0682_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1625_ _0816_ _0817_ _0755_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1487_ t_reg\[7\] _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2730__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2108_ _1248_ _1254_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2039_ _1080_ _1167_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2391__I c\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2566__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer5 _0612_ net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1410_ delta_t\[5\] _0602_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2390_ _0279_ _0280_ _0281_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2726_ _0009_ clknet_1_1__leaf_clk net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2400__A1 _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2657_ _0439_ _0484_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2588_ _0456_ _0457_ _0423_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1539_ _0678_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1608_ _0739_ _0759_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2467__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1442__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_0_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1890_ _1079_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2630__A1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2442_ _0296_ _0299_ _0332_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2511_ _0381_ _0386_ _0399_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2373_ _0260_ _1137_ _0222_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2697__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1375__I _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2621__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2709_ _0285_ _0541_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _0793_ _0972_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ _0884_ _0914_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2356_ _0248_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2425_ _0270_ _0085_ _0906_ _0907_ _0315_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__2134__A3 _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2287_ _0179_ _0180_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2210_ _0091_ _0104_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2072_ _1196_ _1259_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_36_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2141_ delta_t\[3\] _0586_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1925_ _1035_ _1106_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1856_ b\[0\]\[5\] _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2408_ _1082_ _0297_ _0298_ _0293_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2339_ _0216_ _0217_ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input13_I wbs_dat_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__A2 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__A3 _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2690_ _0094_ _0532_ _0533_ _0422_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1793__B2 _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1710_ _0813_ _0824_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1572_ _0700_ _0707_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1641_ _0832_ _0833_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2124_ _1310_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input5_I wbs_cyc_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2055_ _1181_ _1184_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer15 _0880_ net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1908_ _1069_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1839_ _0728_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput51 net51 x_start[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput40 net40 x_end[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ _0025_ clknet_1_0__leaf_clk t_reg\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_14_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ b\[1\]\[4\] _0513_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ _0747_ _0624_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1624_ _0746_ _0749_ _0751_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2191__A1 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2107_ _1250_ _1253_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout63_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1486_ delta_t\[8\] _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2038_ _1169_ _1176_ _1225_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer6 _0254_ net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2725_ _0008_ clknet_1_1__leaf_clk net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2656_ _0507_ _0508_ _0502_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1739__A1 b\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1911__A1 b\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2164__A1 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1538_ _0729_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1607_ _0759_ _0739_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1469_ _0649_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2587_ net20 _0450_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2467__A2 _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0387_ _0390_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_11_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2720__CLK clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2441_ _0301_ _0304_ _0331_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2372_ _0185_ _0263_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_19_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2708_ _0268_ _0532_ _0546_ _0422_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2639_ _0972_ _0486_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1872_ _0970_ _1060_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1941_ _0923_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_16_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1386__I _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2355_ _0207_ _0247_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2286_ _0156_ _0162_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2424_ _0270_ _0085_ _1130_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_39_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2521__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _1319_ _1321_ _1322_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2071_ _1197_ _1258_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1855_ _0967_ _1044_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2714__B _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1924_ _0999_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1786_ _0963_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2407_ _0252_ _0291_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2512__A1 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2338_ _0227_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2269_ _0149_ _0163_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__2579__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1571_ _0726_ _0760_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1640_ _0774_ _0780_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2123_ _1264_ _1307_ _1309_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xrebuffer16 net90 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ _1222_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_17_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1481__A1 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1838_ _0948_ _1025_ _1027_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1907_ _1073_ _1076_ _1096_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_17_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1769_ _0958_ _0941_ _0959_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xoutput52 net52 x_start[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput41 net41 x_end[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _0519_ _0520_ _0516_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2741_ _0024_ clknet_1_0__leaf_clk t_reg\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1554_ delta_t\[7\] _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1485_ _0618_ _0608_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1623_ _0588_ _0600_ _0742_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2191__A2 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

